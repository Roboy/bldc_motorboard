-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Aug 26 2019 01:17:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__37951\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n6111_cascade_\ : std_logic;
signal \c0.n5758_cascade_\ : std_logic;
signal \c0.n5761\ : std_logic;
signal \c0.data_in_frame_18_1\ : std_logic;
signal \c0.data_in_frame_19_1\ : std_logic;
signal \c0.n6303_cascade_\ : std_logic;
signal \c0.n6057_cascade_\ : std_logic;
signal \c0.n6306\ : std_logic;
signal \c0.n6060_cascade_\ : std_logic;
signal \c0.n6087\ : std_logic;
signal \c0.n5770\ : std_logic;
signal \c0.n5788_cascade_\ : std_logic;
signal \c0.n6027_cascade_\ : std_logic;
signal \c0.n5794_cascade_\ : std_logic;
signal \c0.n6015\ : std_logic;
signal \c0.n6072_cascade_\ : std_logic;
signal \c0.n6018\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal \c0.tx2.n6048_cascade_\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_1798_cascade_\ : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal \c0.tx2.n4779\ : std_logic;
signal \c0.tx2.n4780\ : std_logic;
signal \c0.tx2.n318\ : std_logic;
signal \c0.tx2.n4781\ : std_logic;
signal \c0.tx2.n317\ : std_logic;
signal \c0.tx2.n4782\ : std_logic;
signal \c0.tx2.n4783\ : std_logic;
signal \c0.tx2.n4784\ : std_logic;
signal \c0.tx2.n4785\ : std_logic;
signal \c0.tx2.n4786\ : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal n313_adj_1997 : std_logic;
signal \c0.n6135_cascade_\ : std_logic;
signal \c0.n5746_cascade_\ : std_logic;
signal \c0.n6153_cascade_\ : std_logic;
signal \c0.n5740_cascade_\ : std_logic;
signal \c0.n6129\ : std_logic;
signal \c0.n6063\ : std_logic;
signal \c0.n5776\ : std_logic;
signal \c0.n6099\ : std_logic;
signal \c0.tx2.n6006\ : std_logic;
signal \c0.n5375_cascade_\ : std_logic;
signal \c0.n5755\ : std_logic;
signal \c0.n6075_cascade_\ : std_logic;
signal \c0.n5773\ : std_logic;
signal \c0.n5454_cascade_\ : std_logic;
signal \c0.n27_cascade_\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.n52_cascade_\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.n32\ : std_logic;
signal \c0.n24_adj_1879_cascade_\ : std_logic;
signal \c0.n6102\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.tx2.n6045\ : std_logic;
signal \c0.data_in_frame_18_2\ : std_logic;
signal \c0.n6297_cascade_\ : std_logic;
signal \c0.n6300\ : std_logic;
signal \c0.data_in_frame_18_3\ : std_logic;
signal \c0.n6279_cascade_\ : std_logic;
signal \c0.n6282_cascade_\ : std_logic;
signal \c0.n6132\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal \c0.n6069\ : std_logic;
signal \c0.n6249_cascade_\ : std_logic;
signal \c0.n28\ : std_logic;
signal \c0.n3703_cascade_\ : std_logic;
signal \c0.n6117\ : std_logic;
signal \c0.n5536_cascade_\ : std_logic;
signal \c0.n5570_cascade_\ : std_logic;
signal \c0.n27_adj_1910\ : std_logic;
signal \c0.n3689_cascade_\ : std_logic;
signal \c0.tx2.n12\ : std_logic;
signal \c0.n3689\ : std_logic;
signal \c0.n3703\ : std_logic;
signal \c0.tx2.r_Bit_Index_2\ : std_logic;
signal \c0.tx2.n1136\ : std_logic;
signal \n4_adj_1973_cascade_\ : std_logic;
signal tx2_active : std_logic;
signal \c0.r_SM_Main_2_N_1770_0\ : std_logic;
signal tx2_o : std_logic;
signal tx2_enable : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal \r_SM_Main_1_adj_1993\ : std_logic;
signal \c0.tx2.r_SM_Main_2_N_1767_1_cascade_\ : std_logic;
signal \c0.tx2.n315\ : std_logic;
signal \c0.tx2.n5824\ : std_logic;
signal \c0.tx2.n5816\ : std_logic;
signal \c0.tx2.n314\ : std_logic;
signal \c0.tx2.n319\ : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal \c0.tx2.n316\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.n14_adj_1867\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \r_Clock_Count_8_adj_1994\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \c0.tx2.n31\ : std_logic;
signal \c0.tx2.n9\ : std_logic;
signal \c0.tx2.n5631_cascade_\ : std_logic;
signal \c0.tx2.n78\ : std_logic;
signal n4544 : std_logic;
signal \c0.n6159_cascade_\ : std_logic;
signal \c0.n5737\ : std_logic;
signal \c0.n5743\ : std_logic;
signal \c0.n6141\ : std_logic;
signal \c0.n6123_cascade_\ : std_logic;
signal \c0.n5752\ : std_logic;
signal data_in_14_7 : std_logic;
signal \c0.n24_adj_1877\ : std_logic;
signal \c0.data_in_frame_19_2\ : std_logic;
signal \c0.n5381\ : std_logic;
signal \c0.n5381_cascade_\ : std_logic;
signal data_in_13_7 : std_logic;
signal \c0.n2009\ : std_logic;
signal data_in_16_6 : std_logic;
signal \c0.n1942_cascade_\ : std_logic;
signal \c0.n18_adj_1938\ : std_logic;
signal \c0.n5578_cascade_\ : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n5488_cascade_\ : std_logic;
signal \c0.n36_cascade_\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.n12\ : std_logic;
signal \c0.n5488\ : std_logic;
signal \c0.n5489\ : std_logic;
signal \c0.n1886\ : std_logic;
signal \c0.n1942\ : std_logic;
signal \c0.n12_adj_1951\ : std_logic;
signal data_in_14_2 : std_logic;
signal \c0.n5536\ : std_logic;
signal \c0.n5586\ : std_logic;
signal \c0.data_in_frame_19_3\ : std_logic;
signal \c0.n22_adj_1876\ : std_logic;
signal \c0.data_in_field_49\ : std_logic;
signal \c0.n5991_cascade_\ : std_logic;
signal \c0.n6105\ : std_logic;
signal \c0.data_in_frame_18_5\ : std_logic;
signal \c0.n6225_cascade_\ : std_logic;
signal \c0.n6228_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal \c0.n6267_cascade_\ : std_logic;
signal \c0.n6270_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.n6081\ : std_logic;
signal \c0.n6084\ : std_logic;
signal \c0.n5695\ : std_logic;
signal \c0.n6234_cascade_\ : std_logic;
signal \c0.n1081\ : std_logic;
signal \c0.tx2.n1624\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal \c0.tx2.r_Bit_Index_1\ : std_logic;
signal \c0.tx2.n6003\ : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission_N_909\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \c0.n4735\ : std_logic;
signal \c0.n4736\ : std_logic;
signal \c0.n4737\ : std_logic;
signal \c0.n4738\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.n195\ : std_logic;
signal \c0.n2325\ : std_logic;
signal \r_SM_Main_2_adj_1992\ : std_logic;
signal \c0.tx2.n14\ : std_logic;
signal \c0.tx2.r_SM_Main_0\ : std_logic;
signal n2208 : std_logic;
signal n2339 : std_logic;
signal \r_Bit_Index_0_adj_1995\ : std_logic;
signal \c0.tx2.r_SM_Main_2_N_1767_1\ : std_logic;
signal \c0.tx2.n5847\ : std_logic;
signal \c0.rx.n3589\ : std_logic;
signal \c0.rx.n3589_cascade_\ : std_logic;
signal \c0.rx.n17_cascade_\ : std_logic;
signal \c0.rx.n5817\ : std_logic;
signal data_in_15_3 : std_logic;
signal \c0.data_in_field_59\ : std_logic;
signal \c0.data_in_field_123\ : std_logic;
signal data_in_7_3 : std_logic;
signal \c0.data_in_field_11\ : std_logic;
signal data_in_8_3 : std_logic;
signal \c0.data_in_field_67\ : std_logic;
signal data_in_10_3 : std_logic;
signal \c0.n5412_cascade_\ : std_logic;
signal \c0.n16_adj_1880\ : std_logic;
signal \c0.n22_adj_1881_cascade_\ : std_logic;
signal \c0.n24_adj_1884\ : std_logic;
signal \c0.data_in_field_81\ : std_logic;
signal \c0.n5551\ : std_logic;
signal \c0.n5551_cascade_\ : std_logic;
signal \c0.n1892\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.n19_cascade_\ : std_logic;
signal \c0.n5578\ : std_logic;
signal \c0.n6177_cascade_\ : std_logic;
signal \c0.n5728_cascade_\ : std_logic;
signal \c0.n16_adj_1873_cascade_\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n5725\ : std_logic;
signal \c0.n6165\ : std_logic;
signal \c0.n6168\ : std_logic;
signal \c0.n20_adj_1878\ : std_logic;
signal data_in_7_2 : std_logic;
signal \c0.data_in_field_58\ : std_logic;
signal \c0.data_in_frame_19_6\ : std_logic;
signal \c0.n6147_cascade_\ : std_logic;
signal \c0.n6150\ : std_logic;
signal \c0.data_in_frame_19_4\ : std_logic;
signal \c0.data_in_field_14\ : std_logic;
signal \c0.n6255_cascade_\ : std_logic;
signal \c0.n5692\ : std_logic;
signal \c0.data_in_field_119\ : std_logic;
signal \c0.n6273_cascade_\ : std_logic;
signal \c0.data_in_field_111\ : std_logic;
signal \c0.n5994\ : std_logic;
signal \c0.n5686_cascade_\ : std_logic;
signal \c0.n6261_cascade_\ : std_logic;
signal \c0.n6264\ : std_logic;
signal data_in_18_3 : std_logic;
signal \c0.data_in_field_104\ : std_logic;
signal \c0.n6021_cascade_\ : std_logic;
signal \c0.n5797\ : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal \c0.rx.n5860\ : std_logic;
signal \c0.rx.n4772\ : std_logic;
signal \c0.rx.n4773\ : std_logic;
signal \c0.rx.n5856\ : std_logic;
signal \c0.rx.n4774\ : std_logic;
signal \c0.rx.n4775\ : std_logic;
signal \c0.rx.n4776\ : std_logic;
signal \c0.rx.n4777\ : std_logic;
signal \c0.rx.n36\ : std_logic;
signal \c0.rx.n4778\ : std_logic;
signal \c0.rx.n5361\ : std_logic;
signal \c0.rx.n5858\ : std_logic;
signal \c0.rx.n5854\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.n8_cascade_\ : std_logic;
signal \c0.rx.n1724\ : std_logic;
signal \c0.rx.n1724_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n5855\ : std_logic;
signal \c0.rx.r_Clock_Count_0\ : std_logic;
signal \c0.rx.n5857\ : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal tx_enable : std_logic;
signal data_in_16_3 : std_logic;
signal rx_data_3 : std_logic;
signal data_in_18_1 : std_logic;
signal \c0.n6009_cascade_\ : std_logic;
signal \c0.n6012\ : std_logic;
signal \c0.data_in_field_15\ : std_logic;
signal \c0.data_in_field_8\ : std_logic;
signal \c0.n2039\ : std_logic;
signal \c0.n2039_cascade_\ : std_logic;
signal \c0.data_in_field_23\ : std_logic;
signal \c0.data_in_field_138\ : std_logic;
signal \c0.data_in_field_130\ : std_logic;
signal \c0.n6213\ : std_logic;
signal \c0.data_in_field_73\ : std_logic;
signal \c0.n14_adj_1957_cascade_\ : std_logic;
signal \c0.data_in_field_53\ : std_logic;
signal \c0.n22_adj_1903_cascade_\ : std_logic;
signal \c0.n18_adj_1904\ : std_logic;
signal \c0.n20_adj_1905\ : std_logic;
signal \c0.n5589_cascade_\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n5458\ : std_logic;
signal \c0.n1994\ : std_logic;
signal \c0.n5557\ : std_logic;
signal \c0.n17_cascade_\ : std_logic;
signal \c0.n5574\ : std_logic;
signal \c0.n5572\ : std_logic;
signal data_in_8_7 : std_logic;
signal data_in_17_1 : std_logic;
signal \c0.n1973\ : std_logic;
signal data_in_19_3 : std_logic;
signal \c0.n18_adj_1959_cascade_\ : std_logic;
signal \c0.n16\ : std_logic;
signal \c0.n20_adj_1870_cascade_\ : std_logic;
signal \c0.n5577\ : std_logic;
signal \c0.n2101_cascade_\ : std_logic;
signal \c0.n6_adj_1917_cascade_\ : std_logic;
signal \c0.data_in_field_68\ : std_logic;
signal \c0.n5512\ : std_logic;
signal \c0.n5512_cascade_\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.n2155\ : std_logic;
signal \c0.n2155_cascade_\ : std_logic;
signal \c0.n43\ : std_logic;
signal \c0.n2026\ : std_logic;
signal data_in_16_1 : std_logic;
signal \c0.n2080\ : std_logic;
signal \c0.n2012\ : std_logic;
signal data_in_19_6 : std_logic;
signal \c0.data_in_frame_19_0\ : std_logic;
signal \c0.data_in_field_17\ : std_logic;
signal \c0.n6093_cascade_\ : std_logic;
signal \c0.n5767\ : std_logic;
signal data_in_16_2 : std_logic;
signal data_in_18_6 : std_logic;
signal \c0.data_in_frame_18_6\ : std_logic;
signal \c0.data_in_frame_18_7\ : std_logic;
signal data_in_7_1 : std_logic;
signal \n1764_cascade_\ : std_logic;
signal rx_data_5 : std_logic;
signal rx_data_6 : std_logic;
signal \c0.rx.n5822\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal n4_adj_1980 : std_logic;
signal \n4_adj_1980_cascade_\ : std_logic;
signal rx_data_4 : std_logic;
signal \n2198_cascade_\ : std_logic;
signal \c0.rx.n359\ : std_logic;
signal \c0.rx.n5859\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.n5823\ : std_logic;
signal \c0.rx.n6294_cascade_\ : std_logic;
signal \r_SM_Main_2_adj_1989\ : std_logic;
signal \c0.rx.n75_cascade_\ : std_logic;
signal \c0.rx.n5815\ : std_logic;
signal data_in_1_3 : std_logic;
signal data_in_6_3 : std_logic;
signal data_in_12_3 : std_logic;
signal data_in_2_7 : std_logic;
signal \c0.data_in_field_131\ : std_logic;
signal data_in_1_1 : std_logic;
signal \c0.data_in_field_7\ : std_logic;
signal data_in_0_1 : std_logic;
signal \c0.n2104\ : std_logic;
signal \c0.n1835\ : std_logic;
signal \c0.n2104_cascade_\ : std_logic;
signal data_in_8_1 : std_logic;
signal \c0.n20_adj_1958\ : std_logic;
signal \c0.n31_adj_1896_cascade_\ : std_logic;
signal \c0.n41\ : std_logic;
signal \c0.data_in_field_6\ : std_logic;
signal \c0.n10_adj_1915\ : std_logic;
signal \c0.n1913\ : std_logic;
signal \c0.data_in_field_64\ : std_logic;
signal data_in_8_2 : std_logic;
signal data_in_5_3 : std_logic;
signal \c0.n6183\ : std_logic;
signal \c0.n2062_cascade_\ : std_logic;
signal \c0.n44\ : std_logic;
signal \c0.data_in_field_134\ : std_logic;
signal \c0.n5503\ : std_logic;
signal \c0.n2095\ : std_logic;
signal \c0.n16_adj_1871\ : std_logic;
signal data_in_11_3 : std_logic;
signal \c0.n2021\ : std_logic;
signal \c0.data_in_field_10\ : std_logic;
signal \c0.n2021_cascade_\ : std_logic;
signal \c0.data_in_field_41\ : std_logic;
signal \c0.n2074_cascade_\ : std_logic;
signal \c0.n2000\ : std_logic;
signal \c0.data_in_field_26\ : std_logic;
signal \c0.data_in_field_135\ : std_logic;
signal \c0.n1908\ : std_logic;
signal \c0.data_in_field_99\ : std_logic;
signal \c0.data_in_field_65\ : std_logic;
signal \c0.data_in_field_129\ : std_logic;
signal \c0.n5569\ : std_logic;
signal \c0.n5569_cascade_\ : std_logic;
signal \c0.data_in_field_114\ : std_logic;
signal \c0.n20_adj_1882\ : std_logic;
signal \c0.n5388\ : std_logic;
signal \c0.n5418\ : std_logic;
signal \c0.n5491\ : std_logic;
signal \c0.n44_adj_1894\ : std_logic;
signal \c0.data_in_field_112\ : std_logic;
signal \c0.data_in_field_30\ : std_logic;
signal \c0.data_in_field_125\ : std_logic;
signal \c0.n1889\ : std_logic;
signal \c0.data_in_field_76\ : std_logic;
signal \c0.data_in_frame_18_4\ : std_logic;
signal \c0.n6243_cascade_\ : std_logic;
signal \c0.n5698_cascade_\ : std_logic;
signal \c0.n6231\ : std_logic;
signal \c0.n6237\ : std_logic;
signal \c0.data_in_field_102\ : std_logic;
signal \c0.n5701\ : std_logic;
signal data_in_10_6 : std_logic;
signal \c0.data_in_field_86\ : std_logic;
signal data_in_10_1 : std_logic;
signal data_in_9_1 : std_logic;
signal data_in_12_6 : std_logic;
signal n1764 : std_logic;
signal rx_data_7 : std_logic;
signal data_in_15_6 : std_logic;
signal \r_SM_Main_0_adj_1991\ : std_logic;
signal \r_SM_Main_2_N_1824_2\ : std_logic;
signal \c0.rx.n6291\ : std_logic;
signal \c0.rx.n5633\ : std_logic;
signal n3636 : std_logic;
signal \c0.rx.n3850\ : std_logic;
signal \r_SM_Main_1_adj_1990\ : std_logic;
signal \c0.rx.n3850_cascade_\ : std_logic;
signal \c0.rx.n2259\ : std_logic;
signal \c0.rx.n2367\ : std_logic;
signal data_in_2_5 : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.n27_adj_1928\ : std_logic;
signal \c0.n28_adj_1926_cascade_\ : std_logic;
signal \c0.n25_adj_1929\ : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_1_0 : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_1_7 : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.n30_adj_1941\ : std_logic;
signal \c0.n4795\ : std_logic;
signal \c0.n26_adj_1940\ : std_logic;
signal \c0.n1729_cascade_\ : std_logic;
signal \c0.data_in_field_35\ : std_logic;
signal \c0.data_in_field_9\ : std_logic;
signal \c0.data_in_field_54\ : std_logic;
signal \c0.n5369_cascade_\ : std_logic;
signal data_in_0_3 : std_logic;
signal data_in_9_3 : std_logic;
signal \c0.data_in_field_3\ : std_logic;
signal \c0.n2125\ : std_logic;
signal \c0.data_in_field_27\ : std_logic;
signal \c0.n5469\ : std_logic;
signal \c0.data_in_field_83\ : std_logic;
signal \c0.n5454\ : std_logic;
signal \c0.n5469_cascade_\ : std_logic;
signal \c0.n6_adj_1923\ : std_logic;
signal \c0.n5548_cascade_\ : std_logic;
signal data_in_0_4 : std_logic;
signal data_in_7_5 : std_logic;
signal \c0.data_in_field_33\ : std_logic;
signal \c0.data_in_field_140\ : std_logic;
signal data_in_12_7 : std_logic;
signal \c0.data_in_field_126\ : std_logic;
signal \c0.data_in_field_118\ : std_logic;
signal \c0.data_in_field_51\ : std_logic;
signal data_in_16_5 : std_logic;
signal \c0.data_in_field_52\ : std_logic;
signal \c0.data_in_field_103\ : std_logic;
signal \c0.n2152\ : std_logic;
signal \c0.data_in_field_43\ : std_logic;
signal \c0.n2152_cascade_\ : std_logic;
signal \c0.n5397\ : std_logic;
signal data_in_11_6 : std_logic;
signal \c0.data_in_field_75\ : std_logic;
signal data_in_17_6 : std_logic;
signal \c0.data_in_field_142\ : std_logic;
signal \c0.tx2_transmit_N_1031_cascade_\ : std_logic;
signal \c0.data_in_field_29\ : std_logic;
signal \c0.n2030\ : std_logic;
signal \c0.n2030_cascade_\ : std_logic;
signal data_in_15_2 : std_logic;
signal \c0.data_in_field_22\ : std_logic;
signal \c0.n5436\ : std_logic;
signal \c0.n5436_cascade_\ : std_logic;
signal \c0.n5509\ : std_logic;
signal \c0.data_in_field_78\ : std_logic;
signal \c0.n5509_cascade_\ : std_logic;
signal \c0.data_in_field_92\ : std_logic;
signal \c0.data_in_field_36\ : std_logic;
signal \c0.data_in_field_82\ : std_logic;
signal \c0.n1948\ : std_logic;
signal data_in_15_1 : std_logic;
signal data_in_14_1 : std_logic;
signal \c0.data_in_field_127\ : std_logic;
signal n4 : std_logic;
signal data_in_13_1 : std_logic;
signal \c0.data_in_field_105\ : std_logic;
signal \c0.n18_adj_1887\ : std_logic;
signal \c0.n20_adj_1888\ : std_logic;
signal data_in_12_1 : std_logic;
signal \c0.data_in_field_97\ : std_logic;
signal \c0.data_in_frame_19_5\ : std_logic;
signal data_in_14_6 : std_logic;
signal data_in_19_7 : std_logic;
signal \c0.data_in_frame_19_7\ : std_logic;
signal data_in_19_5 : std_logic;
signal data_in_14_0 : std_logic;
signal data_in_13_0 : std_logic;
signal data_in_18_4 : std_logic;
signal \c0.tx.n40_cascade_\ : std_logic;
signal n1760 : std_logic;
signal \c0.tx.n2247\ : std_logic;
signal \c0.tx.n2356\ : std_logic;
signal \c0.rx.r_Bit_Index_2\ : std_logic;
signal \c0.rx.r_Bit_Index_1\ : std_logic;
signal \c0.rx.n1706\ : std_logic;
signal \n1757_cascade_\ : std_logic;
signal rx_data_0 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n1757 : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_0_5 : std_logic;
signal \c0.n22_adj_1924\ : std_logic;
signal \c0.data_in_field_141\ : std_logic;
signal \c0.n5527\ : std_logic;
signal \c0.n5394_cascade_\ : std_logic;
signal \c0.n1926\ : std_logic;
signal \c0.n19_adj_1889\ : std_logic;
signal \c0.n22_adj_1886\ : std_logic;
signal \c0.n5590\ : std_logic;
signal \c0.n40_cascade_\ : std_logic;
signal \c0.n45_adj_1892\ : std_logic;
signal \c0.data_in_field_132\ : std_logic;
signal \c0.n1969\ : std_logic;
signal \c0.n5403\ : std_logic;
signal data_in_19_4 : std_logic;
signal \c0.data_in_field_115\ : std_logic;
signal \c0.n1855_cascade_\ : std_logic;
signal \c0.n1917\ : std_logic;
signal \c0.data_in_field_34\ : std_logic;
signal \c0.n2092\ : std_logic;
signal data_in_17_3 : std_logic;
signal data_in_2_3 : std_logic;
signal data_in_6_7 : std_logic;
signal data_in_6_5 : std_logic;
signal \c0.n25_adj_1948\ : std_logic;
signal \c0.data_in_field_94\ : std_logic;
signal \c0.data_in_field_66\ : std_logic;
signal \c0.data_in_field_79\ : std_logic;
signal \c0.n5545\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.data_in_field_95\ : std_logic;
signal \c0.data_in_field_96\ : std_logic;
signal data_in_15_5 : std_logic;
signal \c0.n6414\ : std_logic;
signal \c0.n5563\ : std_logic;
signal data_in_11_1 : std_logic;
signal \c0.data_in_field_45\ : std_logic;
signal \c0.n2065\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n2149_cascade_\ : std_logic;
signal \c0.n21\ : std_logic;
signal data_in_3_2 : std_logic;
signal \c0.n1955\ : std_logic;
signal data_in_4_2 : std_logic;
signal data_in_18_5 : std_logic;
signal data_in_17_5 : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \c0.n4754\ : std_logic;
signal \c0.n4755\ : std_logic;
signal \c0.n4756\ : std_logic;
signal \c0.n4757\ : std_logic;
signal \c0.n4758\ : std_logic;
signal \c0.n4759\ : std_logic;
signal \c0.n4760\ : std_logic;
signal \c0.n4761\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \c0.n4762\ : std_logic;
signal \c0.n4763\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.data_in_field_116\ : std_logic;
signal \c0.data_in_field_124\ : std_logic;
signal \c0.n6171_cascade_\ : std_logic;
signal \c0.n5731\ : std_logic;
signal \c0.data_in_field_4\ : std_logic;
signal \c0.data_in_field_12\ : std_logic;
signal \c0.n5722\ : std_logic;
signal \c0.tx.n3631_cascade_\ : std_logic;
signal \c0.data_in_field_20\ : std_logic;
signal \c0.n6189\ : std_logic;
signal \c0.tx.n5812_cascade_\ : std_logic;
signal \c0.tx.n14_cascade_\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \c0.tx.n4764\ : std_logic;
signal \c0.tx.n4765\ : std_logic;
signal \c0.tx.n4766\ : std_logic;
signal \c0.tx.n4767\ : std_logic;
signal \c0.tx.n4768\ : std_logic;
signal \c0.tx.n4769\ : std_logic;
signal \c0.tx.n4770\ : std_logic;
signal \c0.tx.n4771\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \c0.tx.n5885\ : std_logic;
signal \c0.tx.n15\ : std_logic;
signal \c0.tx.n5884\ : std_logic;
signal data_in_4_3 : std_logic;
signal data_in_3_3 : std_logic;
signal data_in_2_2 : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.data_in_field_80\ : std_logic;
signal \c0.n42_cascade_\ : std_logic;
signal \c0.n48\ : std_logic;
signal data_in_19_0 : std_logic;
signal data_in_15_7 : std_logic;
signal data_in_16_7 : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.n22_adj_1890\ : std_logic;
signal \c0.data_in_field_61\ : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_0_0 : std_logic;
signal \c0.data_in_field_0\ : std_logic;
signal \c0.data_in_field_117\ : std_logic;
signal \c0.n1855\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.n12_adj_1898_cascade_\ : std_logic;
signal \c0.n47_adj_1897\ : std_logic;
signal \c0.n48_adj_1895\ : std_logic;
signal \c0.n5567_cascade_\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n6219\ : std_logic;
signal \c0.data_in_field_5\ : std_logic;
signal \c0.n1979\ : std_logic;
signal \c0.n1958\ : std_logic;
signal \c0.n2056\ : std_logic;
signal \c0.n5506\ : std_logic;
signal \c0.n5575\ : std_logic;
signal \c0.n5506_cascade_\ : std_logic;
signal \c0.n5539\ : std_logic;
signal \c0.n1779\ : std_logic;
signal \c0.data_in_field_60\ : std_logic;
signal \c0.n5500\ : std_logic;
signal \c0.data_in_field_19\ : std_logic;
signal \c0.data_in_field_139\ : std_logic;
signal data_in_5_5 : std_logic;
signal data_in_6_1 : std_logic;
signal data_in_5_1 : std_logic;
signal data_in_4_1 : std_logic;
signal data_in_18_7 : std_logic;
signal data_in_17_7 : std_logic;
signal \c0.n6_adj_1918\ : std_logic;
signal data_in_1_4 : std_logic;
signal \c0.data_in_field_18\ : std_logic;
signal \c0.n5372\ : std_logic;
signal \c0.n2043_cascade_\ : std_logic;
signal \c0.data_in_field_107\ : std_logic;
signal data_in_13_6 : std_logic;
signal \c0.n5443\ : std_logic;
signal \c0.data_in_field_89\ : std_logic;
signal \c0.data_in_field_90\ : std_logic;
signal data_in_7_7 : std_logic;
signal \c0.data_in_field_37\ : std_logic;
signal \c0.data_in_frame_18_0\ : std_logic;
signal \c0.n2077\ : std_logic;
signal \c0.n5707\ : std_logic;
signal \c0.n5710\ : std_logic;
signal \c0.n6198\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal data_in_5_0 : std_logic;
signal data_in_4_0 : std_logic;
signal data_in_8_4 : std_logic;
signal data_in_7_4 : std_logic;
signal data_in_6_4 : std_logic;
signal data_in_5_6 : std_logic;
signal \n5646_cascade_\ : std_logic;
signal n5645 : std_logic;
signal \LED_c\ : std_logic;
signal \c0.data_in_field_110\ : std_logic;
signal \c0.n5533\ : std_logic;
signal data_out_18_6 : std_logic;
signal \c0.n17_adj_1913_cascade_\ : std_logic;
signal \c0.tx.n5883\ : std_logic;
signal \c0.n1253_cascade_\ : std_logic;
signal \c0.n5830\ : std_logic;
signal \c0.n22_adj_1914_cascade_\ : std_logic;
signal \tx_data_6_N_keep\ : std_logic;
signal \c0.n5827\ : std_logic;
signal \c0.n1253\ : std_logic;
signal \tx_data_7_N_keep\ : std_logic;
signal data_out_18_0 : std_logic;
signal data_out_19_0 : std_logic;
signal \c0.n1198\ : std_logic;
signal \c0.n5810_cascade_\ : std_logic;
signal \c0.tx_data_0_N\ : std_logic;
signal \c0.tx.n14_adj_1869_cascade_\ : std_logic;
signal \c0.tx.r_SM_Main_2_N_1767_1_cascade_\ : std_logic;
signal \c0.tx.n5821\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal n315 : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal n317 : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.tx.n10_adj_1868\ : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal \c0.tx.n5627\ : std_logic;
signal \n11_adj_1979_cascade_\ : std_logic;
signal \c0.tx.n5629\ : std_logic;
signal \c0.tx.n3120\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n3120_cascade_\ : std_logic;
signal n313 : std_logic;
signal \n782_cascade_\ : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal data_in_9_2 : std_logic;
signal \c0.n5384\ : std_logic;
signal \c0.n5476\ : std_logic;
signal \c0.n5427\ : std_logic;
signal \c0.n5521\ : std_logic;
signal \c0.n24_adj_1885\ : std_logic;
signal \c0.n1866\ : std_logic;
signal \c0.data_in_field_113\ : std_logic;
signal \c0.data_in_field_57\ : std_logic;
signal \c0.n10_cascade_\ : std_logic;
signal \c0.n5466\ : std_logic;
signal \c0.n5519\ : std_logic;
signal data_in_7_6 : std_logic;
signal data_in_6_6 : std_logic;
signal data_in_18_0 : std_logic;
signal \c0.n5548\ : std_logic;
signal \c0.n5497\ : std_logic;
signal \c0.n5515\ : std_logic;
signal \c0.data_in_field_44\ : std_logic;
signal \c0.data_in_field_100\ : std_logic;
signal \c0.data_in_field_50\ : std_logic;
signal \c0.n2053\ : std_logic;
signal \c0.n2101\ : std_logic;
signal \c0.n2134\ : std_logic;
signal \c0.n31_adj_1900_cascade_\ : std_logic;
signal \c0.n35\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n5582\ : std_logic;
signal \c0.n13_adj_1899\ : std_logic;
signal \c0.n17_adj_1902\ : std_logic;
signal \c0.n25_adj_1907\ : std_logic;
signal \c0.n4_adj_1920\ : std_logic;
signal \c0.data_in_field_122\ : std_logic;
signal \c0.n5593\ : std_logic;
signal \c0.data_in_field_62\ : std_logic;
signal \c0.n5593_cascade_\ : std_logic;
signal \c0.n5430\ : std_logic;
signal \c0.n33\ : std_logic;
signal \c0.n5430_cascade_\ : std_logic;
signal \c0.n28_adj_1955\ : std_logic;
signal \c0.n37\ : std_logic;
signal data_in_1_5 : std_logic;
signal \c0.data_in_field_13\ : std_logic;
signal \c0.n6_adj_1939\ : std_logic;
signal data_in_12_4 : std_logic;
signal data_in_11_4 : std_logic;
signal \c0.n2089\ : std_logic;
signal \c0.n2074\ : std_logic;
signal \c0.n5581\ : std_logic;
signal \c0.data_in_field_120\ : std_logic;
signal \c0.n2107\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.n6201\ : std_logic;
signal \c0.data_in_field_101\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n5716_cascade_\ : std_logic;
signal \c0.n6195\ : std_logic;
signal \c0.data_in_field_85\ : std_logic;
signal \c0.data_in_field_93\ : std_logic;
signal \c0.data_in_field_77\ : std_logic;
signal \c0.n6207_cascade_\ : std_logic;
signal \c0.data_in_field_69\ : std_logic;
signal \c0.n5713\ : std_logic;
signal data_in_19_2 : std_logic;
signal data_in_9_0 : std_logic;
signal \c0.data_in_field_42\ : std_logic;
signal \c0.data_in_field_72\ : std_logic;
signal data_in_12_0 : std_logic;
signal data_in_18_2 : std_logic;
signal data_in_17_2 : std_logic;
signal data_in_6_2 : std_logic;
signal data_in_5_2 : std_logic;
signal data_in_4_5 : std_logic;
signal data_in_11_7 : std_logic;
signal \n5448_cascade_\ : std_logic;
signal n4_adj_1975 : std_logic;
signal data_out_19_4 : std_logic;
signal data_out_18_4 : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal \c0.n18_adj_1919\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.n20_adj_1922_cascade_\ : std_logic;
signal \c0.n16_adj_1921\ : std_logic;
signal \n4334_cascade_\ : std_logic;
signal n1991 : std_logic;
signal data_out_19_7 : std_logic;
signal \c0.n17_adj_1950\ : std_logic;
signal n4_adj_1982 : std_logic;
signal \c0.n17_adj_1908\ : std_logic;
signal data_out_18_7 : std_logic;
signal \c0.n1508\ : std_logic;
signal data_out_19_2 : std_logic;
signal \c0.n1508_cascade_\ : std_logic;
signal \c0.n5840\ : std_logic;
signal \c0.n6309_cascade_\ : std_logic;
signal data_out_18_2 : std_logic;
signal \c0.n1249\ : std_logic;
signal \tx_data_4_N_keep\ : std_logic;
signal \c0.tx.n3644\ : std_logic;
signal n11_adj_1979 : std_logic;
signal \n5818_cascade_\ : std_logic;
signal n4155 : std_logic;
signal n318 : std_logic;
signal \r_Clock_Count_3\ : std_logic;
signal n321 : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal data_out_18_5 : std_logic;
signal n782 : std_logic;
signal n320 : std_logic;
signal \r_Clock_Count_1\ : std_logic;
signal rx_data_1 : std_logic;
signal data_in_14_3 : std_logic;
signal data_in_13_3 : std_logic;
signal \c0.data_in_field_55\ : std_logic;
signal \c0.data_in_field_63\ : std_logic;
signal data_in_14_4 : std_logic;
signal \c0.data_in_field_48\ : std_logic;
signal \c0.data_in_field_32\ : std_logic;
signal \c0.data_in_field_40\ : std_logic;
signal \c0.n6033_cascade_\ : std_logic;
signal \c0.n5791\ : std_logic;
signal \c0.n1814\ : std_logic;
signal data_in_19_1 : std_logic;
signal \c0.n2143\ : std_logic;
signal \c0.n1814_cascade_\ : std_logic;
signal \c0.data_in_field_109\ : std_logic;
signal \c0.n32_adj_1901\ : std_logic;
signal data_in_8_5 : std_logic;
signal data_in_17_4 : std_logic;
signal data_in_5_4 : std_logic;
signal \c0.n5560\ : std_logic;
signal \c0.data_in_field_106\ : std_logic;
signal \c0.data_in_field_2\ : std_logic;
signal \c0.n5560_cascade_\ : std_logic;
signal \c0.n34\ : std_logic;
signal data_in_5_7 : std_logic;
signal \c0.data_in_field_133\ : std_logic;
signal \c0.data_in_field_21\ : std_logic;
signal \c0.data_in_field_143\ : std_logic;
signal \c0.n5378\ : std_logic;
signal data_in_11_5 : std_logic;
signal data_in_2_0 : std_logic;
signal data_in_13_2 : std_logic;
signal \c0.data_in_field_88\ : std_logic;
signal \c0.data_in_field_98\ : std_logic;
signal \c0.data_in_field_28\ : std_logic;
signal \c0.data_in_field_121\ : std_logic;
signal \c0.n23_adj_1935\ : std_logic;
signal \c0.data_in_field_87\ : std_logic;
signal \c0.data_in_field_128\ : std_logic;
signal \c0.n2068\ : std_logic;
signal \c0.data_in_field_46\ : std_logic;
signal \c0.n1965_cascade_\ : std_logic;
signal \c0.data_in_field_91\ : std_logic;
signal \c0.n24_adj_1930\ : std_logic;
signal data_in_3_5 : std_logic;
signal data_in_3_0 : std_logic;
signal data_in_2_6 : std_logic;
signal \c0.n28_adj_1925\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.data_in_field_24\ : std_logic;
signal \c0.n6039\ : std_logic;
signal \n5_cascade_\ : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.tx.r_SM_Main_2_N_1767_1\ : std_logic;
signal \c0.tx.n2177\ : std_logic;
signal \n4333_cascade_\ : std_logic;
signal \c0.n81_adj_1872_cascade_\ : std_logic;
signal tx_active : std_logic;
signal \c0.tx_transmit\ : std_logic;
signal n135 : std_logic;
signal \n4_adj_1986_cascade_\ : std_logic;
signal data_out_19_6 : std_logic;
signal data_out_19_5 : std_logic;
signal n5440 : std_logic;
signal \c0.n9\ : std_logic;
signal n8_adj_1987 : std_logic;
signal n5400 : std_logic;
signal \tx_data_2_N_keep\ : std_logic;
signal n5364 : std_logic;
signal n5482 : std_logic;
signal n1768 : std_logic;
signal \n5364_cascade_\ : std_logic;
signal n5871 : std_logic;
signal \c0.n6312\ : std_logic;
signal \tx_data_3_N_keep\ : std_logic;
signal \c0.n5853\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \c0.tx.r_Bit_Index_0\ : std_logic;
signal \c0.tx.r_Tx_Data_0\ : std_logic;
signal \c0.tx.n6051_cascade_\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.tx.r_Bit_Index_2\ : std_logic;
signal \c0.tx.n6054\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \c0.tx.o_Tx_Serial_N_1798_cascade_\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.tx.n12_cascade_\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal tx_o : std_logic;
signal data_in_10_5 : std_logic;
signal data_in_9_5 : std_logic;
signal data_in_6_0 : std_logic;
signal data_in_10_4 : std_logic;
signal data_in_9_4 : std_logic;
signal data_in_16_4 : std_logic;
signal data_in_15_4 : std_logic;
signal data_in_13_4 : std_logic;
signal \c0.data_in_field_108\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.data_in_field_47\ : std_logic;
signal \c0.n5997\ : std_logic;
signal \c0.n6000\ : std_logic;
signal \c0.data_in_field_84\ : std_logic;
signal \c0.data_in_field_70\ : std_logic;
signal \c0.data_in_field_56\ : std_logic;
signal \c0.n5494\ : std_logic;
signal \c0.n5554\ : std_logic;
signal \c0.n5524\ : std_logic;
signal \c0.n5494_cascade_\ : std_logic;
signal \c0.n5391\ : std_logic;
signal \c0.n26_adj_1927\ : std_logic;
signal data_in_8_0 : std_logic;
signal data_in_7_0 : std_logic;
signal \c0.data_in_field_74\ : std_logic;
signal \c0.data_in_field_1\ : std_logic;
signal \c0.data_in_field_16\ : std_logic;
signal \c0.n25_adj_1931\ : std_logic;
signal \c0.data_in_field_137\ : std_logic;
signal \c0.data_in_field_25\ : std_logic;
signal \c0.data_in_field_71\ : std_logic;
signal \c0.n5542\ : std_logic;
signal data_in_17_0 : std_logic;
signal data_in_10_2 : std_logic;
signal data_in_4_6 : std_logic;
signal \c0.data_in_field_38\ : std_logic;
signal \c0.data_in_field_136\ : std_logic;
signal \c0.data_in_field_31\ : std_logic;
signal \c0.n2113\ : std_logic;
signal data_in_11_0 : std_logic;
signal data_in_10_0 : std_logic;
signal \c0.FRAME_MATCHER_wait_for_transmission\ : std_logic;
signal \c0.n1729\ : std_logic;
signal data_in_4_7 : std_logic;
signal \c0.data_in_field_39\ : std_logic;
signal data_in_10_7 : std_logic;
signal data_in_9_7 : std_logic;
signal data_in_14_5 : std_logic;
signal data_in_12_2 : std_logic;
signal data_in_11_2 : std_logic;
signal data_in_4_4 : std_logic;
signal data_in_9_6 : std_logic;
signal data_in_8_6 : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.n50_adj_1875\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \c0.n4703\ : std_logic;
signal \c0.n4704\ : std_logic;
signal \c0.n4705\ : std_logic;
signal \c0.n4706\ : std_logic;
signal \c0.byte_transmit_counter_5\ : std_logic;
signal \c0.tx_transmit_N_568_5\ : std_logic;
signal \c0.n4707\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.tx_transmit_N_568_6\ : std_logic;
signal \c0.n4708\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n4709\ : std_logic;
signal \c0.tx_transmit_N_568_7\ : std_logic;
signal \c0.tx_transmit_N_568_3\ : std_logic;
signal \c0.n95\ : std_logic;
signal \c0.n95_cascade_\ : std_logic;
signal \c0.n106\ : std_logic;
signal n4_adj_1981 : std_logic;
signal n7_adj_1988 : std_logic;
signal \c0.n15\ : std_logic;
signal \c0.n81_adj_1872\ : std_logic;
signal \c0.tx_transmit_N_568_4\ : std_logic;
signal \c0.tx_transmit_N_568_2\ : std_logic;
signal \c0.n5833\ : std_logic;
signal \c0.n31_adj_1912\ : std_logic;
signal \c0.n989\ : std_logic;
signal \c0.n9_adj_1906_cascade_\ : std_logic;
signal \c0.n15_adj_1909\ : std_logic;
signal data_out_10_4 : std_logic;
signal \c0.n2293\ : std_logic;
signal n4_adj_1996 : std_logic;
signal n1519 : std_logic;
signal \tx_data_5_N_keep\ : std_logic;
signal n5421 : std_logic;
signal data_out_18_1 : std_logic;
signal data_out_19_3 : std_logic;
signal \c0.n5837\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.tx.r_Bit_Index_1\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.tx.n6285\ : std_logic;
signal \c0.tx.n6288\ : std_logic;
signal n5415 : std_logic;
signal \c0.n1251\ : std_logic;
signal \c0.n5845\ : std_logic;
signal \c0.byte_transmit_counter_4\ : std_logic;
signal \tx_data_1_N_keep\ : std_logic;
signal data_out_11_7 : std_logic;
signal data_in_13_5 : std_logic;
signal data_in_12_5 : std_logic;
signal data_out_10_5 : std_logic;
signal \c0.n9_adj_1911\ : std_logic;
signal data_out_10_0 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.byte_transmit_counter_3\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.n9_adj_1891_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n15_adj_1893\ : std_logic;
signal data_out_11_5 : std_logic;
signal data_out_10_6 : std_logic;
signal n4_adj_1976 : std_logic;
signal n26 : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal n25 : std_logic;
signal n4710 : std_logic;
signal n24 : std_logic;
signal n4711 : std_logic;
signal n23 : std_logic;
signal n4712 : std_logic;
signal n22 : std_logic;
signal n4713 : std_logic;
signal n21 : std_logic;
signal n4714 : std_logic;
signal n20 : std_logic;
signal n4715 : std_logic;
signal n19 : std_logic;
signal n4716 : std_logic;
signal n4717 : std_logic;
signal n18 : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal n17 : std_logic;
signal n4718 : std_logic;
signal n16 : std_logic;
signal n4719 : std_logic;
signal n15 : std_logic;
signal n4720 : std_logic;
signal n14 : std_logic;
signal n4721 : std_logic;
signal n13 : std_logic;
signal n4722 : std_logic;
signal n12 : std_logic;
signal n4723 : std_logic;
signal n11 : std_logic;
signal n4724 : std_logic;
signal n4725 : std_logic;
signal n10 : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal n9 : std_logic;
signal n4726 : std_logic;
signal n8 : std_logic;
signal n4727 : std_logic;
signal n7 : std_logic;
signal n4728 : std_logic;
signal n6 : std_logic;
signal n4729 : std_logic;
signal blink_counter_21 : std_logic;
signal n4730 : std_logic;
signal blink_counter_22 : std_logic;
signal n4731 : std_logic;
signal blink_counter_23 : std_logic;
signal n4732 : std_logic;
signal n4733 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal n4734 : std_logic;
signal blink_counter_25 : std_logic;
signal data_out_10_2 : std_logic;
signal data_out_11_6 : std_logic;
signal rx_data_ready : std_logic;
signal data_in_16_0 : std_logic;
signal data_in_15_0 : std_logic;
signal \c0.n5409\ : std_logic;
signal data_out_11_1 : std_logic;
signal \c0.n5409_cascade_\ : std_logic;
signal data_out_11_4 : std_logic;
signal n4_adj_1978 : std_logic;
signal n4_adj_1983 : std_logic;
signal data_out_11_2 : std_logic;
signal n21_adj_1977 : std_logic;
signal n4333 : std_logic;
signal data_out_10_1 : std_logic;
signal data_out_10_3 : std_logic;
signal n5424 : std_logic;
signal data_out_11_0 : std_logic;
signal data_out_10_7 : std_logic;
signal n5479 : std_logic;
signal data_out_11_3 : std_logic;
signal n8_adj_1984 : std_logic;
signal \n7_adj_1985_cascade_\ : std_logic;
signal data_out_19_1 : std_logic;
signal data_0 : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal data_1 : std_logic;
signal \c0.n4739\ : std_logic;
signal data_2 : std_logic;
signal \c0.n4740\ : std_logic;
signal data_3 : std_logic;
signal \c0.n4741\ : std_logic;
signal data_4 : std_logic;
signal \c0.n4742\ : std_logic;
signal data_5 : std_logic;
signal \c0.n4743\ : std_logic;
signal data_6 : std_logic;
signal \c0.n4744\ : std_logic;
signal data_7 : std_logic;
signal \c0.n4745\ : std_logic;
signal \c0.n4746\ : std_logic;
signal data_8 : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal data_9 : std_logic;
signal \c0.n4747\ : std_logic;
signal data_10 : std_logic;
signal \c0.n4748\ : std_logic;
signal data_11 : std_logic;
signal \c0.n4749\ : std_logic;
signal data_12 : std_logic;
signal \c0.n4750\ : std_logic;
signal data_13 : std_logic;
signal \c0.n4751\ : std_logic;
signal data_14 : std_logic;
signal \c0.n4752\ : std_logic;
signal \c0.n4753\ : std_logic;
signal data_15 : std_logic;
signal n1579 : std_logic;
signal n5433 : std_logic;
signal n4334 : std_logic;
signal data_out_18_3 : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37951\,
            DIN => \N__37950\,
            DOUT => \N__37949\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37951\,
            PADOUT => \N__37950\,
            PADIN => \N__37949\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__23712\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37942\,
            DIN => \N__37941\,
            DOUT => \N__37940\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37942\,
            PADOUT => \N__37941\,
            PADIN => \N__37940\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37933\,
            DIN => \N__37932\,
            DOUT => \N__37931\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37933\,
            PADOUT => \N__37932\,
            PADIN => \N__37931\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__37589\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37924\,
            DIN => \N__37923\,
            DOUT => \N__37922\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37924\,
            PADOUT => \N__37923\,
            PADIN => \N__37922\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12705\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__12675\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__37915\,
            DIN => \N__37914\,
            DOUT => \N__37913\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37915\,
            PADOUT => \N__37914\,
            PADIN => \N__37913\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__28890\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15213\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37906\,
            DIN => \N__37905\,
            DOUT => \N__37904\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__37906\,
            PADOUT => \N__37905\,
            PADIN => \N__37904\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__9581\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37881\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__37881\,
            I => \N__37877\
        );

    \I__9579\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37874\
        );

    \I__9578\ : Odrv12
    port map (
            O => \N__37877\,
            I => data_11
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__37874\,
            I => data_11
        );

    \I__9576\ : InMux
    port map (
            O => \N__37869\,
            I => \c0.n4749\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__37866\,
            I => \N__37863\
        );

    \I__9574\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37860\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__37860\,
            I => \N__37857\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__37857\,
            I => \N__37853\
        );

    \I__9571\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37850\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__37853\,
            I => data_12
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__37850\,
            I => data_12
        );

    \I__9568\ : InMux
    port map (
            O => \N__37845\,
            I => \c0.n4750\
        );

    \I__9567\ : CascadeMux
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__9566\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__37833\,
            I => \N__37829\
        );

    \I__9563\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37826\
        );

    \I__9562\ : Odrv4
    port map (
            O => \N__37829\,
            I => data_13
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__37826\,
            I => data_13
        );

    \I__9560\ : InMux
    port map (
            O => \N__37821\,
            I => \c0.n4751\
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__9558\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37812\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__37812\,
            I => \N__37809\
        );

    \I__9556\ : Span4Mux_v
    port map (
            O => \N__37809\,
            I => \N__37805\
        );

    \I__9555\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37802\
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__37805\,
            I => data_14
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__37802\,
            I => data_14
        );

    \I__9552\ : InMux
    port map (
            O => \N__37797\,
            I => \c0.n4752\
        );

    \I__9551\ : InMux
    port map (
            O => \N__37794\,
            I => \c0.n4753\
        );

    \I__9550\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37787\
        );

    \I__9549\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37784\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__37787\,
            I => \N__37781\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__37784\,
            I => data_15
        );

    \I__9546\ : Odrv12
    port map (
            O => \N__37781\,
            I => data_15
        );

    \I__9545\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37773\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__9543\ : Span4Mux_v
    port map (
            O => \N__37770\,
            I => \N__37767\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__37767\,
            I => n1579
        );

    \I__9541\ : CascadeMux
    port map (
            O => \N__37764\,
            I => \N__37761\
        );

    \I__9540\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37758\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__37758\,
            I => \N__37754\
        );

    \I__9538\ : CascadeMux
    port map (
            O => \N__37757\,
            I => \N__37751\
        );

    \I__9537\ : Span4Mux_v
    port map (
            O => \N__37754\,
            I => \N__37748\
        );

    \I__9536\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37745\
        );

    \I__9535\ : Span4Mux_h
    port map (
            O => \N__37748\,
            I => \N__37740\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37740\
        );

    \I__9533\ : Odrv4
    port map (
            O => \N__37740\,
            I => n5433
        );

    \I__9532\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37731\
        );

    \I__9531\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37728\
        );

    \I__9530\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37721\
        );

    \I__9529\ : InMux
    port map (
            O => \N__37734\,
            I => \N__37721\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__37731\,
            I => \N__37718\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37712\
        );

    \I__9526\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37709\
        );

    \I__9525\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37699\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37696\
        );

    \I__9523\ : Span4Mux_v
    port map (
            O => \N__37718\,
            I => \N__37693\
        );

    \I__9522\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37686\
        );

    \I__9521\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37686\
        );

    \I__9520\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37686\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__37712\,
            I => \N__37681\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__37709\,
            I => \N__37681\
        );

    \I__9517\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37676\
        );

    \I__9516\ : InMux
    port map (
            O => \N__37707\,
            I => \N__37676\
        );

    \I__9515\ : InMux
    port map (
            O => \N__37706\,
            I => \N__37673\
        );

    \I__9514\ : InMux
    port map (
            O => \N__37705\,
            I => \N__37666\
        );

    \I__9513\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37666\
        );

    \I__9512\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37666\
        );

    \I__9511\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37663\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37658\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__37696\,
            I => \N__37658\
        );

    \I__9508\ : Odrv4
    port map (
            O => \N__37693\,
            I => n4334
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__37686\,
            I => n4334
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__37681\,
            I => n4334
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__37676\,
            I => n4334
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__37673\,
            I => n4334
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__37666\,
            I => n4334
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__37663\,
            I => n4334
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__37658\,
            I => n4334
        );

    \I__9500\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37638\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__37638\,
            I => \N__37634\
        );

    \I__9498\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37631\
        );

    \I__9497\ : Span4Mux_h
    port map (
            O => \N__37634\,
            I => \N__37628\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__37631\,
            I => data_out_18_3
        );

    \I__9495\ : Odrv4
    port map (
            O => \N__37628\,
            I => data_out_18_3
        );

    \I__9494\ : ClkMux
    port map (
            O => \N__37623\,
            I => \N__37137\
        );

    \I__9493\ : ClkMux
    port map (
            O => \N__37622\,
            I => \N__37137\
        );

    \I__9492\ : ClkMux
    port map (
            O => \N__37621\,
            I => \N__37137\
        );

    \I__9491\ : ClkMux
    port map (
            O => \N__37620\,
            I => \N__37137\
        );

    \I__9490\ : ClkMux
    port map (
            O => \N__37619\,
            I => \N__37137\
        );

    \I__9489\ : ClkMux
    port map (
            O => \N__37618\,
            I => \N__37137\
        );

    \I__9488\ : ClkMux
    port map (
            O => \N__37617\,
            I => \N__37137\
        );

    \I__9487\ : ClkMux
    port map (
            O => \N__37616\,
            I => \N__37137\
        );

    \I__9486\ : ClkMux
    port map (
            O => \N__37615\,
            I => \N__37137\
        );

    \I__9485\ : ClkMux
    port map (
            O => \N__37614\,
            I => \N__37137\
        );

    \I__9484\ : ClkMux
    port map (
            O => \N__37613\,
            I => \N__37137\
        );

    \I__9483\ : ClkMux
    port map (
            O => \N__37612\,
            I => \N__37137\
        );

    \I__9482\ : ClkMux
    port map (
            O => \N__37611\,
            I => \N__37137\
        );

    \I__9481\ : ClkMux
    port map (
            O => \N__37610\,
            I => \N__37137\
        );

    \I__9480\ : ClkMux
    port map (
            O => \N__37609\,
            I => \N__37137\
        );

    \I__9479\ : ClkMux
    port map (
            O => \N__37608\,
            I => \N__37137\
        );

    \I__9478\ : ClkMux
    port map (
            O => \N__37607\,
            I => \N__37137\
        );

    \I__9477\ : ClkMux
    port map (
            O => \N__37606\,
            I => \N__37137\
        );

    \I__9476\ : ClkMux
    port map (
            O => \N__37605\,
            I => \N__37137\
        );

    \I__9475\ : ClkMux
    port map (
            O => \N__37604\,
            I => \N__37137\
        );

    \I__9474\ : ClkMux
    port map (
            O => \N__37603\,
            I => \N__37137\
        );

    \I__9473\ : ClkMux
    port map (
            O => \N__37602\,
            I => \N__37137\
        );

    \I__9472\ : ClkMux
    port map (
            O => \N__37601\,
            I => \N__37137\
        );

    \I__9471\ : ClkMux
    port map (
            O => \N__37600\,
            I => \N__37137\
        );

    \I__9470\ : ClkMux
    port map (
            O => \N__37599\,
            I => \N__37137\
        );

    \I__9469\ : ClkMux
    port map (
            O => \N__37598\,
            I => \N__37137\
        );

    \I__9468\ : ClkMux
    port map (
            O => \N__37597\,
            I => \N__37137\
        );

    \I__9467\ : ClkMux
    port map (
            O => \N__37596\,
            I => \N__37137\
        );

    \I__9466\ : ClkMux
    port map (
            O => \N__37595\,
            I => \N__37137\
        );

    \I__9465\ : ClkMux
    port map (
            O => \N__37594\,
            I => \N__37137\
        );

    \I__9464\ : ClkMux
    port map (
            O => \N__37593\,
            I => \N__37137\
        );

    \I__9463\ : ClkMux
    port map (
            O => \N__37592\,
            I => \N__37137\
        );

    \I__9462\ : ClkMux
    port map (
            O => \N__37591\,
            I => \N__37137\
        );

    \I__9461\ : ClkMux
    port map (
            O => \N__37590\,
            I => \N__37137\
        );

    \I__9460\ : ClkMux
    port map (
            O => \N__37589\,
            I => \N__37137\
        );

    \I__9459\ : ClkMux
    port map (
            O => \N__37588\,
            I => \N__37137\
        );

    \I__9458\ : ClkMux
    port map (
            O => \N__37587\,
            I => \N__37137\
        );

    \I__9457\ : ClkMux
    port map (
            O => \N__37586\,
            I => \N__37137\
        );

    \I__9456\ : ClkMux
    port map (
            O => \N__37585\,
            I => \N__37137\
        );

    \I__9455\ : ClkMux
    port map (
            O => \N__37584\,
            I => \N__37137\
        );

    \I__9454\ : ClkMux
    port map (
            O => \N__37583\,
            I => \N__37137\
        );

    \I__9453\ : ClkMux
    port map (
            O => \N__37582\,
            I => \N__37137\
        );

    \I__9452\ : ClkMux
    port map (
            O => \N__37581\,
            I => \N__37137\
        );

    \I__9451\ : ClkMux
    port map (
            O => \N__37580\,
            I => \N__37137\
        );

    \I__9450\ : ClkMux
    port map (
            O => \N__37579\,
            I => \N__37137\
        );

    \I__9449\ : ClkMux
    port map (
            O => \N__37578\,
            I => \N__37137\
        );

    \I__9448\ : ClkMux
    port map (
            O => \N__37577\,
            I => \N__37137\
        );

    \I__9447\ : ClkMux
    port map (
            O => \N__37576\,
            I => \N__37137\
        );

    \I__9446\ : ClkMux
    port map (
            O => \N__37575\,
            I => \N__37137\
        );

    \I__9445\ : ClkMux
    port map (
            O => \N__37574\,
            I => \N__37137\
        );

    \I__9444\ : ClkMux
    port map (
            O => \N__37573\,
            I => \N__37137\
        );

    \I__9443\ : ClkMux
    port map (
            O => \N__37572\,
            I => \N__37137\
        );

    \I__9442\ : ClkMux
    port map (
            O => \N__37571\,
            I => \N__37137\
        );

    \I__9441\ : ClkMux
    port map (
            O => \N__37570\,
            I => \N__37137\
        );

    \I__9440\ : ClkMux
    port map (
            O => \N__37569\,
            I => \N__37137\
        );

    \I__9439\ : ClkMux
    port map (
            O => \N__37568\,
            I => \N__37137\
        );

    \I__9438\ : ClkMux
    port map (
            O => \N__37567\,
            I => \N__37137\
        );

    \I__9437\ : ClkMux
    port map (
            O => \N__37566\,
            I => \N__37137\
        );

    \I__9436\ : ClkMux
    port map (
            O => \N__37565\,
            I => \N__37137\
        );

    \I__9435\ : ClkMux
    port map (
            O => \N__37564\,
            I => \N__37137\
        );

    \I__9434\ : ClkMux
    port map (
            O => \N__37563\,
            I => \N__37137\
        );

    \I__9433\ : ClkMux
    port map (
            O => \N__37562\,
            I => \N__37137\
        );

    \I__9432\ : ClkMux
    port map (
            O => \N__37561\,
            I => \N__37137\
        );

    \I__9431\ : ClkMux
    port map (
            O => \N__37560\,
            I => \N__37137\
        );

    \I__9430\ : ClkMux
    port map (
            O => \N__37559\,
            I => \N__37137\
        );

    \I__9429\ : ClkMux
    port map (
            O => \N__37558\,
            I => \N__37137\
        );

    \I__9428\ : ClkMux
    port map (
            O => \N__37557\,
            I => \N__37137\
        );

    \I__9427\ : ClkMux
    port map (
            O => \N__37556\,
            I => \N__37137\
        );

    \I__9426\ : ClkMux
    port map (
            O => \N__37555\,
            I => \N__37137\
        );

    \I__9425\ : ClkMux
    port map (
            O => \N__37554\,
            I => \N__37137\
        );

    \I__9424\ : ClkMux
    port map (
            O => \N__37553\,
            I => \N__37137\
        );

    \I__9423\ : ClkMux
    port map (
            O => \N__37552\,
            I => \N__37137\
        );

    \I__9422\ : ClkMux
    port map (
            O => \N__37551\,
            I => \N__37137\
        );

    \I__9421\ : ClkMux
    port map (
            O => \N__37550\,
            I => \N__37137\
        );

    \I__9420\ : ClkMux
    port map (
            O => \N__37549\,
            I => \N__37137\
        );

    \I__9419\ : ClkMux
    port map (
            O => \N__37548\,
            I => \N__37137\
        );

    \I__9418\ : ClkMux
    port map (
            O => \N__37547\,
            I => \N__37137\
        );

    \I__9417\ : ClkMux
    port map (
            O => \N__37546\,
            I => \N__37137\
        );

    \I__9416\ : ClkMux
    port map (
            O => \N__37545\,
            I => \N__37137\
        );

    \I__9415\ : ClkMux
    port map (
            O => \N__37544\,
            I => \N__37137\
        );

    \I__9414\ : ClkMux
    port map (
            O => \N__37543\,
            I => \N__37137\
        );

    \I__9413\ : ClkMux
    port map (
            O => \N__37542\,
            I => \N__37137\
        );

    \I__9412\ : ClkMux
    port map (
            O => \N__37541\,
            I => \N__37137\
        );

    \I__9411\ : ClkMux
    port map (
            O => \N__37540\,
            I => \N__37137\
        );

    \I__9410\ : ClkMux
    port map (
            O => \N__37539\,
            I => \N__37137\
        );

    \I__9409\ : ClkMux
    port map (
            O => \N__37538\,
            I => \N__37137\
        );

    \I__9408\ : ClkMux
    port map (
            O => \N__37537\,
            I => \N__37137\
        );

    \I__9407\ : ClkMux
    port map (
            O => \N__37536\,
            I => \N__37137\
        );

    \I__9406\ : ClkMux
    port map (
            O => \N__37535\,
            I => \N__37137\
        );

    \I__9405\ : ClkMux
    port map (
            O => \N__37534\,
            I => \N__37137\
        );

    \I__9404\ : ClkMux
    port map (
            O => \N__37533\,
            I => \N__37137\
        );

    \I__9403\ : ClkMux
    port map (
            O => \N__37532\,
            I => \N__37137\
        );

    \I__9402\ : ClkMux
    port map (
            O => \N__37531\,
            I => \N__37137\
        );

    \I__9401\ : ClkMux
    port map (
            O => \N__37530\,
            I => \N__37137\
        );

    \I__9400\ : ClkMux
    port map (
            O => \N__37529\,
            I => \N__37137\
        );

    \I__9399\ : ClkMux
    port map (
            O => \N__37528\,
            I => \N__37137\
        );

    \I__9398\ : ClkMux
    port map (
            O => \N__37527\,
            I => \N__37137\
        );

    \I__9397\ : ClkMux
    port map (
            O => \N__37526\,
            I => \N__37137\
        );

    \I__9396\ : ClkMux
    port map (
            O => \N__37525\,
            I => \N__37137\
        );

    \I__9395\ : ClkMux
    port map (
            O => \N__37524\,
            I => \N__37137\
        );

    \I__9394\ : ClkMux
    port map (
            O => \N__37523\,
            I => \N__37137\
        );

    \I__9393\ : ClkMux
    port map (
            O => \N__37522\,
            I => \N__37137\
        );

    \I__9392\ : ClkMux
    port map (
            O => \N__37521\,
            I => \N__37137\
        );

    \I__9391\ : ClkMux
    port map (
            O => \N__37520\,
            I => \N__37137\
        );

    \I__9390\ : ClkMux
    port map (
            O => \N__37519\,
            I => \N__37137\
        );

    \I__9389\ : ClkMux
    port map (
            O => \N__37518\,
            I => \N__37137\
        );

    \I__9388\ : ClkMux
    port map (
            O => \N__37517\,
            I => \N__37137\
        );

    \I__9387\ : ClkMux
    port map (
            O => \N__37516\,
            I => \N__37137\
        );

    \I__9386\ : ClkMux
    port map (
            O => \N__37515\,
            I => \N__37137\
        );

    \I__9385\ : ClkMux
    port map (
            O => \N__37514\,
            I => \N__37137\
        );

    \I__9384\ : ClkMux
    port map (
            O => \N__37513\,
            I => \N__37137\
        );

    \I__9383\ : ClkMux
    port map (
            O => \N__37512\,
            I => \N__37137\
        );

    \I__9382\ : ClkMux
    port map (
            O => \N__37511\,
            I => \N__37137\
        );

    \I__9381\ : ClkMux
    port map (
            O => \N__37510\,
            I => \N__37137\
        );

    \I__9380\ : ClkMux
    port map (
            O => \N__37509\,
            I => \N__37137\
        );

    \I__9379\ : ClkMux
    port map (
            O => \N__37508\,
            I => \N__37137\
        );

    \I__9378\ : ClkMux
    port map (
            O => \N__37507\,
            I => \N__37137\
        );

    \I__9377\ : ClkMux
    port map (
            O => \N__37506\,
            I => \N__37137\
        );

    \I__9376\ : ClkMux
    port map (
            O => \N__37505\,
            I => \N__37137\
        );

    \I__9375\ : ClkMux
    port map (
            O => \N__37504\,
            I => \N__37137\
        );

    \I__9374\ : ClkMux
    port map (
            O => \N__37503\,
            I => \N__37137\
        );

    \I__9373\ : ClkMux
    port map (
            O => \N__37502\,
            I => \N__37137\
        );

    \I__9372\ : ClkMux
    port map (
            O => \N__37501\,
            I => \N__37137\
        );

    \I__9371\ : ClkMux
    port map (
            O => \N__37500\,
            I => \N__37137\
        );

    \I__9370\ : ClkMux
    port map (
            O => \N__37499\,
            I => \N__37137\
        );

    \I__9369\ : ClkMux
    port map (
            O => \N__37498\,
            I => \N__37137\
        );

    \I__9368\ : ClkMux
    port map (
            O => \N__37497\,
            I => \N__37137\
        );

    \I__9367\ : ClkMux
    port map (
            O => \N__37496\,
            I => \N__37137\
        );

    \I__9366\ : ClkMux
    port map (
            O => \N__37495\,
            I => \N__37137\
        );

    \I__9365\ : ClkMux
    port map (
            O => \N__37494\,
            I => \N__37137\
        );

    \I__9364\ : ClkMux
    port map (
            O => \N__37493\,
            I => \N__37137\
        );

    \I__9363\ : ClkMux
    port map (
            O => \N__37492\,
            I => \N__37137\
        );

    \I__9362\ : ClkMux
    port map (
            O => \N__37491\,
            I => \N__37137\
        );

    \I__9361\ : ClkMux
    port map (
            O => \N__37490\,
            I => \N__37137\
        );

    \I__9360\ : ClkMux
    port map (
            O => \N__37489\,
            I => \N__37137\
        );

    \I__9359\ : ClkMux
    port map (
            O => \N__37488\,
            I => \N__37137\
        );

    \I__9358\ : ClkMux
    port map (
            O => \N__37487\,
            I => \N__37137\
        );

    \I__9357\ : ClkMux
    port map (
            O => \N__37486\,
            I => \N__37137\
        );

    \I__9356\ : ClkMux
    port map (
            O => \N__37485\,
            I => \N__37137\
        );

    \I__9355\ : ClkMux
    port map (
            O => \N__37484\,
            I => \N__37137\
        );

    \I__9354\ : ClkMux
    port map (
            O => \N__37483\,
            I => \N__37137\
        );

    \I__9353\ : ClkMux
    port map (
            O => \N__37482\,
            I => \N__37137\
        );

    \I__9352\ : ClkMux
    port map (
            O => \N__37481\,
            I => \N__37137\
        );

    \I__9351\ : ClkMux
    port map (
            O => \N__37480\,
            I => \N__37137\
        );

    \I__9350\ : ClkMux
    port map (
            O => \N__37479\,
            I => \N__37137\
        );

    \I__9349\ : ClkMux
    port map (
            O => \N__37478\,
            I => \N__37137\
        );

    \I__9348\ : ClkMux
    port map (
            O => \N__37477\,
            I => \N__37137\
        );

    \I__9347\ : ClkMux
    port map (
            O => \N__37476\,
            I => \N__37137\
        );

    \I__9346\ : ClkMux
    port map (
            O => \N__37475\,
            I => \N__37137\
        );

    \I__9345\ : ClkMux
    port map (
            O => \N__37474\,
            I => \N__37137\
        );

    \I__9344\ : ClkMux
    port map (
            O => \N__37473\,
            I => \N__37137\
        );

    \I__9343\ : ClkMux
    port map (
            O => \N__37472\,
            I => \N__37137\
        );

    \I__9342\ : ClkMux
    port map (
            O => \N__37471\,
            I => \N__37137\
        );

    \I__9341\ : ClkMux
    port map (
            O => \N__37470\,
            I => \N__37137\
        );

    \I__9340\ : ClkMux
    port map (
            O => \N__37469\,
            I => \N__37137\
        );

    \I__9339\ : ClkMux
    port map (
            O => \N__37468\,
            I => \N__37137\
        );

    \I__9338\ : ClkMux
    port map (
            O => \N__37467\,
            I => \N__37137\
        );

    \I__9337\ : ClkMux
    port map (
            O => \N__37466\,
            I => \N__37137\
        );

    \I__9336\ : ClkMux
    port map (
            O => \N__37465\,
            I => \N__37137\
        );

    \I__9335\ : ClkMux
    port map (
            O => \N__37464\,
            I => \N__37137\
        );

    \I__9334\ : ClkMux
    port map (
            O => \N__37463\,
            I => \N__37137\
        );

    \I__9333\ : ClkMux
    port map (
            O => \N__37462\,
            I => \N__37137\
        );

    \I__9332\ : GlobalMux
    port map (
            O => \N__37137\,
            I => \N__37134\
        );

    \I__9331\ : gio2CtrlBuf
    port map (
            O => \N__37134\,
            I => \CLK_c\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__37131\,
            I => \N__37128\
        );

    \I__9329\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37125\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__37125\,
            I => \N__37121\
        );

    \I__9327\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37118\
        );

    \I__9326\ : Odrv12
    port map (
            O => \N__37121\,
            I => data_3
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__37118\,
            I => data_3
        );

    \I__9324\ : InMux
    port map (
            O => \N__37113\,
            I => \c0.n4741\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__37110\,
            I => \N__37107\
        );

    \I__9322\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37104\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__37104\,
            I => \N__37101\
        );

    \I__9320\ : Span4Mux_h
    port map (
            O => \N__37101\,
            I => \N__37097\
        );

    \I__9319\ : InMux
    port map (
            O => \N__37100\,
            I => \N__37094\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__37097\,
            I => data_4
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__37094\,
            I => data_4
        );

    \I__9316\ : InMux
    port map (
            O => \N__37089\,
            I => \c0.n4742\
        );

    \I__9315\ : CascadeMux
    port map (
            O => \N__37086\,
            I => \N__37083\
        );

    \I__9314\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37080\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37076\
        );

    \I__9312\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37073\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__37076\,
            I => data_5
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__37073\,
            I => data_5
        );

    \I__9309\ : InMux
    port map (
            O => \N__37068\,
            I => \c0.n4743\
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__37065\,
            I => \N__37062\
        );

    \I__9307\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37059\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__37059\,
            I => \N__37055\
        );

    \I__9305\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37052\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__37055\,
            I => data_6
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__37052\,
            I => data_6
        );

    \I__9302\ : InMux
    port map (
            O => \N__37047\,
            I => \c0.n4744\
        );

    \I__9301\ : CascadeMux
    port map (
            O => \N__37044\,
            I => \N__37041\
        );

    \I__9300\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37038\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__37038\,
            I => \N__37034\
        );

    \I__9298\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37031\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__37034\,
            I => data_7
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__37031\,
            I => data_7
        );

    \I__9295\ : InMux
    port map (
            O => \N__37026\,
            I => \c0.n4745\
        );

    \I__9294\ : InMux
    port map (
            O => \N__37023\,
            I => \N__37020\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__37020\,
            I => \N__37016\
        );

    \I__9292\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37013\
        );

    \I__9291\ : Odrv4
    port map (
            O => \N__37016\,
            I => data_8
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__37013\,
            I => data_8
        );

    \I__9289\ : InMux
    port map (
            O => \N__37008\,
            I => \bfn_15_27_0_\
        );

    \I__9288\ : InMux
    port map (
            O => \N__37005\,
            I => \N__37002\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__37002\,
            I => \N__36999\
        );

    \I__9286\ : Span4Mux_h
    port map (
            O => \N__36999\,
            I => \N__36995\
        );

    \I__9285\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36992\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__36995\,
            I => data_9
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__36992\,
            I => data_9
        );

    \I__9282\ : InMux
    port map (
            O => \N__36987\,
            I => \c0.n4747\
        );

    \I__9281\ : CascadeMux
    port map (
            O => \N__36984\,
            I => \N__36981\
        );

    \I__9280\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36977\
        );

    \I__9279\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36974\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__36977\,
            I => data_10
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__36974\,
            I => data_10
        );

    \I__9276\ : InMux
    port map (
            O => \N__36969\,
            I => \c0.n4748\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__36966\,
            I => \N__36961\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__36965\,
            I => \N__36958\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__36964\,
            I => \N__36955\
        );

    \I__9272\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36949\
        );

    \I__9271\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36949\
        );

    \I__9270\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36946\
        );

    \I__9269\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36942\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__36949\,
            I => \N__36939\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36936\
        );

    \I__9266\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36932\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__36942\,
            I => \N__36929\
        );

    \I__9264\ : Span4Mux_h
    port map (
            O => \N__36939\,
            I => \N__36924\
        );

    \I__9263\ : Span4Mux_h
    port map (
            O => \N__36936\,
            I => \N__36924\
        );

    \I__9262\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36921\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__36932\,
            I => data_out_11_2
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__36929\,
            I => data_out_11_2
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__36924\,
            I => data_out_11_2
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__36921\,
            I => data_out_11_2
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__36912\,
            I => \N__36906\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__36911\,
            I => \N__36903\
        );

    \I__9255\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36887\
        );

    \I__9254\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36887\
        );

    \I__9253\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36884\
        );

    \I__9252\ : InMux
    port map (
            O => \N__36903\,
            I => \N__36877\
        );

    \I__9251\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36877\
        );

    \I__9250\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36877\
        );

    \I__9249\ : InMux
    port map (
            O => \N__36900\,
            I => \N__36874\
        );

    \I__9248\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36871\
        );

    \I__9247\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36868\
        );

    \I__9246\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36865\
        );

    \I__9245\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36862\
        );

    \I__9244\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36855\
        );

    \I__9243\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36855\
        );

    \I__9242\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36855\
        );

    \I__9241\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36852\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__36887\,
            I => \N__36849\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36842\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36842\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__36874\,
            I => \N__36842\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36837\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36837\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36832\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36832\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__36855\,
            I => \N__36829\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__36852\,
            I => \N__36814\
        );

    \I__9230\ : Span4Mux_h
    port map (
            O => \N__36849\,
            I => \N__36814\
        );

    \I__9229\ : Span4Mux_v
    port map (
            O => \N__36842\,
            I => \N__36814\
        );

    \I__9228\ : Span4Mux_v
    port map (
            O => \N__36837\,
            I => \N__36814\
        );

    \I__9227\ : Span4Mux_v
    port map (
            O => \N__36832\,
            I => \N__36814\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__36829\,
            I => \N__36811\
        );

    \I__9225\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36806\
        );

    \I__9224\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36806\
        );

    \I__9223\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36801\
        );

    \I__9222\ : InMux
    port map (
            O => \N__36825\,
            I => \N__36801\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__36814\,
            I => n21_adj_1977
        );

    \I__9220\ : Odrv4
    port map (
            O => \N__36811\,
            I => n21_adj_1977
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__36806\,
            I => n21_adj_1977
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__36801\,
            I => n21_adj_1977
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__36792\,
            I => \N__36780\
        );

    \I__9216\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36777\
        );

    \I__9215\ : InMux
    port map (
            O => \N__36790\,
            I => \N__36772\
        );

    \I__9214\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36772\
        );

    \I__9213\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36763\
        );

    \I__9212\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36763\
        );

    \I__9211\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36756\
        );

    \I__9210\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36756\
        );

    \I__9209\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36756\
        );

    \I__9208\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36753\
        );

    \I__9207\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36749\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__36777\,
            I => \N__36745\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__36772\,
            I => \N__36742\
        );

    \I__9204\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36733\
        );

    \I__9203\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36733\
        );

    \I__9202\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36733\
        );

    \I__9201\ : InMux
    port map (
            O => \N__36768\,
            I => \N__36733\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__36763\,
            I => \N__36724\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__36756\,
            I => \N__36724\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__36753\,
            I => \N__36724\
        );

    \I__9197\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36721\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__36749\,
            I => \N__36718\
        );

    \I__9195\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36715\
        );

    \I__9194\ : Span4Mux_v
    port map (
            O => \N__36745\,
            I => \N__36708\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__36742\,
            I => \N__36708\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__36733\,
            I => \N__36708\
        );

    \I__9191\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36703\
        );

    \I__9190\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36703\
        );

    \I__9189\ : Span4Mux_v
    port map (
            O => \N__36724\,
            I => \N__36696\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__36721\,
            I => \N__36696\
        );

    \I__9187\ : Span4Mux_v
    port map (
            O => \N__36718\,
            I => \N__36696\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__36715\,
            I => n4333
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__36708\,
            I => n4333
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__36703\,
            I => n4333
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__36696\,
            I => n4333
        );

    \I__9182\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36684\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__36684\,
            I => \N__36677\
        );

    \I__9180\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36674\
        );

    \I__9179\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36671\
        );

    \I__9178\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36668\
        );

    \I__9177\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36663\
        );

    \I__9176\ : Span4Mux_v
    port map (
            O => \N__36677\,
            I => \N__36654\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36654\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36654\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36654\
        );

    \I__9172\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36649\
        );

    \I__9171\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36649\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__36663\,
            I => data_out_10_1
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__36654\,
            I => data_out_10_1
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__36649\,
            I => data_out_10_1
        );

    \I__9167\ : InMux
    port map (
            O => \N__36642\,
            I => \N__36636\
        );

    \I__9166\ : InMux
    port map (
            O => \N__36641\,
            I => \N__36632\
        );

    \I__9165\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36629\
        );

    \I__9164\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36626\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__36636\,
            I => \N__36623\
        );

    \I__9162\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36620\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__36632\,
            I => \N__36615\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__36629\,
            I => \N__36615\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__36626\,
            I => \N__36609\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__36623\,
            I => \N__36609\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36606\
        );

    \I__9156\ : Span4Mux_h
    port map (
            O => \N__36615\,
            I => \N__36603\
        );

    \I__9155\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36600\
        );

    \I__9154\ : Odrv4
    port map (
            O => \N__36609\,
            I => data_out_10_3
        );

    \I__9153\ : Odrv4
    port map (
            O => \N__36606\,
            I => data_out_10_3
        );

    \I__9152\ : Odrv4
    port map (
            O => \N__36603\,
            I => data_out_10_3
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__36600\,
            I => data_out_10_3
        );

    \I__9150\ : CascadeMux
    port map (
            O => \N__36591\,
            I => \N__36588\
        );

    \I__9149\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36584\
        );

    \I__9148\ : CascadeMux
    port map (
            O => \N__36587\,
            I => \N__36581\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__36584\,
            I => \N__36578\
        );

    \I__9146\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36575\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__36578\,
            I => \N__36570\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__36575\,
            I => \N__36570\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__36570\,
            I => n5424
        );

    \I__9142\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36561\
        );

    \I__9141\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36558\
        );

    \I__9140\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36555\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__36564\,
            I => \N__36551\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__36561\,
            I => \N__36547\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__36558\,
            I => \N__36542\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__36555\,
            I => \N__36542\
        );

    \I__9135\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36537\
        );

    \I__9134\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36537\
        );

    \I__9133\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36534\
        );

    \I__9132\ : Span4Mux_h
    port map (
            O => \N__36547\,
            I => \N__36531\
        );

    \I__9131\ : Span4Mux_h
    port map (
            O => \N__36542\,
            I => \N__36526\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__36537\,
            I => \N__36526\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__36534\,
            I => data_out_11_0
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__36531\,
            I => data_out_11_0
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__36526\,
            I => data_out_11_0
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__36519\,
            I => \N__36515\
        );

    \I__9125\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36512\
        );

    \I__9124\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36509\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__36512\,
            I => \N__36501\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36501\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__36508\,
            I => \N__36496\
        );

    \I__9120\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36492\
        );

    \I__9119\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36489\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__36501\,
            I => \N__36486\
        );

    \I__9117\ : CascadeMux
    port map (
            O => \N__36500\,
            I => \N__36483\
        );

    \I__9116\ : InMux
    port map (
            O => \N__36499\,
            I => \N__36480\
        );

    \I__9115\ : InMux
    port map (
            O => \N__36496\,
            I => \N__36475\
        );

    \I__9114\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36475\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36472\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__36489\,
            I => \N__36469\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__36486\,
            I => \N__36466\
        );

    \I__9110\ : InMux
    port map (
            O => \N__36483\,
            I => \N__36463\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36458\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__36475\,
            I => \N__36458\
        );

    \I__9107\ : Span4Mux_h
    port map (
            O => \N__36472\,
            I => \N__36455\
        );

    \I__9106\ : Span4Mux_v
    port map (
            O => \N__36469\,
            I => \N__36450\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__36466\,
            I => \N__36450\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__36463\,
            I => data_out_10_7
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__36458\,
            I => data_out_10_7
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__36455\,
            I => data_out_10_7
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__36450\,
            I => data_out_10_7
        );

    \I__9100\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36437\
        );

    \I__9099\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36434\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__36437\,
            I => \N__36431\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36427\
        );

    \I__9096\ : Span4Mux_h
    port map (
            O => \N__36431\,
            I => \N__36424\
        );

    \I__9095\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36421\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__36427\,
            I => n5479
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__36424\,
            I => n5479
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__36421\,
            I => n5479
        );

    \I__9091\ : CascadeMux
    port map (
            O => \N__36414\,
            I => \N__36409\
        );

    \I__9090\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36403\
        );

    \I__9089\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36403\
        );

    \I__9088\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36400\
        );

    \I__9087\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36396\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__36403\,
            I => \N__36393\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__36400\,
            I => \N__36387\
        );

    \I__9084\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36384\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__36396\,
            I => \N__36381\
        );

    \I__9082\ : Span4Mux_h
    port map (
            O => \N__36393\,
            I => \N__36378\
        );

    \I__9081\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36371\
        );

    \I__9080\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36371\
        );

    \I__9079\ : InMux
    port map (
            O => \N__36390\,
            I => \N__36371\
        );

    \I__9078\ : Span4Mux_h
    port map (
            O => \N__36387\,
            I => \N__36368\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__36384\,
            I => data_out_11_3
        );

    \I__9076\ : Odrv4
    port map (
            O => \N__36381\,
            I => data_out_11_3
        );

    \I__9075\ : Odrv4
    port map (
            O => \N__36378\,
            I => data_out_11_3
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__36371\,
            I => data_out_11_3
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__36368\,
            I => data_out_11_3
        );

    \I__9072\ : InMux
    port map (
            O => \N__36357\,
            I => \N__36354\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__36354\,
            I => n8_adj_1984
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__36351\,
            I => \n7_adj_1985_cascade_\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__36348\,
            I => \N__36345\
        );

    \I__9068\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36342\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N__36338\
        );

    \I__9066\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36335\
        );

    \I__9065\ : Span4Mux_h
    port map (
            O => \N__36338\,
            I => \N__36332\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__36335\,
            I => data_out_19_1
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__36332\,
            I => data_out_19_1
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__36327\,
            I => \N__36324\
        );

    \I__9061\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36321\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__36321\,
            I => \N__36318\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__36318\,
            I => \N__36314\
        );

    \I__9058\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36311\
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__36314\,
            I => data_0
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__36311\,
            I => data_0
        );

    \I__9055\ : InMux
    port map (
            O => \N__36306\,
            I => \bfn_15_26_0_\
        );

    \I__9054\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36300\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__36300\,
            I => \N__36297\
        );

    \I__9052\ : Span4Mux_h
    port map (
            O => \N__36297\,
            I => \N__36293\
        );

    \I__9051\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36290\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__36293\,
            I => data_1
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__36290\,
            I => data_1
        );

    \I__9048\ : InMux
    port map (
            O => \N__36285\,
            I => \c0.n4739\
        );

    \I__9047\ : CascadeMux
    port map (
            O => \N__36282\,
            I => \N__36279\
        );

    \I__9046\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__36276\,
            I => \N__36272\
        );

    \I__9044\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36269\
        );

    \I__9043\ : Odrv4
    port map (
            O => \N__36272\,
            I => data_2
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__36269\,
            I => data_2
        );

    \I__9041\ : InMux
    port map (
            O => \N__36264\,
            I => \c0.n4740\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__36261\,
            I => \N__36257\
        );

    \I__9039\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36252\
        );

    \I__9038\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36252\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__36252\,
            I => \N__36249\
        );

    \I__9036\ : Span4Mux_h
    port map (
            O => \N__36249\,
            I => \N__36245\
        );

    \I__9035\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36242\
        );

    \I__9034\ : Odrv4
    port map (
            O => \N__36245\,
            I => blink_counter_23
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__36242\,
            I => blink_counter_23
        );

    \I__9032\ : InMux
    port map (
            O => \N__36237\,
            I => n4732
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__36234\,
            I => \N__36231\
        );

    \I__9030\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36225\
        );

    \I__9029\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36225\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__9027\ : Span12Mux_h
    port map (
            O => \N__36222\,
            I => \N__36218\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36215\
        );

    \I__9025\ : Odrv12
    port map (
            O => \N__36218\,
            I => blink_counter_24
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__36215\,
            I => blink_counter_24
        );

    \I__9023\ : InMux
    port map (
            O => \N__36210\,
            I => \bfn_14_28_0_\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36207\,
            I => n4734
        );

    \I__9021\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36201\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__36201\,
            I => \N__36198\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__36198\,
            I => \N__36195\
        );

    \I__9018\ : Span4Mux_v
    port map (
            O => \N__36195\,
            I => \N__36191\
        );

    \I__9017\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36188\
        );

    \I__9016\ : Odrv4
    port map (
            O => \N__36191\,
            I => blink_counter_25
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__36188\,
            I => blink_counter_25
        );

    \I__9014\ : CascadeMux
    port map (
            O => \N__36183\,
            I => \N__36180\
        );

    \I__9013\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36177\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36170\
        );

    \I__9011\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36166\
        );

    \I__9010\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36163\
        );

    \I__9009\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36160\
        );

    \I__9008\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36157\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__36170\,
            I => \N__36154\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36151\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__36166\,
            I => \N__36147\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36140\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36140\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__36140\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__36154\,
            I => \N__36135\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36135\
        );

    \I__8999\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36132\
        );

    \I__8998\ : Span4Mux_h
    port map (
            O => \N__36147\,
            I => \N__36125\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__36140\,
            I => \N__36125\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__36135\,
            I => \N__36125\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__36132\,
            I => data_out_10_2
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__36125\,
            I => data_out_10_2
        );

    \I__8993\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36116\
        );

    \I__8992\ : InMux
    port map (
            O => \N__36119\,
            I => \N__36113\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__36116\,
            I => \N__36105\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__36113\,
            I => \N__36102\
        );

    \I__8989\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36097\
        );

    \I__8988\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36097\
        );

    \I__8987\ : InMux
    port map (
            O => \N__36110\,
            I => \N__36094\
        );

    \I__8986\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36089\
        );

    \I__8985\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36089\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__36105\,
            I => \N__36082\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__36102\,
            I => \N__36082\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__36097\,
            I => \N__36082\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__36094\,
            I => data_out_11_6
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__36089\,
            I => data_out_11_6
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__36082\,
            I => data_out_11_6
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__36075\,
            I => \N__36065\
        );

    \I__8977\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36059\
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__36073\,
            I => \N__36049\
        );

    \I__8975\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36040\
        );

    \I__8974\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36035\
        );

    \I__8973\ : InMux
    port map (
            O => \N__36070\,
            I => \N__36035\
        );

    \I__8972\ : InMux
    port map (
            O => \N__36069\,
            I => \N__36032\
        );

    \I__8971\ : InMux
    port map (
            O => \N__36068\,
            I => \N__36025\
        );

    \I__8970\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36025\
        );

    \I__8969\ : InMux
    port map (
            O => \N__36064\,
            I => \N__36025\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__36063\,
            I => \N__36016\
        );

    \I__8967\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36011\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__36008\
        );

    \I__8965\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36001\
        );

    \I__8964\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36001\
        );

    \I__8963\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36001\
        );

    \I__8962\ : InMux
    port map (
            O => \N__36055\,
            I => \N__35992\
        );

    \I__8961\ : InMux
    port map (
            O => \N__36054\,
            I => \N__35992\
        );

    \I__8960\ : InMux
    port map (
            O => \N__36053\,
            I => \N__35992\
        );

    \I__8959\ : InMux
    port map (
            O => \N__36052\,
            I => \N__35987\
        );

    \I__8958\ : InMux
    port map (
            O => \N__36049\,
            I => \N__35987\
        );

    \I__8957\ : InMux
    port map (
            O => \N__36048\,
            I => \N__35984\
        );

    \I__8956\ : InMux
    port map (
            O => \N__36047\,
            I => \N__35971\
        );

    \I__8955\ : InMux
    port map (
            O => \N__36046\,
            I => \N__35966\
        );

    \I__8954\ : InMux
    port map (
            O => \N__36045\,
            I => \N__35966\
        );

    \I__8953\ : InMux
    port map (
            O => \N__36044\,
            I => \N__35957\
        );

    \I__8952\ : InMux
    port map (
            O => \N__36043\,
            I => \N__35957\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__36040\,
            I => \N__35948\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__35948\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__35948\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__35948\
        );

    \I__8947\ : InMux
    port map (
            O => \N__36024\,
            I => \N__35945\
        );

    \I__8946\ : CascadeMux
    port map (
            O => \N__36023\,
            I => \N__35936\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__36022\,
            I => \N__35920\
        );

    \I__8944\ : InMux
    port map (
            O => \N__36021\,
            I => \N__35911\
        );

    \I__8943\ : InMux
    port map (
            O => \N__36020\,
            I => \N__35911\
        );

    \I__8942\ : InMux
    port map (
            O => \N__36019\,
            I => \N__35911\
        );

    \I__8941\ : InMux
    port map (
            O => \N__36016\,
            I => \N__35908\
        );

    \I__8940\ : InMux
    port map (
            O => \N__36015\,
            I => \N__35894\
        );

    \I__8939\ : InMux
    port map (
            O => \N__36014\,
            I => \N__35894\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__36011\,
            I => \N__35887\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__36008\,
            I => \N__35887\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35887\
        );

    \I__8935\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35884\
        );

    \I__8934\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35881\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__35992\,
            I => \N__35869\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__35987\,
            I => \N__35869\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__35984\,
            I => \N__35869\
        );

    \I__8930\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35862\
        );

    \I__8929\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35862\
        );

    \I__8928\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35862\
        );

    \I__8927\ : InMux
    port map (
            O => \N__35980\,
            I => \N__35857\
        );

    \I__8926\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35857\
        );

    \I__8925\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35854\
        );

    \I__8924\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35850\
        );

    \I__8923\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35847\
        );

    \I__8922\ : InMux
    port map (
            O => \N__35975\,
            I => \N__35844\
        );

    \I__8921\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35841\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__35971\,
            I => \N__35836\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__35966\,
            I => \N__35836\
        );

    \I__8918\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35831\
        );

    \I__8917\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35831\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__35963\,
            I => \N__35813\
        );

    \I__8915\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35809\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__35957\,
            I => \N__35802\
        );

    \I__8913\ : Span4Mux_v
    port map (
            O => \N__35948\,
            I => \N__35802\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__35945\,
            I => \N__35802\
        );

    \I__8911\ : InMux
    port map (
            O => \N__35944\,
            I => \N__35797\
        );

    \I__8910\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35797\
        );

    \I__8909\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35792\
        );

    \I__8908\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35792\
        );

    \I__8907\ : InMux
    port map (
            O => \N__35940\,
            I => \N__35789\
        );

    \I__8906\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35782\
        );

    \I__8905\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35782\
        );

    \I__8904\ : InMux
    port map (
            O => \N__35935\,
            I => \N__35782\
        );

    \I__8903\ : InMux
    port map (
            O => \N__35934\,
            I => \N__35775\
        );

    \I__8902\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35775\
        );

    \I__8901\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35775\
        );

    \I__8900\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35766\
        );

    \I__8899\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35766\
        );

    \I__8898\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35766\
        );

    \I__8897\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35766\
        );

    \I__8896\ : InMux
    port map (
            O => \N__35927\,
            I => \N__35761\
        );

    \I__8895\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35761\
        );

    \I__8894\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35757\
        );

    \I__8893\ : InMux
    port map (
            O => \N__35924\,
            I => \N__35754\
        );

    \I__8892\ : InMux
    port map (
            O => \N__35923\,
            I => \N__35751\
        );

    \I__8891\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35744\
        );

    \I__8890\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35744\
        );

    \I__8889\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35744\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__35911\,
            I => \N__35741\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35738\
        );

    \I__8886\ : InMux
    port map (
            O => \N__35907\,
            I => \N__35731\
        );

    \I__8885\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35731\
        );

    \I__8884\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35731\
        );

    \I__8883\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35728\
        );

    \I__8882\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35725\
        );

    \I__8881\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35720\
        );

    \I__8880\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35720\
        );

    \I__8879\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35716\
        );

    \I__8878\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35713\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35704\
        );

    \I__8876\ : Span4Mux_v
    port map (
            O => \N__35887\,
            I => \N__35704\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__35884\,
            I => \N__35704\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__35881\,
            I => \N__35704\
        );

    \I__8873\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35699\
        );

    \I__8872\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35699\
        );

    \I__8871\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35694\
        );

    \I__8870\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35694\
        );

    \I__8869\ : CascadeMux
    port map (
            O => \N__35876\,
            I => \N__35690\
        );

    \I__8868\ : Span4Mux_v
    port map (
            O => \N__35869\,
            I => \N__35674\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__35862\,
            I => \N__35674\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__35857\,
            I => \N__35674\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35671\
        );

    \I__8864\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35668\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__35850\,
            I => \N__35659\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35659\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__35844\,
            I => \N__35659\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__35841\,
            I => \N__35659\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__35836\,
            I => \N__35654\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__35831\,
            I => \N__35654\
        );

    \I__8857\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35651\
        );

    \I__8856\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35642\
        );

    \I__8855\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35642\
        );

    \I__8854\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35642\
        );

    \I__8853\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35642\
        );

    \I__8852\ : CascadeMux
    port map (
            O => \N__35825\,
            I => \N__35637\
        );

    \I__8851\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35623\
        );

    \I__8850\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35623\
        );

    \I__8849\ : InMux
    port map (
            O => \N__35822\,
            I => \N__35616\
        );

    \I__8848\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35616\
        );

    \I__8847\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35616\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35607\
        );

    \I__8845\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35607\
        );

    \I__8844\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35607\
        );

    \I__8843\ : InMux
    port map (
            O => \N__35816\,
            I => \N__35607\
        );

    \I__8842\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35604\
        );

    \I__8841\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35601\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35594\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__35802\,
            I => \N__35594\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35594\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35591\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35584\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__35782\,
            I => \N__35584\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35584\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35581\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__35761\,
            I => \N__35578\
        );

    \I__8831\ : InMux
    port map (
            O => \N__35760\,
            I => \N__35575\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35570\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__35754\,
            I => \N__35570\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35559\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__35744\,
            I => \N__35559\
        );

    \I__8826\ : Span4Mux_v
    port map (
            O => \N__35741\,
            I => \N__35559\
        );

    \I__8825\ : Span4Mux_v
    port map (
            O => \N__35738\,
            I => \N__35559\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__35731\,
            I => \N__35559\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__35728\,
            I => \N__35550\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35550\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35550\
        );

    \I__8820\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35547\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35536\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35536\
        );

    \I__8817\ : Span4Mux_h
    port map (
            O => \N__35704\,
            I => \N__35536\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__35699\,
            I => \N__35536\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__35694\,
            I => \N__35536\
        );

    \I__8814\ : InMux
    port map (
            O => \N__35693\,
            I => \N__35533\
        );

    \I__8813\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35524\
        );

    \I__8812\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35524\
        );

    \I__8811\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35524\
        );

    \I__8810\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35524\
        );

    \I__8809\ : InMux
    port map (
            O => \N__35686\,
            I => \N__35519\
        );

    \I__8808\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35519\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__35684\,
            I => \N__35512\
        );

    \I__8806\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35506\
        );

    \I__8805\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35503\
        );

    \I__8804\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35496\
        );

    \I__8803\ : Span4Mux_h
    port map (
            O => \N__35674\,
            I => \N__35489\
        );

    \I__8802\ : Span4Mux_v
    port map (
            O => \N__35671\,
            I => \N__35489\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__35668\,
            I => \N__35489\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__35659\,
            I => \N__35486\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__35654\,
            I => \N__35479\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35479\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35479\
        );

    \I__8796\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35474\
        );

    \I__8795\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35471\
        );

    \I__8794\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35466\
        );

    \I__8793\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35466\
        );

    \I__8792\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35457\
        );

    \I__8791\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35457\
        );

    \I__8790\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35457\
        );

    \I__8789\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35457\
        );

    \I__8788\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35454\
        );

    \I__8787\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35451\
        );

    \I__8786\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35443\
        );

    \I__8785\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35443\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__35623\,
            I => \N__35436\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__35616\,
            I => \N__35436\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__35607\,
            I => \N__35436\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35433\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__35601\,
            I => \N__35430\
        );

    \I__8779\ : Span4Mux_v
    port map (
            O => \N__35594\,
            I => \N__35427\
        );

    \I__8778\ : Span4Mux_s3_h
    port map (
            O => \N__35591\,
            I => \N__35422\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__35584\,
            I => \N__35422\
        );

    \I__8776\ : Span4Mux_v
    port map (
            O => \N__35581\,
            I => \N__35419\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__35578\,
            I => \N__35416\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__35575\,
            I => \N__35413\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__35570\,
            I => \N__35408\
        );

    \I__8772\ : Span4Mux_v
    port map (
            O => \N__35559\,
            I => \N__35408\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__35558\,
            I => \N__35402\
        );

    \I__8770\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35398\
        );

    \I__8769\ : Span4Mux_v
    port map (
            O => \N__35550\,
            I => \N__35385\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35385\
        );

    \I__8767\ : Span4Mux_v
    port map (
            O => \N__35536\,
            I => \N__35385\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__35533\,
            I => \N__35385\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35385\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35385\
        );

    \I__8763\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35381\
        );

    \I__8762\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35378\
        );

    \I__8761\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35373\
        );

    \I__8760\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35373\
        );

    \I__8759\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35368\
        );

    \I__8758\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35368\
        );

    \I__8757\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35363\
        );

    \I__8756\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35363\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__35506\,
            I => \N__35358\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35358\
        );

    \I__8753\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35353\
        );

    \I__8752\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35353\
        );

    \I__8751\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35350\
        );

    \I__8750\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35339\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__35496\,
            I => \N__35330\
        );

    \I__8748\ : Span4Mux_h
    port map (
            O => \N__35489\,
            I => \N__35330\
        );

    \I__8747\ : Span4Mux_s1_h
    port map (
            O => \N__35486\,
            I => \N__35330\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35330\
        );

    \I__8745\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35325\
        );

    \I__8744\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35325\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__35474\,
            I => \N__35322\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35311\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__35466\,
            I => \N__35311\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__35457\,
            I => \N__35311\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__35454\,
            I => \N__35311\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__35451\,
            I => \N__35311\
        );

    \I__8737\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35306\
        );

    \I__8736\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35306\
        );

    \I__8735\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35303\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__35443\,
            I => \N__35296\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__35436\,
            I => \N__35296\
        );

    \I__8732\ : Span4Mux_v
    port map (
            O => \N__35433\,
            I => \N__35296\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__35430\,
            I => \N__35289\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__35427\,
            I => \N__35289\
        );

    \I__8729\ : Span4Mux_v
    port map (
            O => \N__35422\,
            I => \N__35289\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__35419\,
            I => \N__35284\
        );

    \I__8727\ : Span4Mux_v
    port map (
            O => \N__35416\,
            I => \N__35284\
        );

    \I__8726\ : Span4Mux_v
    port map (
            O => \N__35413\,
            I => \N__35279\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__35408\,
            I => \N__35279\
        );

    \I__8724\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35270\
        );

    \I__8723\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35270\
        );

    \I__8722\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35270\
        );

    \I__8721\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35270\
        );

    \I__8720\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35267\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__35398\,
            I => \N__35262\
        );

    \I__8718\ : Span4Mux_h
    port map (
            O => \N__35385\,
            I => \N__35262\
        );

    \I__8717\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35252\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__35381\,
            I => \N__35245\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__35378\,
            I => \N__35245\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__35373\,
            I => \N__35245\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__35368\,
            I => \N__35242\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__35363\,
            I => \N__35237\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__35358\,
            I => \N__35237\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35234\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__35350\,
            I => \N__35231\
        );

    \I__8708\ : InMux
    port map (
            O => \N__35349\,
            I => \N__35228\
        );

    \I__8707\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35225\
        );

    \I__8706\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35220\
        );

    \I__8705\ : InMux
    port map (
            O => \N__35346\,
            I => \N__35220\
        );

    \I__8704\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35211\
        );

    \I__8703\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35211\
        );

    \I__8702\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35211\
        );

    \I__8701\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35211\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__35339\,
            I => \N__35208\
        );

    \I__8699\ : Sp12to4
    port map (
            O => \N__35330\,
            I => \N__35205\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__35325\,
            I => \N__35196\
        );

    \I__8697\ : Sp12to4
    port map (
            O => \N__35322\,
            I => \N__35196\
        );

    \I__8696\ : Span12Mux_h
    port map (
            O => \N__35311\,
            I => \N__35196\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__35306\,
            I => \N__35196\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35185\
        );

    \I__8693\ : Span4Mux_v
    port map (
            O => \N__35296\,
            I => \N__35185\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__35289\,
            I => \N__35185\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__35284\,
            I => \N__35185\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__35279\,
            I => \N__35185\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35178\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35178\
        );

    \I__8687\ : Sp12to4
    port map (
            O => \N__35262\,
            I => \N__35178\
        );

    \I__8686\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35175\
        );

    \I__8685\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35170\
        );

    \I__8684\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35170\
        );

    \I__8683\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35163\
        );

    \I__8682\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35163\
        );

    \I__8681\ : InMux
    port map (
            O => \N__35256\,
            I => \N__35163\
        );

    \I__8680\ : InMux
    port map (
            O => \N__35255\,
            I => \N__35160\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__35252\,
            I => \N__35157\
        );

    \I__8678\ : Span4Mux_v
    port map (
            O => \N__35245\,
            I => \N__35154\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__35242\,
            I => \N__35145\
        );

    \I__8676\ : Span4Mux_s1_h
    port map (
            O => \N__35237\,
            I => \N__35145\
        );

    \I__8675\ : Span4Mux_v
    port map (
            O => \N__35234\,
            I => \N__35145\
        );

    \I__8674\ : Span4Mux_v
    port map (
            O => \N__35231\,
            I => \N__35145\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35132\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35132\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__35220\,
            I => \N__35132\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35132\
        );

    \I__8669\ : Span12Mux_h
    port map (
            O => \N__35208\,
            I => \N__35132\
        );

    \I__8668\ : Span12Mux_s4_h
    port map (
            O => \N__35205\,
            I => \N__35132\
        );

    \I__8667\ : Span12Mux_v
    port map (
            O => \N__35196\,
            I => \N__35129\
        );

    \I__8666\ : Sp12to4
    port map (
            O => \N__35185\,
            I => \N__35124\
        );

    \I__8665\ : Span12Mux_v
    port map (
            O => \N__35178\,
            I => \N__35124\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__35175\,
            I => rx_data_ready
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__35170\,
            I => rx_data_ready
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__35163\,
            I => rx_data_ready
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__35160\,
            I => rx_data_ready
        );

    \I__8660\ : Odrv4
    port map (
            O => \N__35157\,
            I => rx_data_ready
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__35154\,
            I => rx_data_ready
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__35145\,
            I => rx_data_ready
        );

    \I__8657\ : Odrv12
    port map (
            O => \N__35132\,
            I => rx_data_ready
        );

    \I__8656\ : Odrv12
    port map (
            O => \N__35129\,
            I => rx_data_ready
        );

    \I__8655\ : Odrv12
    port map (
            O => \N__35124\,
            I => rx_data_ready
        );

    \I__8654\ : CascadeMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__8653\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35096\
        );

    \I__8652\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__35096\,
            I => \N__35090\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__35087\
        );

    \I__8649\ : Span4Mux_v
    port map (
            O => \N__35090\,
            I => \N__35081\
        );

    \I__8648\ : Span4Mux_v
    port map (
            O => \N__35087\,
            I => \N__35081\
        );

    \I__8647\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35078\
        );

    \I__8646\ : Odrv4
    port map (
            O => \N__35081\,
            I => data_in_16_0
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__35078\,
            I => data_in_16_0
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__8643\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35066\
        );

    \I__8642\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35063\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35057\
        );

    \I__8639\ : Span4Mux_v
    port map (
            O => \N__35060\,
            I => \N__35052\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__35057\,
            I => \N__35052\
        );

    \I__8637\ : Span4Mux_h
    port map (
            O => \N__35052\,
            I => \N__35048\
        );

    \I__8636\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35045\
        );

    \I__8635\ : Odrv4
    port map (
            O => \N__35048\,
            I => data_in_15_0
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__35045\,
            I => data_in_15_0
        );

    \I__8633\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35031\
        );

    \I__8632\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35031\
        );

    \I__8631\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35031\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__8629\ : Span4Mux_h
    port map (
            O => \N__35028\,
            I => \N__35025\
        );

    \I__8628\ : Span4Mux_h
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__35022\,
            I => \c0.n5409\
        );

    \I__8626\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35015\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__35018\,
            I => \N__35009\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__35004\
        );

    \I__8623\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35001\
        );

    \I__8622\ : InMux
    port map (
            O => \N__35013\,
            I => \N__34998\
        );

    \I__8621\ : InMux
    port map (
            O => \N__35012\,
            I => \N__34993\
        );

    \I__8620\ : InMux
    port map (
            O => \N__35009\,
            I => \N__34993\
        );

    \I__8619\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34988\
        );

    \I__8618\ : InMux
    port map (
            O => \N__35007\,
            I => \N__34988\
        );

    \I__8617\ : Span4Mux_h
    port map (
            O => \N__35004\,
            I => \N__34983\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34983\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__34998\,
            I => data_out_11_1
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__34993\,
            I => data_out_11_1
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__34988\,
            I => data_out_11_1
        );

    \I__8612\ : Odrv4
    port map (
            O => \N__34983\,
            I => data_out_11_1
        );

    \I__8611\ : CascadeMux
    port map (
            O => \N__34974\,
            I => \c0.n5409_cascade_\
        );

    \I__8610\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34963\
        );

    \I__8609\ : InMux
    port map (
            O => \N__34970\,
            I => \N__34963\
        );

    \I__8608\ : CascadeMux
    port map (
            O => \N__34969\,
            I => \N__34958\
        );

    \I__8607\ : CascadeMux
    port map (
            O => \N__34968\,
            I => \N__34955\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34952\
        );

    \I__8605\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34949\
        );

    \I__8604\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34946\
        );

    \I__8603\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34940\
        );

    \I__8602\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34940\
        );

    \I__8601\ : Span4Mux_h
    port map (
            O => \N__34952\,
            I => \N__34937\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34932\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__34946\,
            I => \N__34932\
        );

    \I__8598\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34929\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34926\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__34937\,
            I => data_out_11_4
        );

    \I__8595\ : Odrv4
    port map (
            O => \N__34932\,
            I => data_out_11_4
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__34929\,
            I => data_out_11_4
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__34926\,
            I => data_out_11_4
        );

    \I__8592\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34914\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__8590\ : Span4Mux_h
    port map (
            O => \N__34911\,
            I => \N__34908\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__34908\,
            I => n4_adj_1978
        );

    \I__8588\ : CascadeMux
    port map (
            O => \N__34905\,
            I => \N__34902\
        );

    \I__8587\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__8585\ : Span4Mux_v
    port map (
            O => \N__34896\,
            I => \N__34893\
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__34893\,
            I => n4_adj_1983
        );

    \I__8583\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34887\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__34887\,
            I => n11
        );

    \I__8581\ : InMux
    port map (
            O => \N__34884\,
            I => n4724
        );

    \I__8580\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__34878\,
            I => n10
        );

    \I__8578\ : InMux
    port map (
            O => \N__34875\,
            I => \bfn_14_27_0_\
        );

    \I__8577\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__34869\,
            I => n9
        );

    \I__8575\ : InMux
    port map (
            O => \N__34866\,
            I => n4726
        );

    \I__8574\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__34860\,
            I => n8
        );

    \I__8572\ : InMux
    port map (
            O => \N__34857\,
            I => n4727
        );

    \I__8571\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__34851\,
            I => n7
        );

    \I__8569\ : InMux
    port map (
            O => \N__34848\,
            I => n4728
        );

    \I__8568\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__34842\,
            I => n6
        );

    \I__8566\ : InMux
    port map (
            O => \N__34839\,
            I => n4729
        );

    \I__8565\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34830\
        );

    \I__8564\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34830\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__8562\ : Span4Mux_v
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__34824\,
            I => \N__34820\
        );

    \I__8560\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34817\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__34820\,
            I => blink_counter_21
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__34817\,
            I => blink_counter_21
        );

    \I__8557\ : InMux
    port map (
            O => \N__34812\,
            I => n4730
        );

    \I__8556\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34803\
        );

    \I__8555\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34803\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__34800\,
            I => \N__34797\
        );

    \I__8552\ : Sp12to4
    port map (
            O => \N__34797\,
            I => \N__34793\
        );

    \I__8551\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34790\
        );

    \I__8550\ : Odrv12
    port map (
            O => \N__34793\,
            I => blink_counter_22
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__34790\,
            I => blink_counter_22
        );

    \I__8548\ : InMux
    port map (
            O => \N__34785\,
            I => n4731
        );

    \I__8547\ : InMux
    port map (
            O => \N__34782\,
            I => n4715
        );

    \I__8546\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__34776\,
            I => n19
        );

    \I__8544\ : InMux
    port map (
            O => \N__34773\,
            I => n4716
        );

    \I__8543\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34767\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__34767\,
            I => n18
        );

    \I__8541\ : InMux
    port map (
            O => \N__34764\,
            I => \bfn_14_26_0_\
        );

    \I__8540\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34758\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__34758\,
            I => n17
        );

    \I__8538\ : InMux
    port map (
            O => \N__34755\,
            I => n4718
        );

    \I__8537\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34749\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__34749\,
            I => n16
        );

    \I__8535\ : InMux
    port map (
            O => \N__34746\,
            I => n4719
        );

    \I__8534\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34740\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__34740\,
            I => n15
        );

    \I__8532\ : InMux
    port map (
            O => \N__34737\,
            I => n4720
        );

    \I__8531\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__34731\,
            I => n14
        );

    \I__8529\ : InMux
    port map (
            O => \N__34728\,
            I => n4721
        );

    \I__8528\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34722\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__34722\,
            I => n13
        );

    \I__8526\ : InMux
    port map (
            O => \N__34719\,
            I => n4722
        );

    \I__8525\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34713\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__34713\,
            I => n12
        );

    \I__8523\ : InMux
    port map (
            O => \N__34710\,
            I => n4723
        );

    \I__8522\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34702\
        );

    \I__8521\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34697\
        );

    \I__8520\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34697\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34691\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34688\
        );

    \I__8517\ : InMux
    port map (
            O => \N__34696\,
            I => \N__34683\
        );

    \I__8516\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34683\
        );

    \I__8515\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34679\
        );

    \I__8514\ : Span4Mux_v
    port map (
            O => \N__34691\,
            I => \N__34676\
        );

    \I__8513\ : Span4Mux_v
    port map (
            O => \N__34688\,
            I => \N__34671\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__34683\,
            I => \N__34671\
        );

    \I__8511\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34668\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__34679\,
            I => data_out_11_5
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__34676\,
            I => data_out_11_5
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__34671\,
            I => data_out_11_5
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__34668\,
            I => data_out_11_5
        );

    \I__8506\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34654\
        );

    \I__8505\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34651\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34646\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__34654\,
            I => \N__34643\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__34651\,
            I => \N__34638\
        );

    \I__8501\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34635\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34632\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__34646\,
            I => \N__34629\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__34643\,
            I => \N__34626\
        );

    \I__8497\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34621\
        );

    \I__8496\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34621\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__34638\,
            I => \N__34618\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__34635\,
            I => \N__34613\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__34632\,
            I => \N__34613\
        );

    \I__8492\ : Odrv12
    port map (
            O => \N__34629\,
            I => data_out_10_6
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__34626\,
            I => data_out_10_6
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__34621\,
            I => data_out_10_6
        );

    \I__8489\ : Odrv4
    port map (
            O => \N__34618\,
            I => data_out_10_6
        );

    \I__8488\ : Odrv4
    port map (
            O => \N__34613\,
            I => data_out_10_6
        );

    \I__8487\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34599\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34596\
        );

    \I__8485\ : Odrv12
    port map (
            O => \N__34596\,
            I => n4_adj_1976
        );

    \I__8484\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34590\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__34590\,
            I => n26
        );

    \I__8482\ : InMux
    port map (
            O => \N__34587\,
            I => \bfn_14_25_0_\
        );

    \I__8481\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34581\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__34581\,
            I => n25
        );

    \I__8479\ : InMux
    port map (
            O => \N__34578\,
            I => n4710
        );

    \I__8478\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34572\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__34572\,
            I => n24
        );

    \I__8476\ : InMux
    port map (
            O => \N__34569\,
            I => n4711
        );

    \I__8475\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34563\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__34563\,
            I => n23
        );

    \I__8473\ : InMux
    port map (
            O => \N__34560\,
            I => n4712
        );

    \I__8472\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34554\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__34554\,
            I => n22
        );

    \I__8470\ : InMux
    port map (
            O => \N__34551\,
            I => n4713
        );

    \I__8469\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__34545\,
            I => n21
        );

    \I__8467\ : InMux
    port map (
            O => \N__34542\,
            I => n4714
        );

    \I__8466\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__34536\,
            I => n20
        );

    \I__8464\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34528\
        );

    \I__8463\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34525\
        );

    \I__8462\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34522\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__34528\,
            I => \N__34515\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__34525\,
            I => \N__34512\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__34522\,
            I => \N__34509\
        );

    \I__8458\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34500\
        );

    \I__8457\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34500\
        );

    \I__8456\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34500\
        );

    \I__8455\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34500\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__34515\,
            I => data_out_11_7
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__34512\,
            I => data_out_11_7
        );

    \I__8452\ : Odrv4
    port map (
            O => \N__34509\,
            I => data_out_11_7
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__34500\,
            I => data_out_11_7
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__34491\,
            I => \N__34488\
        );

    \I__8449\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34485\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__34485\,
            I => \N__34482\
        );

    \I__8447\ : Span4Mux_h
    port map (
            O => \N__34482\,
            I => \N__34479\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__34479\,
            I => \N__34474\
        );

    \I__8445\ : InMux
    port map (
            O => \N__34478\,
            I => \N__34471\
        );

    \I__8444\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34468\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__34474\,
            I => data_in_13_5
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__34471\,
            I => data_in_13_5
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__34468\,
            I => data_in_13_5
        );

    \I__8440\ : CascadeMux
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__8439\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34454\
        );

    \I__8438\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34451\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34448\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__34451\,
            I => \N__34445\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__34448\,
            I => \N__34439\
        );

    \I__8434\ : Span4Mux_h
    port map (
            O => \N__34445\,
            I => \N__34439\
        );

    \I__8433\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34436\
        );

    \I__8432\ : Odrv4
    port map (
            O => \N__34439\,
            I => data_in_12_5
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__34436\,
            I => data_in_12_5
        );

    \I__8430\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34426\
        );

    \I__8429\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34423\
        );

    \I__8428\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34420\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34412\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__34423\,
            I => \N__34412\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34412\
        );

    \I__8424\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34408\
        );

    \I__8423\ : Span4Mux_v
    port map (
            O => \N__34412\,
            I => \N__34405\
        );

    \I__8422\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34402\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__34408\,
            I => data_out_10_5
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__34405\,
            I => data_out_10_5
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__34402\,
            I => data_out_10_5
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__34395\,
            I => \N__34392\
        );

    \I__8417\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__8415\ : Odrv4
    port map (
            O => \N__34386\,
            I => \c0.n9_adj_1911\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__34383\,
            I => \N__34376\
        );

    \I__8413\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34370\
        );

    \I__8412\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34370\
        );

    \I__8411\ : InMux
    port map (
            O => \N__34380\,
            I => \N__34367\
        );

    \I__8410\ : InMux
    port map (
            O => \N__34379\,
            I => \N__34364\
        );

    \I__8409\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34361\
        );

    \I__8408\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34358\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__34370\,
            I => \N__34355\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__34367\,
            I => \N__34352\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__34364\,
            I => \N__34349\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__34361\,
            I => \N__34342\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__34358\,
            I => \N__34342\
        );

    \I__8402\ : Span4Mux_h
    port map (
            O => \N__34355\,
            I => \N__34342\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__34352\,
            I => \N__34339\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__34349\,
            I => data_out_10_0
        );

    \I__8399\ : Odrv4
    port map (
            O => \N__34342\,
            I => data_out_10_0
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__34339\,
            I => data_out_10_0
        );

    \I__8397\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34316\
        );

    \I__8396\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34309\
        );

    \I__8395\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34309\
        );

    \I__8394\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34309\
        );

    \I__8393\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34304\
        );

    \I__8392\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34304\
        );

    \I__8391\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34296\
        );

    \I__8390\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34296\
        );

    \I__8389\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34291\
        );

    \I__8388\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34291\
        );

    \I__8387\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34286\
        );

    \I__8386\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34286\
        );

    \I__8385\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34283\
        );

    \I__8384\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34280\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34271\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__34309\,
            I => \N__34271\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__34304\,
            I => \N__34271\
        );

    \I__8380\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34262\
        );

    \I__8379\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34262\
        );

    \I__8378\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34262\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34257\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__34291\,
            I => \N__34257\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__34286\,
            I => \N__34250\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__34283\,
            I => \N__34250\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34250\
        );

    \I__8372\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34247\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__34278\,
            I => \N__34244\
        );

    \I__8370\ : Span4Mux_v
    port map (
            O => \N__34271\,
            I => \N__34241\
        );

    \I__8369\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34238\
        );

    \I__8368\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34235\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34226\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__34257\,
            I => \N__34226\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__34250\,
            I => \N__34226\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34226\
        );

    \I__8363\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34223\
        );

    \I__8362\ : Odrv4
    port map (
            O => \N__34241\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__34238\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__34235\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__34226\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__34223\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8357\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34208\
        );

    \I__8356\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34201\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34198\
        );

    \I__8354\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34188\
        );

    \I__8353\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34188\
        );

    \I__8352\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34188\
        );

    \I__8351\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34188\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__34201\,
            I => \N__34183\
        );

    \I__8349\ : Span4Mux_h
    port map (
            O => \N__34198\,
            I => \N__34180\
        );

    \I__8348\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34177\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__34188\,
            I => \N__34174\
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__34187\,
            I => \N__34168\
        );

    \I__8345\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34165\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__34183\,
            I => \N__34162\
        );

    \I__8343\ : Span4Mux_h
    port map (
            O => \N__34180\,
            I => \N__34155\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__34177\,
            I => \N__34155\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__34174\,
            I => \N__34155\
        );

    \I__8340\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34148\
        );

    \I__8339\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34148\
        );

    \I__8338\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34148\
        );

    \I__8337\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34145\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__34165\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__34162\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8334\ : Odrv4
    port map (
            O => \N__34155\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__34148\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__34145\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8331\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34123\
        );

    \I__8330\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34123\
        );

    \I__8329\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34123\
        );

    \I__8328\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34118\
        );

    \I__8327\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34118\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__34123\,
            I => \N__34109\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34118\,
            I => \N__34109\
        );

    \I__8324\ : InMux
    port map (
            O => \N__34117\,
            I => \N__34105\
        );

    \I__8323\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34098\
        );

    \I__8322\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34098\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34098\
        );

    \I__8320\ : Span4Mux_h
    port map (
            O => \N__34109\,
            I => \N__34095\
        );

    \I__8319\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34092\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__34105\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__34098\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__34095\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__34092\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__34083\,
            I => \c0.n9_adj_1891_cascade_\
        );

    \I__8313\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34076\
        );

    \I__8312\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34073\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__34076\,
            I => \N__34061\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__34073\,
            I => \N__34061\
        );

    \I__8309\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34050\
        );

    \I__8308\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34050\
        );

    \I__8307\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34050\
        );

    \I__8306\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34043\
        );

    \I__8305\ : InMux
    port map (
            O => \N__34068\,
            I => \N__34043\
        );

    \I__8304\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34043\
        );

    \I__8303\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34040\
        );

    \I__8302\ : Span4Mux_v
    port map (
            O => \N__34061\,
            I => \N__34037\
        );

    \I__8301\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34031\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34031\
        );

    \I__8299\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34026\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34057\,
            I => \N__34026\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__34050\,
            I => \N__34023\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34018\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34018\
        );

    \I__8294\ : Span4Mux_h
    port map (
            O => \N__34037\,
            I => \N__34014\
        );

    \I__8293\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34011\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34008\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__34026\,
            I => \N__34003\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__34023\,
            I => \N__34003\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__34018\,
            I => \N__34000\
        );

    \I__8288\ : InMux
    port map (
            O => \N__34017\,
            I => \N__33997\
        );

    \I__8287\ : Odrv4
    port map (
            O => \N__34014\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__34011\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8285\ : Odrv12
    port map (
            O => \N__34008\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8284\ : Odrv4
    port map (
            O => \N__34003\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__34000\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__33997\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8281\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__8279\ : Span4Mux_v
    port map (
            O => \N__33978\,
            I => \N__33975\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__33975\,
            I => \c0.n15_adj_1893\
        );

    \I__8277\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33968\
        );

    \I__8276\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33964\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__33968\,
            I => \N__33961\
        );

    \I__8274\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33958\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__33964\,
            I => n5421
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__33961\,
            I => n5421
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__33958\,
            I => n5421
        );

    \I__8270\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33947\
        );

    \I__8269\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33944\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__33947\,
            I => \N__33941\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__33944\,
            I => data_out_18_1
        );

    \I__8266\ : Odrv4
    port map (
            O => \N__33941\,
            I => data_out_18_1
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__8264\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33927\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__33927\,
            I => \N__33923\
        );

    \I__8261\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33920\
        );

    \I__8260\ : Sp12to4
    port map (
            O => \N__33923\,
            I => \N__33917\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__33920\,
            I => data_out_19_3
        );

    \I__8258\ : Odrv12
    port map (
            O => \N__33917\,
            I => data_out_19_3
        );

    \I__8257\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__33909\,
            I => \c0.n5837\
        );

    \I__8255\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33902\
        );

    \I__8254\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33899\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__33902\,
            I => \r_Tx_Data_5\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__33899\,
            I => \r_Tx_Data_5\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__33894\,
            I => \N__33889\
        );

    \I__8250\ : CascadeMux
    port map (
            O => \N__33893\,
            I => \N__33885\
        );

    \I__8249\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33878\
        );

    \I__8248\ : InMux
    port map (
            O => \N__33889\,
            I => \N__33878\
        );

    \I__8247\ : InMux
    port map (
            O => \N__33888\,
            I => \N__33873\
        );

    \I__8246\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33873\
        );

    \I__8245\ : CascadeMux
    port map (
            O => \N__33884\,
            I => \N__33870\
        );

    \I__8244\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33865\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__33878\,
            I => \N__33862\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__33873\,
            I => \N__33859\
        );

    \I__8241\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33854\
        );

    \I__8240\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33854\
        );

    \I__8239\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33851\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33848\
        );

    \I__8237\ : Span4Mux_h
    port map (
            O => \N__33862\,
            I => \N__33843\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__33859\,
            I => \N__33843\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__33854\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__33851\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__33848\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__33843\,
            I => \c0.tx.r_Bit_Index_1\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__33834\,
            I => \N__33830\
        );

    \I__8230\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33827\
        );

    \I__8229\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33824\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33819\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33819\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__33819\,
            I => \r_Tx_Data_4\
        );

    \I__8225\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__8222\ : Odrv4
    port map (
            O => \N__33807\,
            I => \c0.tx.n6285\
        );

    \I__8221\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33801\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__33801\,
            I => \c0.tx.n6288\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__8218\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33792\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33789\
        );

    \I__8216\ : Span4Mux_h
    port map (
            O => \N__33789\,
            I => \N__33786\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__33786\,
            I => n5415
        );

    \I__8214\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33777\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__33782\,
            I => \N__33774\
        );

    \I__8212\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33769\
        );

    \I__8211\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33769\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33766\
        );

    \I__8209\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33763\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__33769\,
            I => \N__33760\
        );

    \I__8207\ : Odrv12
    port map (
            O => \N__33766\,
            I => \c0.n1251\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__33763\,
            I => \c0.n1251\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__33760\,
            I => \c0.n1251\
        );

    \I__8204\ : CascadeMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__8203\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33747\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__33747\,
            I => \c0.n5845\
        );

    \I__8201\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33733\
        );

    \I__8199\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33724\
        );

    \I__8198\ : InMux
    port map (
            O => \N__33739\,
            I => \N__33724\
        );

    \I__8197\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33724\
        );

    \I__8196\ : InMux
    port map (
            O => \N__33737\,
            I => \N__33724\
        );

    \I__8195\ : InMux
    port map (
            O => \N__33736\,
            I => \N__33719\
        );

    \I__8194\ : Span4Mux_h
    port map (
            O => \N__33733\,
            I => \N__33714\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__33724\,
            I => \N__33714\
        );

    \I__8192\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33710\
        );

    \I__8191\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33707\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33704\
        );

    \I__8189\ : Span4Mux_v
    port map (
            O => \N__33714\,
            I => \N__33701\
        );

    \I__8188\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33698\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__33710\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__33707\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8185\ : Odrv4
    port map (
            O => \N__33704\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__33701\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__33698\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8182\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__33684\,
            I => \tx_data_1_N_keep\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__33681\,
            I => \c0.n9_adj_1906_cascade_\
        );

    \I__8179\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33675\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__33675\,
            I => \N__33672\
        );

    \I__8177\ : Odrv4
    port map (
            O => \N__33672\,
            I => \c0.n15_adj_1909\
        );

    \I__8176\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33661\
        );

    \I__8174\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33658\
        );

    \I__8173\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33652\
        );

    \I__8172\ : Span12Mux_v
    port map (
            O => \N__33661\,
            I => \N__33647\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__33658\,
            I => \N__33647\
        );

    \I__8170\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33640\
        );

    \I__8169\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33640\
        );

    \I__8168\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33640\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__33652\,
            I => data_out_10_4
        );

    \I__8166\ : Odrv12
    port map (
            O => \N__33647\,
            I => data_out_10_4
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__33640\,
            I => data_out_10_4
        );

    \I__8164\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__8162\ : Odrv12
    port map (
            O => \N__33627\,
            I => \c0.n2293\
        );

    \I__8161\ : InMux
    port map (
            O => \N__33624\,
            I => \N__33621\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__33621\,
            I => \N__33618\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__33615\,
            I => n4_adj_1996
        );

    \I__8157\ : CascadeMux
    port map (
            O => \N__33612\,
            I => \N__33606\
        );

    \I__8156\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33602\
        );

    \I__8155\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33599\
        );

    \I__8154\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33595\
        );

    \I__8153\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33592\
        );

    \I__8152\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33589\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__33602\,
            I => \N__33586\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33583\
        );

    \I__8149\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33580\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__33595\,
            I => \N__33577\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33572\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33572\
        );

    \I__8145\ : Span4Mux_v
    port map (
            O => \N__33586\,
            I => \N__33563\
        );

    \I__8144\ : Span4Mux_v
    port map (
            O => \N__33583\,
            I => \N__33563\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33563\
        );

    \I__8142\ : Span4Mux_v
    port map (
            O => \N__33577\,
            I => \N__33558\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__33572\,
            I => \N__33558\
        );

    \I__8140\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33555\
        );

    \I__8139\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33552\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__33563\,
            I => \N__33549\
        );

    \I__8137\ : Sp12to4
    port map (
            O => \N__33558\,
            I => \N__33544\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__33555\,
            I => \N__33544\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__33552\,
            I => \N__33541\
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__33549\,
            I => n1519
        );

    \I__8133\ : Odrv12
    port map (
            O => \N__33544\,
            I => n1519
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__33541\,
            I => n1519
        );

    \I__8131\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__33531\,
            I => \tx_data_5_N_keep\
        );

    \I__8129\ : CascadeMux
    port map (
            O => \N__33528\,
            I => \c0.n95_cascade_\
        );

    \I__8128\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33519\
        );

    \I__8127\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33519\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__33519\,
            I => \c0.n106\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__8124\ : InMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__8122\ : Odrv12
    port map (
            O => \N__33507\,
            I => n4_adj_1981
        );

    \I__8121\ : CascadeMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__8120\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33498\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__33495\,
            I => n7_adj_1988
        );

    \I__8117\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33483\
        );

    \I__8116\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33483\
        );

    \I__8115\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33476\
        );

    \I__8114\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33476\
        );

    \I__8113\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33476\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__33483\,
            I => \c0.n15\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__33476\,
            I => \c0.n15\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__33471\,
            I => \N__33468\
        );

    \I__8109\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33461\
        );

    \I__8108\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33461\
        );

    \I__8107\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33458\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33451\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33451\
        );

    \I__8104\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33448\
        );

    \I__8103\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33445\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__33451\,
            I => \c0.n81_adj_1872\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__33448\,
            I => \c0.n81_adj_1872\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__33445\,
            I => \c0.n81_adj_1872\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__33438\,
            I => \N__33433\
        );

    \I__8098\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33429\
        );

    \I__8097\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33422\
        );

    \I__8096\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33422\
        );

    \I__8095\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33422\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__33429\,
            I => \c0.tx_transmit_N_568_4\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__33422\,
            I => \c0.tx_transmit_N_568_4\
        );

    \I__8092\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33411\
        );

    \I__8091\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33411\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__33411\,
            I => \c0.tx_transmit_N_568_2\
        );

    \I__8089\ : CascadeMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__8088\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33402\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__8086\ : Odrv12
    port map (
            O => \N__33399\,
            I => \c0.n5833\
        );

    \I__8085\ : CascadeMux
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__8084\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33390\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__8082\ : Span4Mux_h
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__33384\,
            I => \c0.n31_adj_1912\
        );

    \I__8080\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33378\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__33378\,
            I => \c0.n989\
        );

    \I__8078\ : InMux
    port map (
            O => \N__33375\,
            I => \c0.n4703\
        );

    \I__8077\ : InMux
    port map (
            O => \N__33372\,
            I => \c0.n4704\
        );

    \I__8076\ : InMux
    port map (
            O => \N__33369\,
            I => \c0.n4705\
        );

    \I__8075\ : InMux
    port map (
            O => \N__33366\,
            I => \c0.n4706\
        );

    \I__8074\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33360\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__33360\,
            I => \c0.byte_transmit_counter_5\
        );

    \I__8072\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33351\
        );

    \I__8071\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33351\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__33351\,
            I => \c0.tx_transmit_N_568_5\
        );

    \I__8069\ : InMux
    port map (
            O => \N__33348\,
            I => \c0.n4707\
        );

    \I__8068\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33342\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33339\
        );

    \I__8066\ : Odrv4
    port map (
            O => \N__33339\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__8065\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33333\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33329\
        );

    \I__8063\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33326\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__33329\,
            I => \c0.tx_transmit_N_568_6\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__33326\,
            I => \c0.tx_transmit_N_568_6\
        );

    \I__8060\ : InMux
    port map (
            O => \N__33321\,
            I => \c0.n4708\
        );

    \I__8059\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__33315\,
            I => \N__33312\
        );

    \I__8057\ : Odrv4
    port map (
            O => \N__33312\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__8056\ : InMux
    port map (
            O => \N__33309\,
            I => \c0.n4709\
        );

    \I__8055\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33299\
        );

    \I__8053\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33296\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__33299\,
            I => \c0.tx_transmit_N_568_7\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__33296\,
            I => \c0.tx_transmit_N_568_7\
        );

    \I__8050\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33285\
        );

    \I__8049\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33285\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__33285\,
            I => \c0.tx_transmit_N_568_3\
        );

    \I__8047\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__33279\,
            I => \c0.n95\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__33276\,
            I => \N__33264\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33258\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__33274\,
            I => \N__33255\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__33273\,
            I => \N__33247\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__33272\,
            I => \N__33235\
        );

    \I__8040\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33220\
        );

    \I__8039\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33220\
        );

    \I__8038\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33220\
        );

    \I__8037\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33212\
        );

    \I__8036\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33212\
        );

    \I__8035\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33203\
        );

    \I__8034\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33203\
        );

    \I__8033\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33203\
        );

    \I__8032\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33203\
        );

    \I__8031\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33198\
        );

    \I__8030\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33198\
        );

    \I__8029\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33191\
        );

    \I__8028\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33191\
        );

    \I__8027\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33191\
        );

    \I__8026\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33186\
        );

    \I__8025\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33186\
        );

    \I__8024\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33183\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33180\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__33245\,
            I => \N__33177\
        );

    \I__8021\ : CascadeMux
    port map (
            O => \N__33244\,
            I => \N__33170\
        );

    \I__8020\ : CascadeMux
    port map (
            O => \N__33243\,
            I => \N__33167\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__33242\,
            I => \N__33160\
        );

    \I__8018\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33144\
        );

    \I__8017\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33144\
        );

    \I__8016\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33144\
        );

    \I__8015\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33144\
        );

    \I__8014\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33139\
        );

    \I__8013\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33139\
        );

    \I__8012\ : CascadeMux
    port map (
            O => \N__33233\,
            I => \N__33132\
        );

    \I__8011\ : CascadeMux
    port map (
            O => \N__33232\,
            I => \N__33126\
        );

    \I__8010\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33112\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33112\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__33229\,
            I => \N__33109\
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__33228\,
            I => \N__33099\
        );

    \I__8006\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33091\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33088\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__33219\,
            I => \N__33078\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__33218\,
            I => \N__33071\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__33217\,
            I => \N__33065\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33062\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__33203\,
            I => \N__33055\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__33198\,
            I => \N__33055\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33055\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33050\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33050\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__33180\,
            I => \N__33047\
        );

    \I__7994\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33038\
        );

    \I__7993\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33038\
        );

    \I__7992\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33038\
        );

    \I__7991\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33038\
        );

    \I__7990\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33027\
        );

    \I__7989\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33027\
        );

    \I__7988\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33027\
        );

    \I__7987\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33027\
        );

    \I__7986\ : InMux
    port map (
            O => \N__33165\,
            I => \N__33027\
        );

    \I__7985\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33015\
        );

    \I__7984\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33015\
        );

    \I__7983\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33015\
        );

    \I__7982\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33015\
        );

    \I__7981\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33015\
        );

    \I__7980\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33010\
        );

    \I__7979\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33010\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__33155\,
            I => \N__33007\
        );

    \I__7977\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33000\
        );

    \I__7976\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33000\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__33144\,
            I => \N__32995\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__33139\,
            I => \N__32995\
        );

    \I__7973\ : InMux
    port map (
            O => \N__33138\,
            I => \N__32979\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__33137\,
            I => \N__32974\
        );

    \I__7971\ : CascadeMux
    port map (
            O => \N__33136\,
            I => \N__32971\
        );

    \I__7970\ : InMux
    port map (
            O => \N__33135\,
            I => \N__32958\
        );

    \I__7969\ : InMux
    port map (
            O => \N__33132\,
            I => \N__32958\
        );

    \I__7968\ : InMux
    port map (
            O => \N__33131\,
            I => \N__32958\
        );

    \I__7967\ : InMux
    port map (
            O => \N__33130\,
            I => \N__32958\
        );

    \I__7966\ : InMux
    port map (
            O => \N__33129\,
            I => \N__32958\
        );

    \I__7965\ : InMux
    port map (
            O => \N__33126\,
            I => \N__32953\
        );

    \I__7964\ : InMux
    port map (
            O => \N__33125\,
            I => \N__32953\
        );

    \I__7963\ : InMux
    port map (
            O => \N__33124\,
            I => \N__32944\
        );

    \I__7962\ : InMux
    port map (
            O => \N__33123\,
            I => \N__32944\
        );

    \I__7961\ : InMux
    port map (
            O => \N__33122\,
            I => \N__32944\
        );

    \I__7960\ : InMux
    port map (
            O => \N__33121\,
            I => \N__32944\
        );

    \I__7959\ : InMux
    port map (
            O => \N__33120\,
            I => \N__32935\
        );

    \I__7958\ : InMux
    port map (
            O => \N__33119\,
            I => \N__32935\
        );

    \I__7957\ : InMux
    port map (
            O => \N__33118\,
            I => \N__32935\
        );

    \I__7956\ : InMux
    port map (
            O => \N__33117\,
            I => \N__32935\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__32932\
        );

    \I__7954\ : InMux
    port map (
            O => \N__33109\,
            I => \N__32925\
        );

    \I__7953\ : InMux
    port map (
            O => \N__33108\,
            I => \N__32925\
        );

    \I__7952\ : InMux
    port map (
            O => \N__33107\,
            I => \N__32925\
        );

    \I__7951\ : InMux
    port map (
            O => \N__33106\,
            I => \N__32920\
        );

    \I__7950\ : InMux
    port map (
            O => \N__33105\,
            I => \N__32920\
        );

    \I__7949\ : InMux
    port map (
            O => \N__33104\,
            I => \N__32917\
        );

    \I__7948\ : InMux
    port map (
            O => \N__33103\,
            I => \N__32913\
        );

    \I__7947\ : InMux
    port map (
            O => \N__33102\,
            I => \N__32910\
        );

    \I__7946\ : InMux
    port map (
            O => \N__33099\,
            I => \N__32905\
        );

    \I__7945\ : InMux
    port map (
            O => \N__33098\,
            I => \N__32905\
        );

    \I__7944\ : InMux
    port map (
            O => \N__33097\,
            I => \N__32896\
        );

    \I__7943\ : InMux
    port map (
            O => \N__33096\,
            I => \N__32896\
        );

    \I__7942\ : InMux
    port map (
            O => \N__33095\,
            I => \N__32896\
        );

    \I__7941\ : InMux
    port map (
            O => \N__33094\,
            I => \N__32896\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__33091\,
            I => \N__32891\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__33088\,
            I => \N__32888\
        );

    \I__7938\ : InMux
    port map (
            O => \N__33087\,
            I => \N__32881\
        );

    \I__7937\ : InMux
    port map (
            O => \N__33086\,
            I => \N__32881\
        );

    \I__7936\ : InMux
    port map (
            O => \N__33085\,
            I => \N__32881\
        );

    \I__7935\ : InMux
    port map (
            O => \N__33084\,
            I => \N__32878\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33083\,
            I => \N__32875\
        );

    \I__7933\ : InMux
    port map (
            O => \N__33082\,
            I => \N__32870\
        );

    \I__7932\ : InMux
    port map (
            O => \N__33081\,
            I => \N__32870\
        );

    \I__7931\ : InMux
    port map (
            O => \N__33078\,
            I => \N__32865\
        );

    \I__7930\ : InMux
    port map (
            O => \N__33077\,
            I => \N__32862\
        );

    \I__7929\ : InMux
    port map (
            O => \N__33076\,
            I => \N__32853\
        );

    \I__7928\ : InMux
    port map (
            O => \N__33075\,
            I => \N__32853\
        );

    \I__7927\ : InMux
    port map (
            O => \N__33074\,
            I => \N__32853\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33071\,
            I => \N__32848\
        );

    \I__7925\ : InMux
    port map (
            O => \N__33070\,
            I => \N__32848\
        );

    \I__7924\ : CascadeMux
    port map (
            O => \N__33069\,
            I => \N__32843\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__33068\,
            I => \N__32840\
        );

    \I__7922\ : InMux
    port map (
            O => \N__33065\,
            I => \N__32835\
        );

    \I__7921\ : Span4Mux_v
    port map (
            O => \N__33062\,
            I => \N__32824\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__33055\,
            I => \N__32824\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__33050\,
            I => \N__32824\
        );

    \I__7918\ : Span4Mux_v
    port map (
            O => \N__33047\,
            I => \N__32824\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__32824\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__33027\,
            I => \N__32821\
        );

    \I__7915\ : InMux
    port map (
            O => \N__33026\,
            I => \N__32818\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__32813\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__33010\,
            I => \N__32813\
        );

    \I__7912\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32808\
        );

    \I__7911\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32808\
        );

    \I__7910\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32801\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32798\
        );

    \I__7908\ : Span4Mux_h
    port map (
            O => \N__32995\,
            I => \N__32795\
        );

    \I__7907\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32784\
        );

    \I__7906\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32784\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32784\
        );

    \I__7904\ : InMux
    port map (
            O => \N__32991\,
            I => \N__32784\
        );

    \I__7903\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32784\
        );

    \I__7902\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32781\
        );

    \I__7901\ : CascadeMux
    port map (
            O => \N__32988\,
            I => \N__32774\
        );

    \I__7900\ : CascadeMux
    port map (
            O => \N__32987\,
            I => \N__32770\
        );

    \I__7899\ : CascadeMux
    port map (
            O => \N__32986\,
            I => \N__32764\
        );

    \I__7898\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32747\
        );

    \I__7897\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32747\
        );

    \I__7896\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32747\
        );

    \I__7895\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32747\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32744\
        );

    \I__7893\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32739\
        );

    \I__7892\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32739\
        );

    \I__7891\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32734\
        );

    \I__7890\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32734\
        );

    \I__7889\ : InMux
    port map (
            O => \N__32970\,
            I => \N__32729\
        );

    \I__7888\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32729\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32726\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__32953\,
            I => \N__32723\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__32944\,
            I => \N__32718\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32718\
        );

    \I__7883\ : Span4Mux_v
    port map (
            O => \N__32932\,
            I => \N__32709\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32709\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32709\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32709\
        );

    \I__7879\ : CascadeMux
    port map (
            O => \N__32916\,
            I => \N__32706\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32695\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__32910\,
            I => \N__32695\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32695\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__32896\,
            I => \N__32695\
        );

    \I__7874\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32690\
        );

    \I__7873\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32690\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__32891\,
            I => \N__32681\
        );

    \I__7871\ : Span4Mux_v
    port map (
            O => \N__32888\,
            I => \N__32681\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32681\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32681\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32676\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__32870\,
            I => \N__32676\
        );

    \I__7866\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32671\
        );

    \I__7865\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32671\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32666\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32666\
        );

    \I__7862\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32661\
        );

    \I__7861\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32661\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32656\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32656\
        );

    \I__7858\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32649\
        );

    \I__7857\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32649\
        );

    \I__7856\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32649\
        );

    \I__7855\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32644\
        );

    \I__7854\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32644\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__32838\,
            I => \N__32640\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32632\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__32824\,
            I => \N__32632\
        );

    \I__7850\ : Span4Mux_h
    port map (
            O => \N__32821\,
            I => \N__32623\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__32818\,
            I => \N__32623\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__32813\,
            I => \N__32623\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__32808\,
            I => \N__32623\
        );

    \I__7846\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32614\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32614\
        );

    \I__7844\ : InMux
    port map (
            O => \N__32805\,
            I => \N__32614\
        );

    \I__7843\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32614\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32603\
        );

    \I__7841\ : Span4Mux_v
    port map (
            O => \N__32798\,
            I => \N__32603\
        );

    \I__7840\ : Span4Mux_h
    port map (
            O => \N__32795\,
            I => \N__32603\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32603\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32603\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__32780\,
            I => \N__32599\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__32779\,
            I => \N__32595\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__32778\,
            I => \N__32592\
        );

    \I__7834\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32582\
        );

    \I__7833\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32582\
        );

    \I__7832\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32575\
        );

    \I__7831\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32575\
        );

    \I__7830\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32575\
        );

    \I__7829\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32572\
        );

    \I__7828\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32563\
        );

    \I__7827\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32563\
        );

    \I__7826\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32563\
        );

    \I__7825\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32563\
        );

    \I__7824\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32554\
        );

    \I__7823\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32554\
        );

    \I__7822\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32554\
        );

    \I__7821\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32554\
        );

    \I__7820\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32549\
        );

    \I__7819\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32549\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__32747\,
            I => \N__32542\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32542\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__32739\,
            I => \N__32542\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__32734\,
            I => \N__32531\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32531\
        );

    \I__7813\ : Span4Mux_v
    port map (
            O => \N__32726\,
            I => \N__32531\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__32723\,
            I => \N__32531\
        );

    \I__7811\ : Span4Mux_v
    port map (
            O => \N__32718\,
            I => \N__32531\
        );

    \I__7810\ : Span4Mux_v
    port map (
            O => \N__32709\,
            I => \N__32528\
        );

    \I__7809\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32521\
        );

    \I__7808\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32521\
        );

    \I__7807\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32521\
        );

    \I__7806\ : Span4Mux_h
    port map (
            O => \N__32695\,
            I => \N__32516\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32516\
        );

    \I__7804\ : Span4Mux_h
    port map (
            O => \N__32681\,
            I => \N__32505\
        );

    \I__7803\ : Span4Mux_h
    port map (
            O => \N__32676\,
            I => \N__32505\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__32671\,
            I => \N__32505\
        );

    \I__7801\ : Span4Mux_v
    port map (
            O => \N__32666\,
            I => \N__32505\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32505\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__32656\,
            I => \N__32502\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__32649\,
            I => \N__32497\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__32644\,
            I => \N__32497\
        );

    \I__7796\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32494\
        );

    \I__7795\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32485\
        );

    \I__7794\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32485\
        );

    \I__7793\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32485\
        );

    \I__7792\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32485\
        );

    \I__7791\ : Span4Mux_s1_h
    port map (
            O => \N__32632\,
            I => \N__32480\
        );

    \I__7790\ : Span4Mux_h
    port map (
            O => \N__32623\,
            I => \N__32480\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__32614\,
            I => \N__32475\
        );

    \I__7788\ : Span4Mux_h
    port map (
            O => \N__32603\,
            I => \N__32475\
        );

    \I__7787\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32469\
        );

    \I__7786\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32469\
        );

    \I__7785\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32462\
        );

    \I__7784\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32462\
        );

    \I__7783\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32462\
        );

    \I__7782\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32459\
        );

    \I__7781\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32454\
        );

    \I__7780\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32454\
        );

    \I__7779\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32449\
        );

    \I__7778\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32449\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__32582\,
            I => \N__32444\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32444\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32439\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__32563\,
            I => \N__32439\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32434\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32429\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__32542\,
            I => \N__32429\
        );

    \I__7770\ : Span4Mux_v
    port map (
            O => \N__32531\,
            I => \N__32426\
        );

    \I__7769\ : Span4Mux_v
    port map (
            O => \N__32528\,
            I => \N__32423\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32420\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__32516\,
            I => \N__32417\
        );

    \I__7766\ : Span4Mux_v
    port map (
            O => \N__32505\,
            I => \N__32414\
        );

    \I__7765\ : Span4Mux_v
    port map (
            O => \N__32502\,
            I => \N__32411\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__32497\,
            I => \N__32400\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32400\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32400\
        );

    \I__7761\ : Span4Mux_v
    port map (
            O => \N__32480\,
            I => \N__32400\
        );

    \I__7760\ : Span4Mux_h
    port map (
            O => \N__32475\,
            I => \N__32400\
        );

    \I__7759\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32397\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__32469\,
            I => \N__32394\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__32462\,
            I => \N__32391\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__32459\,
            I => \N__32380\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32380\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__32449\,
            I => \N__32380\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__32444\,
            I => \N__32380\
        );

    \I__7752\ : Span4Mux_v
    port map (
            O => \N__32439\,
            I => \N__32380\
        );

    \I__7751\ : CascadeMux
    port map (
            O => \N__32438\,
            I => \N__32376\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__32437\,
            I => \N__32373\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__32434\,
            I => \N__32363\
        );

    \I__7748\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32363\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__32426\,
            I => \N__32363\
        );

    \I__7746\ : Span4Mux_h
    port map (
            O => \N__32423\,
            I => \N__32363\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__32420\,
            I => \N__32354\
        );

    \I__7744\ : Span4Mux_v
    port map (
            O => \N__32417\,
            I => \N__32354\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__32414\,
            I => \N__32354\
        );

    \I__7742\ : Span4Mux_h
    port map (
            O => \N__32411\,
            I => \N__32354\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__32400\,
            I => \N__32351\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32348\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__32394\,
            I => \N__32343\
        );

    \I__7738\ : Span4Mux_v
    port map (
            O => \N__32391\,
            I => \N__32343\
        );

    \I__7737\ : Span4Mux_v
    port map (
            O => \N__32380\,
            I => \N__32340\
        );

    \I__7736\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32333\
        );

    \I__7735\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32333\
        );

    \I__7734\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32333\
        );

    \I__7733\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32330\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__32363\,
            I => \N__32327\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__32354\,
            I => \N__32324\
        );

    \I__7730\ : Span4Mux_v
    port map (
            O => \N__32351\,
            I => \N__32321\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__32348\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7728\ : Odrv4
    port map (
            O => \N__32343\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7727\ : Odrv4
    port map (
            O => \N__32340\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__32333\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__32330\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__32327\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__32324\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__32321\,
            I => \c0.FRAME_MATCHER_wait_for_transmission\
        );

    \I__7721\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32300\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__32303\,
            I => \N__32297\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__32300\,
            I => \N__32279\
        );

    \I__7718\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32276\
        );

    \I__7717\ : InMux
    port map (
            O => \N__32296\,
            I => \N__32273\
        );

    \I__7716\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32268\
        );

    \I__7715\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32268\
        );

    \I__7714\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32265\
        );

    \I__7713\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32258\
        );

    \I__7712\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32258\
        );

    \I__7711\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32258\
        );

    \I__7710\ : InMux
    port map (
            O => \N__32289\,
            I => \N__32251\
        );

    \I__7709\ : InMux
    port map (
            O => \N__32288\,
            I => \N__32251\
        );

    \I__7708\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32251\
        );

    \I__7707\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32246\
        );

    \I__7706\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32246\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__32284\,
            I => \N__32223\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__32283\,
            I => \N__32213\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__32282\,
            I => \N__32208\
        );

    \I__7702\ : Span4Mux_h
    port map (
            O => \N__32279\,
            I => \N__32184\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32184\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__32273\,
            I => \N__32184\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__32268\,
            I => \N__32184\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32184\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__32258\,
            I => \N__32184\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__32251\,
            I => \N__32184\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__32246\,
            I => \N__32184\
        );

    \I__7694\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32179\
        );

    \I__7693\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32179\
        );

    \I__7692\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32174\
        );

    \I__7691\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32174\
        );

    \I__7690\ : CascadeMux
    port map (
            O => \N__32241\,
            I => \N__32166\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32157\
        );

    \I__7688\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32148\
        );

    \I__7687\ : InMux
    port map (
            O => \N__32238\,
            I => \N__32148\
        );

    \I__7686\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32148\
        );

    \I__7685\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32148\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32145\
        );

    \I__7683\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32139\
        );

    \I__7682\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32136\
        );

    \I__7681\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32117\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32117\
        );

    \I__7679\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32112\
        );

    \I__7678\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32112\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32106\
        );

    \I__7676\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32106\
        );

    \I__7675\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32101\
        );

    \I__7674\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32101\
        );

    \I__7673\ : CascadeMux
    port map (
            O => \N__32222\,
            I => \N__32096\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__32221\,
            I => \N__32093\
        );

    \I__7671\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32077\
        );

    \I__7670\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32077\
        );

    \I__7669\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32077\
        );

    \I__7668\ : CascadeMux
    port map (
            O => \N__32217\,
            I => \N__32073\
        );

    \I__7667\ : CascadeMux
    port map (
            O => \N__32216\,
            I => \N__32060\
        );

    \I__7666\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32049\
        );

    \I__7665\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32044\
        );

    \I__7664\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32044\
        );

    \I__7663\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32039\
        );

    \I__7662\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32039\
        );

    \I__7661\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32030\
        );

    \I__7660\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32030\
        );

    \I__7659\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32030\
        );

    \I__7658\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32030\
        );

    \I__7657\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32025\
        );

    \I__7656\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32025\
        );

    \I__7655\ : Span4Mux_v
    port map (
            O => \N__32184\,
            I => \N__32021\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__32179\,
            I => \N__32016\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__32174\,
            I => \N__32016\
        );

    \I__7652\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32011\
        );

    \I__7651\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32011\
        );

    \I__7650\ : CascadeMux
    port map (
            O => \N__32171\,
            I => \N__32008\
        );

    \I__7649\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \N__32001\
        );

    \I__7648\ : InMux
    port map (
            O => \N__32169\,
            I => \N__31991\
        );

    \I__7647\ : InMux
    port map (
            O => \N__32166\,
            I => \N__31986\
        );

    \I__7646\ : InMux
    port map (
            O => \N__32165\,
            I => \N__31986\
        );

    \I__7645\ : InMux
    port map (
            O => \N__32164\,
            I => \N__31975\
        );

    \I__7644\ : InMux
    port map (
            O => \N__32163\,
            I => \N__31975\
        );

    \I__7643\ : InMux
    port map (
            O => \N__32162\,
            I => \N__31975\
        );

    \I__7642\ : InMux
    port map (
            O => \N__32161\,
            I => \N__31975\
        );

    \I__7641\ : InMux
    port map (
            O => \N__32160\,
            I => \N__31975\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__31970\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__31970\
        );

    \I__7638\ : InMux
    port map (
            O => \N__32145\,
            I => \N__31967\
        );

    \I__7637\ : InMux
    port map (
            O => \N__32144\,
            I => \N__31964\
        );

    \I__7636\ : InMux
    port map (
            O => \N__32143\,
            I => \N__31961\
        );

    \I__7635\ : InMux
    port map (
            O => \N__32142\,
            I => \N__31958\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__32139\,
            I => \N__31953\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__31953\
        );

    \I__7632\ : InMux
    port map (
            O => \N__32135\,
            I => \N__31948\
        );

    \I__7631\ : InMux
    port map (
            O => \N__32134\,
            I => \N__31948\
        );

    \I__7630\ : InMux
    port map (
            O => \N__32133\,
            I => \N__31945\
        );

    \I__7629\ : CascadeMux
    port map (
            O => \N__32132\,
            I => \N__31933\
        );

    \I__7628\ : InMux
    port map (
            O => \N__32131\,
            I => \N__31927\
        );

    \I__7627\ : InMux
    port map (
            O => \N__32130\,
            I => \N__31924\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32129\,
            I => \N__31919\
        );

    \I__7625\ : InMux
    port map (
            O => \N__32128\,
            I => \N__31919\
        );

    \I__7624\ : InMux
    port map (
            O => \N__32127\,
            I => \N__31916\
        );

    \I__7623\ : InMux
    port map (
            O => \N__32126\,
            I => \N__31912\
        );

    \I__7622\ : InMux
    port map (
            O => \N__32125\,
            I => \N__31909\
        );

    \I__7621\ : InMux
    port map (
            O => \N__32124\,
            I => \N__31906\
        );

    \I__7620\ : InMux
    port map (
            O => \N__32123\,
            I => \N__31901\
        );

    \I__7619\ : InMux
    port map (
            O => \N__32122\,
            I => \N__31901\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__31896\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__31896\
        );

    \I__7616\ : InMux
    port map (
            O => \N__32111\,
            I => \N__31893\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__31888\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__31888\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__32100\,
            I => \N__31884\
        );

    \I__7612\ : InMux
    port map (
            O => \N__32099\,
            I => \N__31877\
        );

    \I__7611\ : InMux
    port map (
            O => \N__32096\,
            I => \N__31877\
        );

    \I__7610\ : InMux
    port map (
            O => \N__32093\,
            I => \N__31868\
        );

    \I__7609\ : InMux
    port map (
            O => \N__32092\,
            I => \N__31868\
        );

    \I__7608\ : InMux
    port map (
            O => \N__32091\,
            I => \N__31868\
        );

    \I__7607\ : InMux
    port map (
            O => \N__32090\,
            I => \N__31868\
        );

    \I__7606\ : InMux
    port map (
            O => \N__32089\,
            I => \N__31863\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32088\,
            I => \N__31863\
        );

    \I__7604\ : InMux
    port map (
            O => \N__32087\,
            I => \N__31854\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32086\,
            I => \N__31854\
        );

    \I__7602\ : InMux
    port map (
            O => \N__32085\,
            I => \N__31854\
        );

    \I__7601\ : InMux
    port map (
            O => \N__32084\,
            I => \N__31854\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__31851\
        );

    \I__7599\ : InMux
    port map (
            O => \N__32076\,
            I => \N__31840\
        );

    \I__7598\ : InMux
    port map (
            O => \N__32073\,
            I => \N__31840\
        );

    \I__7597\ : InMux
    port map (
            O => \N__32072\,
            I => \N__31835\
        );

    \I__7596\ : InMux
    port map (
            O => \N__32071\,
            I => \N__31835\
        );

    \I__7595\ : InMux
    port map (
            O => \N__32070\,
            I => \N__31830\
        );

    \I__7594\ : InMux
    port map (
            O => \N__32069\,
            I => \N__31830\
        );

    \I__7593\ : InMux
    port map (
            O => \N__32068\,
            I => \N__31821\
        );

    \I__7592\ : InMux
    port map (
            O => \N__32067\,
            I => \N__31821\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32066\,
            I => \N__31821\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32065\,
            I => \N__31821\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32064\,
            I => \N__31818\
        );

    \I__7588\ : InMux
    port map (
            O => \N__32063\,
            I => \N__31815\
        );

    \I__7587\ : InMux
    port map (
            O => \N__32060\,
            I => \N__31804\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32059\,
            I => \N__31804\
        );

    \I__7585\ : InMux
    port map (
            O => \N__32058\,
            I => \N__31804\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32057\,
            I => \N__31804\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32056\,
            I => \N__31804\
        );

    \I__7582\ : InMux
    port map (
            O => \N__32055\,
            I => \N__31795\
        );

    \I__7581\ : InMux
    port map (
            O => \N__32054\,
            I => \N__31795\
        );

    \I__7580\ : InMux
    port map (
            O => \N__32053\,
            I => \N__31795\
        );

    \I__7579\ : InMux
    port map (
            O => \N__32052\,
            I => \N__31795\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__32049\,
            I => \N__31788\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__31788\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__32039\,
            I => \N__31788\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__31785\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__31782\
        );

    \I__7573\ : InMux
    port map (
            O => \N__32024\,
            I => \N__31779\
        );

    \I__7572\ : Span4Mux_h
    port map (
            O => \N__32021\,
            I => \N__31772\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__32016\,
            I => \N__31772\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__31772\
        );

    \I__7569\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31769\
        );

    \I__7568\ : InMux
    port map (
            O => \N__32007\,
            I => \N__31762\
        );

    \I__7567\ : InMux
    port map (
            O => \N__32006\,
            I => \N__31762\
        );

    \I__7566\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31762\
        );

    \I__7565\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31751\
        );

    \I__7564\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31751\
        );

    \I__7563\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31751\
        );

    \I__7562\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31751\
        );

    \I__7561\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31751\
        );

    \I__7560\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31746\
        );

    \I__7559\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31746\
        );

    \I__7558\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31741\
        );

    \I__7557\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31741\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__31991\,
            I => \N__31734\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__31986\,
            I => \N__31734\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__31975\,
            I => \N__31734\
        );

    \I__7553\ : Span4Mux_h
    port map (
            O => \N__31970\,
            I => \N__31721\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31721\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__31964\,
            I => \N__31721\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31721\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__31958\,
            I => \N__31721\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__31953\,
            I => \N__31721\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__31948\,
            I => \N__31716\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__31945\,
            I => \N__31716\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__31944\,
            I => \N__31701\
        );

    \I__7544\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31694\
        );

    \I__7543\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31694\
        );

    \I__7542\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31689\
        );

    \I__7541\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31689\
        );

    \I__7540\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31680\
        );

    \I__7539\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31680\
        );

    \I__7538\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31680\
        );

    \I__7537\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31680\
        );

    \I__7536\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31671\
        );

    \I__7535\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31671\
        );

    \I__7534\ : InMux
    port map (
            O => \N__31931\,
            I => \N__31671\
        );

    \I__7533\ : InMux
    port map (
            O => \N__31930\,
            I => \N__31671\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31662\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__31924\,
            I => \N__31662\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__31919\,
            I => \N__31662\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__31916\,
            I => \N__31662\
        );

    \I__7528\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31659\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__31912\,
            I => \N__31656\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31651\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__31906\,
            I => \N__31651\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__31901\,
            I => \N__31646\
        );

    \I__7523\ : Span4Mux_v
    port map (
            O => \N__31896\,
            I => \N__31646\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31641\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__31888\,
            I => \N__31641\
        );

    \I__7520\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31632\
        );

    \I__7519\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31632\
        );

    \I__7518\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31632\
        );

    \I__7517\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31632\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__31877\,
            I => \N__31621\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__31868\,
            I => \N__31621\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31621\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__31854\,
            I => \N__31621\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__31851\,
            I => \N__31621\
        );

    \I__7511\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31618\
        );

    \I__7510\ : InMux
    port map (
            O => \N__31849\,
            I => \N__31615\
        );

    \I__7509\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31606\
        );

    \I__7508\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31606\
        );

    \I__7507\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31606\
        );

    \I__7506\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31606\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31595\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31595\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31595\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__31821\,
            I => \N__31595\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31818\,
            I => \N__31595\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31592\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31581\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__31795\,
            I => \N__31581\
        );

    \I__7497\ : Span4Mux_h
    port map (
            O => \N__31788\,
            I => \N__31581\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__31785\,
            I => \N__31581\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__31782\,
            I => \N__31581\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31578\
        );

    \I__7493\ : Span4Mux_v
    port map (
            O => \N__31772\,
            I => \N__31575\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31562\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31562\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__31751\,
            I => \N__31562\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__31746\,
            I => \N__31562\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__31741\,
            I => \N__31562\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__31734\,
            I => \N__31562\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__31721\,
            I => \N__31559\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__31716\,
            I => \N__31556\
        );

    \I__7484\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31551\
        );

    \I__7483\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31551\
        );

    \I__7482\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31548\
        );

    \I__7481\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31541\
        );

    \I__7480\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31541\
        );

    \I__7479\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31541\
        );

    \I__7478\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31530\
        );

    \I__7477\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31530\
        );

    \I__7476\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31530\
        );

    \I__7475\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31530\
        );

    \I__7474\ : InMux
    port map (
            O => \N__31705\,
            I => \N__31530\
        );

    \I__7473\ : InMux
    port map (
            O => \N__31704\,
            I => \N__31521\
        );

    \I__7472\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31521\
        );

    \I__7471\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31521\
        );

    \I__7470\ : InMux
    port map (
            O => \N__31699\,
            I => \N__31521\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__31694\,
            I => \N__31512\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__31689\,
            I => \N__31512\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__31680\,
            I => \N__31512\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__31671\,
            I => \N__31512\
        );

    \I__7465\ : Span4Mux_v
    port map (
            O => \N__31662\,
            I => \N__31509\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__31659\,
            I => \N__31498\
        );

    \I__7463\ : Span4Mux_v
    port map (
            O => \N__31656\,
            I => \N__31498\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__31651\,
            I => \N__31498\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__31646\,
            I => \N__31498\
        );

    \I__7460\ : Span4Mux_h
    port map (
            O => \N__31641\,
            I => \N__31498\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__31632\,
            I => \N__31493\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__31621\,
            I => \N__31493\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31482\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31482\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__31606\,
            I => \N__31482\
        );

    \I__7454\ : Span12Mux_v
    port map (
            O => \N__31595\,
            I => \N__31482\
        );

    \I__7453\ : Span12Mux_v
    port map (
            O => \N__31592\,
            I => \N__31482\
        );

    \I__7452\ : Span4Mux_v
    port map (
            O => \N__31581\,
            I => \N__31479\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__31578\,
            I => \N__31468\
        );

    \I__7450\ : Span4Mux_h
    port map (
            O => \N__31575\,
            I => \N__31468\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__31562\,
            I => \N__31468\
        );

    \I__7448\ : Span4Mux_h
    port map (
            O => \N__31559\,
            I => \N__31468\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__31556\,
            I => \N__31468\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__31551\,
            I => \c0.n1729\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__31548\,
            I => \c0.n1729\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__31541\,
            I => \c0.n1729\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__31530\,
            I => \c0.n1729\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__31521\,
            I => \c0.n1729\
        );

    \I__7441\ : Odrv12
    port map (
            O => \N__31512\,
            I => \c0.n1729\
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__31509\,
            I => \c0.n1729\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__31498\,
            I => \c0.n1729\
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__31493\,
            I => \c0.n1729\
        );

    \I__7437\ : Odrv12
    port map (
            O => \N__31482\,
            I => \c0.n1729\
        );

    \I__7436\ : Odrv4
    port map (
            O => \N__31479\,
            I => \c0.n1729\
        );

    \I__7435\ : Odrv4
    port map (
            O => \N__31468\,
            I => \c0.n1729\
        );

    \I__7434\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31440\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31437\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__31437\,
            I => \N__31433\
        );

    \I__7431\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31429\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__31433\,
            I => \N__31426\
        );

    \I__7429\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31423\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__31429\,
            I => data_in_4_7
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__31426\,
            I => data_in_4_7
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__31423\,
            I => data_in_4_7
        );

    \I__7425\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31408\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__31412\,
            I => \N__31404\
        );

    \I__7422\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31401\
        );

    \I__7421\ : Span4Mux_v
    port map (
            O => \N__31408\,
            I => \N__31397\
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__31407\,
            I => \N__31394\
        );

    \I__7419\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31391\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31388\
        );

    \I__7417\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31385\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__31397\,
            I => \N__31382\
        );

    \I__7415\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31379\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__31391\,
            I => \c0.data_in_field_39\
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__31388\,
            I => \c0.data_in_field_39\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__31385\,
            I => \c0.data_in_field_39\
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__31382\,
            I => \c0.data_in_field_39\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__31379\,
            I => \c0.data_in_field_39\
        );

    \I__7409\ : InMux
    port map (
            O => \N__31368\,
            I => \N__31364\
        );

    \I__7408\ : InMux
    port map (
            O => \N__31367\,
            I => \N__31361\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31358\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__31361\,
            I => \N__31354\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__31358\,
            I => \N__31351\
        );

    \I__7404\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31348\
        );

    \I__7403\ : Odrv12
    port map (
            O => \N__31354\,
            I => data_in_10_7
        );

    \I__7402\ : Odrv4
    port map (
            O => \N__31351\,
            I => data_in_10_7
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__31348\,
            I => data_in_10_7
        );

    \I__7400\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__31338\,
            I => \N__31334\
        );

    \I__7398\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31331\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__31334\,
            I => \N__31326\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31326\
        );

    \I__7395\ : Sp12to4
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__7394\ : Span12Mux_s11_v
    port map (
            O => \N__31323\,
            I => \N__31319\
        );

    \I__7393\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31316\
        );

    \I__7392\ : Odrv12
    port map (
            O => \N__31319\,
            I => data_in_9_7
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__31316\,
            I => data_in_9_7
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__31311\,
            I => \N__31307\
        );

    \I__7389\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31304\
        );

    \I__7388\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31301\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31298\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31294\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__31298\,
            I => \N__31291\
        );

    \I__7384\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31288\
        );

    \I__7383\ : Odrv12
    port map (
            O => \N__31294\,
            I => data_in_14_5
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__31291\,
            I => data_in_14_5
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__31288\,
            I => data_in_14_5
        );

    \I__7380\ : CascadeMux
    port map (
            O => \N__31281\,
            I => \N__31278\
        );

    \I__7379\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31271\
        );

    \I__7378\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31271\
        );

    \I__7377\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31268\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31265\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__31268\,
            I => data_in_12_2
        );

    \I__7374\ : Odrv4
    port map (
            O => \N__31265\,
            I => data_in_12_2
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__31260\,
            I => \N__31257\
        );

    \I__7372\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31250\
        );

    \I__7370\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31247\
        );

    \I__7369\ : Span4Mux_v
    port map (
            O => \N__31250\,
            I => \N__31243\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__31247\,
            I => \N__31240\
        );

    \I__7367\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31237\
        );

    \I__7366\ : Odrv4
    port map (
            O => \N__31243\,
            I => data_in_11_2
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__31240\,
            I => data_in_11_2
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__31237\,
            I => data_in_11_2
        );

    \I__7363\ : CascadeMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__7362\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__31224\,
            I => \N__31220\
        );

    \I__7360\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31217\
        );

    \I__7359\ : Span4Mux_h
    port map (
            O => \N__31220\,
            I => \N__31214\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31211\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__31214\,
            I => \N__31205\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__31211\,
            I => \N__31205\
        );

    \I__7355\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31202\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__31205\,
            I => data_in_4_4
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__31202\,
            I => data_in_4_4
        );

    \I__7352\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31190\
        );

    \I__7350\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31187\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__31190\,
            I => \N__31184\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__31187\,
            I => \N__31178\
        );

    \I__7347\ : Sp12to4
    port map (
            O => \N__31184\,
            I => \N__31178\
        );

    \I__7346\ : InMux
    port map (
            O => \N__31183\,
            I => \N__31175\
        );

    \I__7345\ : Odrv12
    port map (
            O => \N__31178\,
            I => data_in_9_6
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__31175\,
            I => data_in_9_6
        );

    \I__7343\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31166\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__31169\,
            I => \N__31163\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__31166\,
            I => \N__31160\
        );

    \I__7340\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31157\
        );

    \I__7339\ : Span4Mux_v
    port map (
            O => \N__31160\,
            I => \N__31154\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31150\
        );

    \I__7337\ : Span4Mux_h
    port map (
            O => \N__31154\,
            I => \N__31147\
        );

    \I__7336\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31144\
        );

    \I__7335\ : Odrv12
    port map (
            O => \N__31150\,
            I => data_in_8_6
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__31147\,
            I => data_in_8_6
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__31144\,
            I => data_in_8_6
        );

    \I__7332\ : CascadeMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__7331\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31127\
        );

    \I__7329\ : CascadeMux
    port map (
            O => \N__31130\,
            I => \N__31122\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__31127\,
            I => \N__31119\
        );

    \I__7327\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31114\
        );

    \I__7326\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31114\
        );

    \I__7325\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31111\
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__31119\,
            I => data_in_3_4
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__31114\,
            I => data_in_3_4
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__31111\,
            I => data_in_3_4
        );

    \I__7321\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31099\
        );

    \I__7320\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31096\
        );

    \I__7319\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31093\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__31099\,
            I => \N__31090\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__31096\,
            I => \N__31084\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31084\
        );

    \I__7315\ : Span4Mux_v
    port map (
            O => \N__31090\,
            I => \N__31081\
        );

    \I__7314\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31078\
        );

    \I__7313\ : Span4Mux_h
    port map (
            O => \N__31084\,
            I => \N__31075\
        );

    \I__7312\ : Odrv4
    port map (
            O => \N__31081\,
            I => data_in_2_4
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__31078\,
            I => data_in_2_4
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__31075\,
            I => data_in_2_4
        );

    \I__7309\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__31065\,
            I => \c0.n50_adj_1875\
        );

    \I__7307\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__31059\,
            I => \N__31055\
        );

    \I__7305\ : InMux
    port map (
            O => \N__31058\,
            I => \N__31052\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__31055\,
            I => \N__31049\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__31052\,
            I => \N__31046\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__7301\ : Span4Mux_h
    port map (
            O => \N__31046\,
            I => \N__31040\
        );

    \I__7300\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31037\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__31040\,
            I => data_in_8_0
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__31037\,
            I => data_in_8_0
        );

    \I__7297\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31028\
        );

    \I__7296\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31024\
        );

    \I__7295\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31019\
        );

    \I__7294\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31019\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__31024\,
            I => data_in_7_0
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__31019\,
            I => data_in_7_0
        );

    \I__7291\ : InMux
    port map (
            O => \N__31014\,
            I => \N__31010\
        );

    \I__7290\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31007\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__31004\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__31007\,
            I => \N__31001\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__31004\,
            I => \N__30997\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__31001\,
            I => \N__30994\
        );

    \I__7285\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30990\
        );

    \I__7284\ : Span4Mux_h
    port map (
            O => \N__30997\,
            I => \N__30985\
        );

    \I__7283\ : Span4Mux_h
    port map (
            O => \N__30994\,
            I => \N__30985\
        );

    \I__7282\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30982\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__30990\,
            I => \c0.data_in_field_74\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__30985\,
            I => \c0.data_in_field_74\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__30982\,
            I => \c0.data_in_field_74\
        );

    \I__7278\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30971\
        );

    \I__7277\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30968\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__30971\,
            I => \N__30963\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30960\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__30967\,
            I => \N__30957\
        );

    \I__7273\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30954\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__30963\,
            I => \N__30951\
        );

    \I__7271\ : Span12Mux_h
    port map (
            O => \N__30960\,
            I => \N__30948\
        );

    \I__7270\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30945\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__30954\,
            I => \c0.data_in_field_1\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__30951\,
            I => \c0.data_in_field_1\
        );

    \I__7267\ : Odrv12
    port map (
            O => \N__30948\,
            I => \c0.data_in_field_1\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__30945\,
            I => \c0.data_in_field_1\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__30936\,
            I => \N__30930\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__30935\,
            I => \N__30927\
        );

    \I__7263\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30923\
        );

    \I__7262\ : InMux
    port map (
            O => \N__30933\,
            I => \N__30920\
        );

    \I__7261\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30917\
        );

    \I__7260\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30912\
        );

    \I__7259\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30912\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__30923\,
            I => \c0.data_in_field_16\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__30920\,
            I => \c0.data_in_field_16\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__30917\,
            I => \c0.data_in_field_16\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30912\,
            I => \c0.data_in_field_16\
        );

    \I__7254\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__30900\,
            I => \c0.n25_adj_1931\
        );

    \I__7252\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30893\
        );

    \I__7251\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30889\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__30893\,
            I => \N__30886\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30883\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30878\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__30886\,
            I => \N__30875\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__30883\,
            I => \N__30872\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__30882\,
            I => \N__30869\
        );

    \I__7244\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30866\
        );

    \I__7243\ : Span4Mux_v
    port map (
            O => \N__30878\,
            I => \N__30863\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__30875\,
            I => \N__30858\
        );

    \I__7241\ : Span4Mux_v
    port map (
            O => \N__30872\,
            I => \N__30858\
        );

    \I__7240\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30855\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__30866\,
            I => \c0.data_in_field_137\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__30863\,
            I => \c0.data_in_field_137\
        );

    \I__7237\ : Odrv4
    port map (
            O => \N__30858\,
            I => \c0.data_in_field_137\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30855\,
            I => \c0.data_in_field_137\
        );

    \I__7235\ : CascadeMux
    port map (
            O => \N__30846\,
            I => \N__30842\
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__7233\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30836\
        );

    \I__7232\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30833\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__30836\,
            I => \N__30830\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__30833\,
            I => \N__30825\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__30830\,
            I => \N__30822\
        );

    \I__7228\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30818\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__30828\,
            I => \N__30815\
        );

    \I__7226\ : Span4Mux_v
    port map (
            O => \N__30825\,
            I => \N__30812\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__30822\,
            I => \N__30809\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__30821\,
            I => \N__30806\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30803\
        );

    \I__7222\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30800\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__30812\,
            I => \N__30795\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__30809\,
            I => \N__30795\
        );

    \I__7219\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30792\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__30803\,
            I => \N__30789\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__30800\,
            I => \c0.data_in_field_25\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__30795\,
            I => \c0.data_in_field_25\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__30792\,
            I => \c0.data_in_field_25\
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__30789\,
            I => \c0.data_in_field_25\
        );

    \I__7213\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30776\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30772\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30769\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__30775\,
            I => \N__30765\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__30772\,
            I => \N__30762\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__30769\,
            I => \N__30759\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30756\
        );

    \I__7206\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30753\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__30762\,
            I => \N__30750\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__30759\,
            I => \N__30747\
        );

    \I__7203\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30744\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__30753\,
            I => \c0.data_in_field_71\
        );

    \I__7201\ : Odrv4
    port map (
            O => \N__30750\,
            I => \c0.data_in_field_71\
        );

    \I__7200\ : Odrv4
    port map (
            O => \N__30747\,
            I => \c0.data_in_field_71\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__30744\,
            I => \c0.data_in_field_71\
        );

    \I__7198\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30731\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__30734\,
            I => \N__30728\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__30731\,
            I => \N__30725\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30722\
        );

    \I__7194\ : Span4Mux_h
    port map (
            O => \N__30725\,
            I => \N__30719\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30716\
        );

    \I__7192\ : Span4Mux_h
    port map (
            O => \N__30719\,
            I => \N__30713\
        );

    \I__7191\ : Span4Mux_h
    port map (
            O => \N__30716\,
            I => \N__30710\
        );

    \I__7190\ : Odrv4
    port map (
            O => \N__30713\,
            I => \c0.n5542\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__30710\,
            I => \c0.n5542\
        );

    \I__7188\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__30696\,
            I => \N__30691\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30688\
        );

    \I__7183\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30685\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__30691\,
            I => data_in_17_0
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__30688\,
            I => data_in_17_0
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__30685\,
            I => data_in_17_0
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30668\
        );

    \I__7176\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__7175\ : Span4Mux_h
    port map (
            O => \N__30668\,
            I => \N__30662\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30659\
        );

    \I__7173\ : Span4Mux_h
    port map (
            O => \N__30662\,
            I => \N__30655\
        );

    \I__7172\ : Span12Mux_v
    port map (
            O => \N__30659\,
            I => \N__30652\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__30655\,
            I => data_in_10_2
        );

    \I__7169\ : Odrv12
    port map (
            O => \N__30652\,
            I => data_in_10_2
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__30649\,
            I => data_in_10_2
        );

    \I__7167\ : CascadeMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__7166\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__7164\ : Span4Mux_h
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__30630\,
            I => \N__30625\
        );

    \I__7162\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30620\
        );

    \I__7161\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30620\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__30625\,
            I => data_in_4_6
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30620\,
            I => data_in_4_6
        );

    \I__7158\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30611\
        );

    \I__7157\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30608\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__30611\,
            I => \N__30600\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30600\
        );

    \I__7154\ : InMux
    port map (
            O => \N__30607\,
            I => \N__30597\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__30606\,
            I => \N__30594\
        );

    \I__7152\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30590\
        );

    \I__7151\ : Span12Mux_v
    port map (
            O => \N__30600\,
            I => \N__30585\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__30597\,
            I => \N__30585\
        );

    \I__7149\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30580\
        );

    \I__7148\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30580\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__30590\,
            I => \c0.data_in_field_38\
        );

    \I__7146\ : Odrv12
    port map (
            O => \N__30585\,
            I => \c0.data_in_field_38\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__30580\,
            I => \c0.data_in_field_38\
        );

    \I__7144\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__30570\,
            I => \N__30565\
        );

    \I__7142\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30562\
        );

    \I__7141\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30557\
        );

    \I__7140\ : Span12Mux_h
    port map (
            O => \N__30565\,
            I => \N__30554\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__30562\,
            I => \N__30551\
        );

    \I__7138\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30548\
        );

    \I__7137\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30545\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__30557\,
            I => \c0.data_in_field_136\
        );

    \I__7135\ : Odrv12
    port map (
            O => \N__30554\,
            I => \c0.data_in_field_136\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__30551\,
            I => \c0.data_in_field_136\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__30548\,
            I => \c0.data_in_field_136\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__30545\,
            I => \c0.data_in_field_136\
        );

    \I__7131\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__30531\,
            I => \N__30526\
        );

    \I__7129\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30523\
        );

    \I__7128\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30519\
        );

    \I__7127\ : Span4Mux_v
    port map (
            O => \N__30526\,
            I => \N__30515\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30512\
        );

    \I__7125\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30509\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30506\
        );

    \I__7123\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30503\
        );

    \I__7122\ : Sp12to4
    port map (
            O => \N__30515\,
            I => \N__30498\
        );

    \I__7121\ : Sp12to4
    port map (
            O => \N__30512\,
            I => \N__30498\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__30509\,
            I => \c0.data_in_field_31\
        );

    \I__7119\ : Odrv12
    port map (
            O => \N__30506\,
            I => \c0.data_in_field_31\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__30503\,
            I => \c0.data_in_field_31\
        );

    \I__7117\ : Odrv12
    port map (
            O => \N__30498\,
            I => \c0.data_in_field_31\
        );

    \I__7116\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__30486\,
            I => \c0.n2113\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__30483\,
            I => \N__30479\
        );

    \I__7113\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30476\
        );

    \I__7112\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30473\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30470\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__30473\,
            I => \N__30466\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__30470\,
            I => \N__30463\
        );

    \I__7108\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30460\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__30466\,
            I => data_in_11_0
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__30463\,
            I => data_in_11_0
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__30460\,
            I => data_in_11_0
        );

    \I__7104\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30449\
        );

    \I__7103\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30446\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30443\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__30446\,
            I => \N__30440\
        );

    \I__7100\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30434\
        );

    \I__7099\ : Span4Mux_v
    port map (
            O => \N__30440\,
            I => \N__30434\
        );

    \I__7098\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30431\
        );

    \I__7097\ : Span4Mux_h
    port map (
            O => \N__30434\,
            I => \N__30428\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__30431\,
            I => data_in_10_0
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__30428\,
            I => data_in_10_0
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__7093\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30416\
        );

    \I__7092\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__30416\,
            I => \N__30410\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__30413\,
            I => \N__30407\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__30410\,
            I => \N__30403\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__30407\,
            I => \N__30400\
        );

    \I__7087\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30397\
        );

    \I__7086\ : Odrv4
    port map (
            O => \N__30403\,
            I => data_in_10_4
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__30400\,
            I => data_in_10_4
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__30397\,
            I => data_in_10_4
        );

    \I__7083\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30387\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30383\
        );

    \I__7081\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30380\
        );

    \I__7080\ : Span4Mux_h
    port map (
            O => \N__30383\,
            I => \N__30377\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30374\
        );

    \I__7078\ : Span4Mux_h
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__30374\,
            I => \N__30368\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__30371\,
            I => \N__30364\
        );

    \I__7075\ : Span4Mux_h
    port map (
            O => \N__30368\,
            I => \N__30361\
        );

    \I__7074\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30358\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__30364\,
            I => data_in_9_4
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__30361\,
            I => data_in_9_4
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__30358\,
            I => data_in_9_4
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__7069\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__30342\,
            I => \N__30337\
        );

    \I__7066\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30334\
        );

    \I__7065\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30331\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__30337\,
            I => data_in_16_4
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__30334\,
            I => data_in_16_4
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__30331\,
            I => data_in_16_4
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__7060\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__7058\ : Span4Mux_h
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__7057\ : Span4Mux_h
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__30309\,
            I => \N__30304\
        );

    \I__7055\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30301\
        );

    \I__7054\ : InMux
    port map (
            O => \N__30307\,
            I => \N__30298\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__30304\,
            I => data_in_15_4
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__30301\,
            I => data_in_15_4
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__30298\,
            I => data_in_15_4
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__30291\,
            I => \N__30287\
        );

    \I__7049\ : CascadeMux
    port map (
            O => \N__30290\,
            I => \N__30284\
        );

    \I__7048\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30281\
        );

    \I__7047\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30277\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__30281\,
            I => \N__30274\
        );

    \I__7045\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30271\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__30277\,
            I => data_in_13_4
        );

    \I__7043\ : Odrv4
    port map (
            O => \N__30274\,
            I => data_in_13_4
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__30271\,
            I => data_in_13_4
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__7040\ : InMux
    port map (
            O => \N__30261\,
            I => \N__30257\
        );

    \I__7039\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30254\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30251\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__30254\,
            I => \N__30247\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__30251\,
            I => \N__30244\
        );

    \I__7035\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30240\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__30247\,
            I => \N__30237\
        );

    \I__7033\ : Span4Mux_v
    port map (
            O => \N__30244\,
            I => \N__30234\
        );

    \I__7032\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30231\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30225\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__30237\,
            I => \N__30225\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__30234\,
            I => \N__30220\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__30231\,
            I => \N__30220\
        );

    \I__7027\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30217\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__30225\,
            I => \c0.data_in_field_108\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__30220\,
            I => \c0.data_in_field_108\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__30217\,
            I => \c0.data_in_field_108\
        );

    \I__7023\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30201\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__30209\,
            I => \N__30195\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__30208\,
            I => \N__30190\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__30207\,
            I => \N__30187\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__30206\,
            I => \N__30181\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__30205\,
            I => \N__30177\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__30204\,
            I => \N__30167\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__30201\,
            I => \N__30164\
        );

    \I__7015\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30161\
        );

    \I__7014\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30154\
        );

    \I__7013\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30154\
        );

    \I__7012\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30154\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__30194\,
            I => \N__30150\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__30193\,
            I => \N__30141\
        );

    \I__7009\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30136\
        );

    \I__7008\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30136\
        );

    \I__7007\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30133\
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__30185\,
            I => \N__30129\
        );

    \I__7005\ : CascadeMux
    port map (
            O => \N__30184\,
            I => \N__30122\
        );

    \I__7004\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30114\
        );

    \I__7003\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30114\
        );

    \I__7002\ : InMux
    port map (
            O => \N__30177\,
            I => \N__30114\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__30176\,
            I => \N__30106\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30102\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__30174\,
            I => \N__30097\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__30173\,
            I => \N__30094\
        );

    \I__6997\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30090\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__30171\,
            I => \N__30086\
        );

    \I__6995\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30081\
        );

    \I__6994\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30081\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__30164\,
            I => \N__30074\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__30161\,
            I => \N__30074\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30074\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__30153\,
            I => \N__30071\
        );

    \I__6989\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30066\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__30149\,
            I => \N__30062\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__30148\,
            I => \N__30056\
        );

    \I__6986\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30050\
        );

    \I__6985\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30047\
        );

    \I__6984\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30040\
        );

    \I__6983\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30040\
        );

    \I__6982\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30040\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__30136\,
            I => \N__30035\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30035\
        );

    \I__6979\ : InMux
    port map (
            O => \N__30132\,
            I => \N__30030\
        );

    \I__6978\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30030\
        );

    \I__6977\ : CascadeMux
    port map (
            O => \N__30128\,
            I => \N__30026\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__30127\,
            I => \N__30022\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__30126\,
            I => \N__30019\
        );

    \I__6974\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30009\
        );

    \I__6973\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30009\
        );

    \I__6972\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30009\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30006\
        );

    \I__6970\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30003\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__30112\,
            I => \N__30000\
        );

    \I__6968\ : InMux
    port map (
            O => \N__30111\,
            I => \N__29994\
        );

    \I__6967\ : InMux
    port map (
            O => \N__30110\,
            I => \N__29994\
        );

    \I__6966\ : InMux
    port map (
            O => \N__30109\,
            I => \N__29989\
        );

    \I__6965\ : InMux
    port map (
            O => \N__30106\,
            I => \N__29989\
        );

    \I__6964\ : InMux
    port map (
            O => \N__30105\,
            I => \N__29986\
        );

    \I__6963\ : InMux
    port map (
            O => \N__30102\,
            I => \N__29981\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30101\,
            I => \N__29981\
        );

    \I__6961\ : InMux
    port map (
            O => \N__30100\,
            I => \N__29978\
        );

    \I__6960\ : InMux
    port map (
            O => \N__30097\,
            I => \N__29975\
        );

    \I__6959\ : InMux
    port map (
            O => \N__30094\,
            I => \N__29972\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__30093\,
            I => \N__29967\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__30090\,
            I => \N__29964\
        );

    \I__6956\ : InMux
    port map (
            O => \N__30089\,
            I => \N__29959\
        );

    \I__6955\ : InMux
    port map (
            O => \N__30086\,
            I => \N__29959\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__30081\,
            I => \N__29956\
        );

    \I__6953\ : Span4Mux_h
    port map (
            O => \N__30074\,
            I => \N__29953\
        );

    \I__6952\ : InMux
    port map (
            O => \N__30071\,
            I => \N__29950\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__30070\,
            I => \N__29944\
        );

    \I__6950\ : CascadeMux
    port map (
            O => \N__30069\,
            I => \N__29940\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__29935\
        );

    \I__6948\ : InMux
    port map (
            O => \N__30065\,
            I => \N__29930\
        );

    \I__6947\ : InMux
    port map (
            O => \N__30062\,
            I => \N__29930\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__30061\,
            I => \N__29926\
        );

    \I__6945\ : CascadeMux
    port map (
            O => \N__30060\,
            I => \N__29921\
        );

    \I__6944\ : CascadeMux
    port map (
            O => \N__30059\,
            I => \N__29918\
        );

    \I__6943\ : InMux
    port map (
            O => \N__30056\,
            I => \N__29911\
        );

    \I__6942\ : InMux
    port map (
            O => \N__30055\,
            I => \N__29911\
        );

    \I__6941\ : InMux
    port map (
            O => \N__30054\,
            I => \N__29911\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30053\,
            I => \N__29908\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__29897\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__30047\,
            I => \N__29897\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__30040\,
            I => \N__29897\
        );

    \I__6936\ : Span4Mux_h
    port map (
            O => \N__30035\,
            I => \N__29897\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__29897\
        );

    \I__6934\ : InMux
    port map (
            O => \N__30029\,
            I => \N__29892\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30026\,
            I => \N__29892\
        );

    \I__6932\ : InMux
    port map (
            O => \N__30025\,
            I => \N__29883\
        );

    \I__6931\ : InMux
    port map (
            O => \N__30022\,
            I => \N__29883\
        );

    \I__6930\ : InMux
    port map (
            O => \N__30019\,
            I => \N__29883\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29883\
        );

    \I__6928\ : InMux
    port map (
            O => \N__30017\,
            I => \N__29878\
        );

    \I__6927\ : InMux
    port map (
            O => \N__30016\,
            I => \N__29878\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__30009\,
            I => \N__29875\
        );

    \I__6925\ : Span4Mux_v
    port map (
            O => \N__30006\,
            I => \N__29870\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__30003\,
            I => \N__29870\
        );

    \I__6923\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29867\
        );

    \I__6922\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29864\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29857\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29857\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__29986\,
            I => \N__29857\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29854\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__29978\,
            I => \N__29847\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__29975\,
            I => \N__29847\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__29972\,
            I => \N__29847\
        );

    \I__6914\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29842\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29842\
        );

    \I__6912\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29839\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__29964\,
            I => \N__29828\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29828\
        );

    \I__6909\ : Span4Mux_v
    port map (
            O => \N__29956\,
            I => \N__29828\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__29953\,
            I => \N__29828\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__29950\,
            I => \N__29828\
        );

    \I__6906\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29818\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29818\
        );

    \I__6904\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29813\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29813\
        );

    \I__6902\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29810\
        );

    \I__6901\ : InMux
    port map (
            O => \N__29940\,
            I => \N__29807\
        );

    \I__6900\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29804\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__29938\,
            I => \N__29799\
        );

    \I__6898\ : Span4Mux_h
    port map (
            O => \N__29935\,
            I => \N__29796\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__29930\,
            I => \N__29793\
        );

    \I__6896\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29787\
        );

    \I__6895\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29787\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__29925\,
            I => \N__29783\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__29924\,
            I => \N__29779\
        );

    \I__6892\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29776\
        );

    \I__6891\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29773\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29770\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29765\
        );

    \I__6888\ : Span4Mux_v
    port map (
            O => \N__29897\,
            I => \N__29765\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__29892\,
            I => \N__29752\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29752\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__29878\,
            I => \N__29752\
        );

    \I__6884\ : Span4Mux_v
    port map (
            O => \N__29875\,
            I => \N__29752\
        );

    \I__6883\ : Span4Mux_h
    port map (
            O => \N__29870\,
            I => \N__29752\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__29867\,
            I => \N__29752\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__29864\,
            I => \N__29745\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__29857\,
            I => \N__29745\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__29854\,
            I => \N__29745\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__29847\,
            I => \N__29742\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__29842\,
            I => \N__29735\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__29839\,
            I => \N__29735\
        );

    \I__6875\ : Span4Mux_v
    port map (
            O => \N__29828\,
            I => \N__29735\
        );

    \I__6874\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29732\
        );

    \I__6873\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29723\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29723\
        );

    \I__6871\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29723\
        );

    \I__6870\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29723\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__29818\,
            I => \N__29718\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__29813\,
            I => \N__29718\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29713\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__29807\,
            I => \N__29713\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__29804\,
            I => \N__29710\
        );

    \I__6864\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29703\
        );

    \I__6863\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29703\
        );

    \I__6862\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29703\
        );

    \I__6861\ : Span4Mux_h
    port map (
            O => \N__29796\,
            I => \N__29698\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__29793\,
            I => \N__29698\
        );

    \I__6859\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29695\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__29787\,
            I => \N__29692\
        );

    \I__6857\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29689\
        );

    \I__6856\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29686\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29683\
        );

    \I__6854\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29680\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__29776\,
            I => \N__29675\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__29773\,
            I => \N__29675\
        );

    \I__6851\ : Span4Mux_s2_h
    port map (
            O => \N__29770\,
            I => \N__29668\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__29765\,
            I => \N__29668\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__29752\,
            I => \N__29668\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__29745\,
            I => \N__29661\
        );

    \I__6847\ : Span4Mux_h
    port map (
            O => \N__29742\,
            I => \N__29661\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__29735\,
            I => \N__29661\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__29732\,
            I => \N__29646\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29646\
        );

    \I__6843\ : Span4Mux_s2_h
    port map (
            O => \N__29718\,
            I => \N__29646\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__29713\,
            I => \N__29646\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__29710\,
            I => \N__29646\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29646\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29646\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__29695\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__29692\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__29689\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__29686\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__29683\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__29680\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6832\ : Odrv12
    port map (
            O => \N__29675\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6831\ : Odrv4
    port map (
            O => \N__29668\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__29661\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__29646\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6828\ : CascadeMux
    port map (
            O => \N__29625\,
            I => \N__29622\
        );

    \I__6827\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29619\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29616\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__29613\,
            I => \N__29609\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29604\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__29609\,
            I => \N__29601\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29598\
        );

    \I__6820\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29595\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__29604\,
            I => \c0.data_in_field_47\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__29601\,
            I => \c0.data_in_field_47\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__29598\,
            I => \c0.data_in_field_47\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__29595\,
            I => \c0.data_in_field_47\
        );

    \I__6815\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__29583\,
            I => \c0.n5997\
        );

    \I__6813\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29577\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__6811\ : Span4Mux_v
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__6809\ : Span4Mux_h
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__29565\,
            I => \c0.n6000\
        );

    \I__6807\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29559\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__29559\,
            I => \N__29555\
        );

    \I__6805\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29552\
        );

    \I__6804\ : Span4Mux_v
    port map (
            O => \N__29555\,
            I => \N__29549\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__29552\,
            I => \N__29546\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__29549\,
            I => \N__29543\
        );

    \I__6801\ : Span4Mux_v
    port map (
            O => \N__29546\,
            I => \N__29539\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__29543\,
            I => \N__29536\
        );

    \I__6799\ : InMux
    port map (
            O => \N__29542\,
            I => \N__29532\
        );

    \I__6798\ : Span4Mux_h
    port map (
            O => \N__29539\,
            I => \N__29529\
        );

    \I__6797\ : Span4Mux_v
    port map (
            O => \N__29536\,
            I => \N__29526\
        );

    \I__6796\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29523\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__29532\,
            I => \c0.data_in_field_84\
        );

    \I__6794\ : Odrv4
    port map (
            O => \N__29529\,
            I => \c0.data_in_field_84\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__29526\,
            I => \c0.data_in_field_84\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__29523\,
            I => \c0.data_in_field_84\
        );

    \I__6791\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29510\
        );

    \I__6790\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29507\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__29510\,
            I => \N__29504\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__29507\,
            I => \N__29500\
        );

    \I__6787\ : Span4Mux_h
    port map (
            O => \N__29504\,
            I => \N__29497\
        );

    \I__6786\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29494\
        );

    \I__6785\ : Sp12to4
    port map (
            O => \N__29500\,
            I => \N__29491\
        );

    \I__6784\ : Span4Mux_h
    port map (
            O => \N__29497\,
            I => \N__29488\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__29494\,
            I => \N__29485\
        );

    \I__6782\ : Span12Mux_v
    port map (
            O => \N__29491\,
            I => \N__29480\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__29488\,
            I => \N__29477\
        );

    \I__6780\ : Span4Mux_h
    port map (
            O => \N__29485\,
            I => \N__29474\
        );

    \I__6779\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29469\
        );

    \I__6778\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29469\
        );

    \I__6777\ : Odrv12
    port map (
            O => \N__29480\,
            I => \c0.data_in_field_70\
        );

    \I__6776\ : Odrv4
    port map (
            O => \N__29477\,
            I => \c0.data_in_field_70\
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__29474\,
            I => \c0.data_in_field_70\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__29469\,
            I => \c0.data_in_field_70\
        );

    \I__6773\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29455\
        );

    \I__6772\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29450\
        );

    \I__6771\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29450\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__29455\,
            I => \c0.data_in_field_56\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__29450\,
            I => \c0.data_in_field_56\
        );

    \I__6768\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__29436\,
            I => \c0.n5494\
        );

    \I__6764\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29426\
        );

    \I__6762\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29423\
        );

    \I__6761\ : Span4Mux_s3_h
    port map (
            O => \N__29426\,
            I => \N__29420\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29417\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__29420\,
            I => \c0.n5554\
        );

    \I__6758\ : Odrv12
    port map (
            O => \N__29417\,
            I => \c0.n5554\
        );

    \I__6757\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29405\
        );

    \I__6755\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29402\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__29405\,
            I => \N__29399\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__29402\,
            I => \N__29396\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29393\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__29396\,
            I => \N__29388\
        );

    \I__6750\ : Span4Mux_h
    port map (
            O => \N__29393\,
            I => \N__29388\
        );

    \I__6749\ : Odrv4
    port map (
            O => \N__29388\,
            I => \c0.n5524\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__29385\,
            I => \c0.n5494_cascade_\
        );

    \I__6747\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29379\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__29379\,
            I => \N__29375\
        );

    \I__6745\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29372\
        );

    \I__6744\ : Span4Mux_v
    port map (
            O => \N__29375\,
            I => \N__29369\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__29372\,
            I => \N__29366\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__29369\,
            I => \c0.n5391\
        );

    \I__6741\ : Odrv12
    port map (
            O => \N__29366\,
            I => \c0.n5391\
        );

    \I__6740\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__29358\,
            I => \c0.n26_adj_1927\
        );

    \I__6738\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29349\
        );

    \I__6737\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29349\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__29349\,
            I => \r_Tx_Data_3\
        );

    \I__6735\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29342\
        );

    \I__6734\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29339\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__29342\,
            I => \r_Tx_Data_2\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__29339\,
            I => \r_Tx_Data_2\
        );

    \I__6731\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29328\
        );

    \I__6730\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29328\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__29328\,
            I => \N__29322\
        );

    \I__6728\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29318\
        );

    \I__6727\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29312\
        );

    \I__6726\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29312\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__29322\,
            I => \N__29309\
        );

    \I__6724\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29306\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__29318\,
            I => \N__29303\
        );

    \I__6722\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29300\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__29312\,
            I => \N__29297\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__29309\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__29306\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__6718\ : Odrv12
    port map (
            O => \N__29303\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__29300\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__29297\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__6715\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29283\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__29283\,
            I => \N__29279\
        );

    \I__6713\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29276\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__29279\,
            I => \N__29273\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__29276\,
            I => \c0.tx.r_Tx_Data_0\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__29273\,
            I => \c0.tx.r_Tx_Data_0\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__29268\,
            I => \c0.tx.n6051_cascade_\
        );

    \I__6708\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29261\
        );

    \I__6707\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29258\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__29261\,
            I => \r_Tx_Data_1\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__29258\,
            I => \r_Tx_Data_1\
        );

    \I__6704\ : CascadeMux
    port map (
            O => \N__29253\,
            I => \N__29249\
        );

    \I__6703\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__6702\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29243\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29240\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29235\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__29240\,
            I => \N__29232\
        );

    \I__6698\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29229\
        );

    \I__6697\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29226\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__29235\,
            I => \N__29223\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__29232\,
            I => \N__29220\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__29229\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__29226\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__6692\ : Odrv4
    port map (
            O => \N__29223\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__29220\,
            I => \c0.tx.r_Bit_Index_2\
        );

    \I__6690\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29208\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__29208\,
            I => \c0.tx.n6054\
        );

    \I__6688\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29193\
        );

    \I__6687\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29193\
        );

    \I__6686\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29190\
        );

    \I__6685\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29185\
        );

    \I__6684\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29185\
        );

    \I__6683\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29182\
        );

    \I__6682\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29179\
        );

    \I__6681\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29176\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__29193\,
            I => \N__29170\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__29190\,
            I => \N__29167\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29164\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__29182\,
            I => \N__29161\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__29179\,
            I => \N__29156\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__29176\,
            I => \N__29156\
        );

    \I__6674\ : InMux
    port map (
            O => \N__29175\,
            I => \N__29153\
        );

    \I__6673\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29150\
        );

    \I__6672\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29147\
        );

    \I__6671\ : Span4Mux_v
    port map (
            O => \N__29170\,
            I => \N__29138\
        );

    \I__6670\ : Span4Mux_v
    port map (
            O => \N__29167\,
            I => \N__29138\
        );

    \I__6669\ : Span4Mux_v
    port map (
            O => \N__29164\,
            I => \N__29138\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__29161\,
            I => \N__29138\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__29156\,
            I => \N__29135\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__29153\,
            I => \r_SM_Main_0\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__29150\,
            I => \r_SM_Main_0\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__29147\,
            I => \r_SM_Main_0\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__29138\,
            I => \r_SM_Main_0\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__29135\,
            I => \r_SM_Main_0\
        );

    \I__6661\ : CascadeMux
    port map (
            O => \N__29124\,
            I => \c0.tx.o_Tx_Serial_N_1798_cascade_\
        );

    \I__6660\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29109\
        );

    \I__6658\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29106\
        );

    \I__6657\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29101\
        );

    \I__6656\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29101\
        );

    \I__6655\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29098\
        );

    \I__6654\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29093\
        );

    \I__6653\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29093\
        );

    \I__6652\ : Span4Mux_h
    port map (
            O => \N__29109\,
            I => \N__29082\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__29106\,
            I => \N__29082\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29101\,
            I => \N__29079\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29074\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29074\
        );

    \I__6647\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29071\
        );

    \I__6646\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29067\
        );

    \I__6645\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29064\
        );

    \I__6644\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29061\
        );

    \I__6643\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29056\
        );

    \I__6642\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29056\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__29082\,
            I => \N__29053\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__29079\,
            I => \N__29050\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__29074\,
            I => \N__29045\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29045\
        );

    \I__6637\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29042\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__29067\,
            I => \r_SM_Main_1\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__29064\,
            I => \r_SM_Main_1\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__29061\,
            I => \r_SM_Main_1\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__29056\,
            I => \r_SM_Main_1\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__29053\,
            I => \r_SM_Main_1\
        );

    \I__6631\ : Odrv4
    port map (
            O => \N__29050\,
            I => \r_SM_Main_1\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__29045\,
            I => \r_SM_Main_1\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__29042\,
            I => \r_SM_Main_1\
        );

    \I__6628\ : CascadeMux
    port map (
            O => \N__29025\,
            I => \c0.tx.n12_cascade_\
        );

    \I__6627\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \N__29018\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__29021\,
            I => \N__29012\
        );

    \I__6625\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29006\
        );

    \I__6624\ : InMux
    port map (
            O => \N__29017\,
            I => \N__29001\
        );

    \I__6623\ : InMux
    port map (
            O => \N__29016\,
            I => \N__28998\
        );

    \I__6622\ : InMux
    port map (
            O => \N__29015\,
            I => \N__28993\
        );

    \I__6621\ : InMux
    port map (
            O => \N__29012\,
            I => \N__28993\
        );

    \I__6620\ : InMux
    port map (
            O => \N__29011\,
            I => \N__28986\
        );

    \I__6619\ : InMux
    port map (
            O => \N__29010\,
            I => \N__28986\
        );

    \I__6618\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28986\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__29006\,
            I => \N__28983\
        );

    \I__6616\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28980\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__29004\,
            I => \N__28970\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__29001\,
            I => \N__28965\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28998\,
            I => \N__28962\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28959\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__28986\,
            I => \N__28949\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__28983\,
            I => \N__28949\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__28980\,
            I => \N__28949\
        );

    \I__6608\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28946\
        );

    \I__6607\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28937\
        );

    \I__6606\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28937\
        );

    \I__6605\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28937\
        );

    \I__6604\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28937\
        );

    \I__6603\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28934\
        );

    \I__6602\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28925\
        );

    \I__6601\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28925\
        );

    \I__6600\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28925\
        );

    \I__6599\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28925\
        );

    \I__6598\ : Span4Mux_h
    port map (
            O => \N__28965\,
            I => \N__28922\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__28962\,
            I => \N__28917\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__28959\,
            I => \N__28917\
        );

    \I__6595\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28910\
        );

    \I__6594\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28910\
        );

    \I__6593\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28910\
        );

    \I__6592\ : Span4Mux_h
    port map (
            O => \N__28949\,
            I => \N__28907\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__28946\,
            I => \r_SM_Main_2\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__28937\,
            I => \r_SM_Main_2\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__28934\,
            I => \r_SM_Main_2\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__28925\,
            I => \r_SM_Main_2\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__28922\,
            I => \r_SM_Main_2\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__28917\,
            I => \r_SM_Main_2\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28910\,
            I => \r_SM_Main_2\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__28907\,
            I => \r_SM_Main_2\
        );

    \I__6583\ : IoInMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__6581\ : IoSpan4Mux
    port map (
            O => \N__28884\,
            I => \N__28880\
        );

    \I__6580\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28877\
        );

    \I__6579\ : Span4Mux_s0_v
    port map (
            O => \N__28880\,
            I => \N__28872\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__28877\,
            I => \N__28872\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__28872\,
            I => \N__28869\
        );

    \I__6576\ : Span4Mux_h
    port map (
            O => \N__28869\,
            I => \N__28865\
        );

    \I__6575\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28862\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__28865\,
            I => tx_o
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__28862\,
            I => tx_o
        );

    \I__6572\ : CascadeMux
    port map (
            O => \N__28857\,
            I => \N__28854\
        );

    \I__6571\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28851\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__6568\ : Span4Mux_h
    port map (
            O => \N__28845\,
            I => \N__28842\
        );

    \I__6567\ : Span4Mux_v
    port map (
            O => \N__28842\,
            I => \N__28837\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28834\
        );

    \I__6565\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28831\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__28837\,
            I => data_in_10_5
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__28834\,
            I => data_in_10_5
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__28831\,
            I => data_in_10_5
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__28824\,
            I => \N__28821\
        );

    \I__6560\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28813\
        );

    \I__6558\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28810\
        );

    \I__6557\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28807\
        );

    \I__6556\ : Odrv12
    port map (
            O => \N__28813\,
            I => data_in_9_5
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__28810\,
            I => data_in_9_5
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__28807\,
            I => data_in_9_5
        );

    \I__6553\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28796\
        );

    \I__6552\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28793\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__28796\,
            I => \N__28790\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__28793\,
            I => \N__28787\
        );

    \I__6549\ : Span4Mux_v
    port map (
            O => \N__28790\,
            I => \N__28782\
        );

    \I__6548\ : Span4Mux_v
    port map (
            O => \N__28787\,
            I => \N__28782\
        );

    \I__6547\ : Span4Mux_h
    port map (
            O => \N__28782\,
            I => \N__28778\
        );

    \I__6546\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__28778\,
            I => data_in_6_0
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__28775\,
            I => data_in_6_0
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__28770\,
            I => \N__28767\
        );

    \I__6542\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28764\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__28761\,
            I => \c0.n9\
        );

    \I__6539\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28755\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__28749\,
            I => n8_adj_1987
        );

    \I__6535\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28740\
        );

    \I__6534\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28740\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__28737\,
            I => n5400
        );

    \I__6531\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28731\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__6529\ : Odrv4
    port map (
            O => \N__28728\,
            I => \tx_data_2_N_keep\
        );

    \I__6528\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__6526\ : Span4Mux_h
    port map (
            O => \N__28719\,
            I => \N__28716\
        );

    \I__6525\ : Odrv4
    port map (
            O => \N__28716\,
            I => n5364
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28710\,
            I => \N__28706\
        );

    \I__6522\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28703\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28700\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__28703\,
            I => \N__28697\
        );

    \I__6519\ : Odrv12
    port map (
            O => \N__28700\,
            I => n5482
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__28697\,
            I => n5482
        );

    \I__6517\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__28689\,
            I => \N__28685\
        );

    \I__6515\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28682\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__28685\,
            I => n1768
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28682\,
            I => n1768
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \n5364_cascade_\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28671\
        );

    \I__6510\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28668\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__28668\,
            I => n5871
        );

    \I__6508\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28662\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__28662\,
            I => \c0.n6312\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__28659\,
            I => \N__28656\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28653\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__28653\,
            I => \tx_data_3_N_keep\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28644\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__28644\,
            I => \c0.n5853\
        );

    \I__6500\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28629\
        );

    \I__6499\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28629\
        );

    \I__6498\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28629\
        );

    \I__6497\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28622\
        );

    \I__6496\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28622\
        );

    \I__6495\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28622\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__28629\,
            I => tx_active
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__28622\,
            I => tx_active
        );

    \I__6492\ : CascadeMux
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28610\
        );

    \I__6490\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28605\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__28610\,
            I => \N__28602\
        );

    \I__6488\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28599\
        );

    \I__6487\ : CascadeMux
    port map (
            O => \N__28608\,
            I => \N__28594\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__28605\,
            I => \N__28587\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__28602\,
            I => \N__28587\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28587\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__28598\,
            I => \N__28584\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28580\
        );

    \I__6481\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28577\
        );

    \I__6480\ : Span4Mux_v
    port map (
            O => \N__28587\,
            I => \N__28574\
        );

    \I__6479\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28567\
        );

    \I__6478\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28567\
        );

    \I__6477\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28567\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__28577\,
            I => \c0.tx_transmit\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__28574\,
            I => \c0.tx_transmit\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__28567\,
            I => \c0.tx_transmit\
        );

    \I__6473\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__28554\,
            I => n135
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__28551\,
            I => \n4_adj_1986_cascade_\
        );

    \I__6469\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28544\
        );

    \I__6468\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28541\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28538\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__28541\,
            I => data_out_19_6
        );

    \I__6465\ : Odrv12
    port map (
            O => \N__28538\,
            I => data_out_19_6
        );

    \I__6464\ : CascadeMux
    port map (
            O => \N__28533\,
            I => \N__28529\
        );

    \I__6463\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28526\
        );

    \I__6462\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28523\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__28526\,
            I => data_out_19_5
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__28523\,
            I => data_out_19_5
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__28518\,
            I => \N__28514\
        );

    \I__6458\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28509\
        );

    \I__6457\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28509\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__28509\,
            I => n5440
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__28506\,
            I => \n5_cascade_\
        );

    \I__6454\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28500\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__28500\,
            I => \c0.tx_active_prev\
        );

    \I__6452\ : InMux
    port map (
            O => \N__28497\,
            I => \N__28490\
        );

    \I__6451\ : InMux
    port map (
            O => \N__28496\,
            I => \N__28490\
        );

    \I__6450\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28487\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28482\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__28487\,
            I => \N__28479\
        );

    \I__6447\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28472\
        );

    \I__6446\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28472\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__28482\,
            I => \N__28469\
        );

    \I__6444\ : Span4Mux_h
    port map (
            O => \N__28479\,
            I => \N__28466\
        );

    \I__6443\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28461\
        );

    \I__6442\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28461\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__28472\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__28469\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__28466\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__28461\,
            I => \c0.tx.r_SM_Main_2_N_1767_1\
        );

    \I__6437\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28449\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__28446\,
            I => \c0.tx.n2177\
        );

    \I__6434\ : CascadeMux
    port map (
            O => \N__28443\,
            I => \n4333_cascade_\
        );

    \I__6433\ : CascadeMux
    port map (
            O => \N__28440\,
            I => \c0.n81_adj_1872_cascade_\
        );

    \I__6432\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28429\
        );

    \I__6430\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28426\
        );

    \I__6429\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28423\
        );

    \I__6428\ : Span4Mux_v
    port map (
            O => \N__28429\,
            I => \N__28420\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__28426\,
            I => \N__28416\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28413\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__28420\,
            I => \N__28410\
        );

    \I__6424\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28407\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28402\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__28413\,
            I => \N__28402\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__28410\,
            I => data_in_2_0
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__28407\,
            I => data_in_2_0
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__28402\,
            I => data_in_2_0
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \N__28392\
        );

    \I__6417\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28388\
        );

    \I__6416\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28385\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28382\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__28379\,
            I => \N__28373\
        );

    \I__6411\ : Span4Mux_h
    port map (
            O => \N__28376\,
            I => \N__28368\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__28373\,
            I => \N__28368\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__28368\,
            I => \N__28364\
        );

    \I__6408\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28361\
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__28364\,
            I => data_in_13_2
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__28361\,
            I => data_in_13_2
        );

    \I__6405\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__6403\ : Span4Mux_v
    port map (
            O => \N__28350\,
            I => \N__28345\
        );

    \I__6402\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28340\
        );

    \I__6401\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28340\
        );

    \I__6400\ : Sp12to4
    port map (
            O => \N__28345\,
            I => \N__28333\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28333\
        );

    \I__6398\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28329\
        );

    \I__6397\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28326\
        );

    \I__6396\ : Span12Mux_s10_h
    port map (
            O => \N__28333\,
            I => \N__28323\
        );

    \I__6395\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28320\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__28329\,
            I => \c0.data_in_field_88\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__28326\,
            I => \c0.data_in_field_88\
        );

    \I__6392\ : Odrv12
    port map (
            O => \N__28323\,
            I => \c0.data_in_field_88\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__28320\,
            I => \c0.data_in_field_88\
        );

    \I__6390\ : CascadeMux
    port map (
            O => \N__28311\,
            I => \N__28307\
        );

    \I__6389\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28303\
        );

    \I__6388\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28300\
        );

    \I__6387\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28296\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__28303\,
            I => \N__28291\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__28300\,
            I => \N__28291\
        );

    \I__6384\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28288\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28285\
        );

    \I__6382\ : Span4Mux_s3_h
    port map (
            O => \N__28291\,
            I => \N__28282\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28278\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__28285\,
            I => \N__28274\
        );

    \I__6379\ : Span4Mux_h
    port map (
            O => \N__28282\,
            I => \N__28271\
        );

    \I__6378\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28267\
        );

    \I__6377\ : Span4Mux_h
    port map (
            O => \N__28278\,
            I => \N__28264\
        );

    \I__6376\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28261\
        );

    \I__6375\ : Span4Mux_h
    port map (
            O => \N__28274\,
            I => \N__28258\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__28271\,
            I => \N__28255\
        );

    \I__6373\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28252\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__28267\,
            I => \c0.data_in_field_98\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__28264\,
            I => \c0.data_in_field_98\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__28261\,
            I => \c0.data_in_field_98\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__28258\,
            I => \c0.data_in_field_98\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__28255\,
            I => \c0.data_in_field_98\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__28252\,
            I => \c0.data_in_field_98\
        );

    \I__6366\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28235\
        );

    \I__6365\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28231\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28228\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__28234\,
            I => \N__28225\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28221\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__28228\,
            I => \N__28218\
        );

    \I__6360\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28215\
        );

    \I__6359\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28212\
        );

    \I__6358\ : Span4Mux_v
    port map (
            O => \N__28221\,
            I => \N__28209\
        );

    \I__6357\ : Span4Mux_h
    port map (
            O => \N__28218\,
            I => \N__28204\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__28215\,
            I => \N__28204\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__28212\,
            I => \c0.data_in_field_28\
        );

    \I__6354\ : Odrv4
    port map (
            O => \N__28209\,
            I => \c0.data_in_field_28\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__28204\,
            I => \c0.data_in_field_28\
        );

    \I__6352\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28192\
        );

    \I__6351\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28189\
        );

    \I__6350\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28185\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28182\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__28189\,
            I => \N__28179\
        );

    \I__6347\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28176\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28173\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__28182\,
            I => \N__28170\
        );

    \I__6344\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28165\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28162\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__28173\,
            I => \N__28157\
        );

    \I__6341\ : Span4Mux_h
    port map (
            O => \N__28170\,
            I => \N__28157\
        );

    \I__6340\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28152\
        );

    \I__6339\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28152\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__28165\,
            I => \c0.data_in_field_121\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__28162\,
            I => \c0.data_in_field_121\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__28157\,
            I => \c0.data_in_field_121\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__28152\,
            I => \c0.data_in_field_121\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__6333\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28137\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__28134\,
            I => \c0.n23_adj_1935\
        );

    \I__6330\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28127\
        );

    \I__6329\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28123\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28118\
        );

    \I__6327\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28115\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__28123\,
            I => \N__28111\
        );

    \I__6325\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28108\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__28121\,
            I => \N__28105\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__28118\,
            I => \N__28100\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__28115\,
            I => \N__28100\
        );

    \I__6321\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28097\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__28111\,
            I => \N__28093\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28090\
        );

    \I__6318\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28087\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__28100\,
            I => \N__28082\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__28097\,
            I => \N__28082\
        );

    \I__6315\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28079\
        );

    \I__6314\ : Span4Mux_h
    port map (
            O => \N__28093\,
            I => \N__28074\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__28090\,
            I => \N__28074\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__28087\,
            I => \c0.data_in_field_87\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__28082\,
            I => \c0.data_in_field_87\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__28079\,
            I => \c0.data_in_field_87\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__28074\,
            I => \c0.data_in_field_87\
        );

    \I__6308\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28062\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__6306\ : Span4Mux_v
    port map (
            O => \N__28059\,
            I => \N__28055\
        );

    \I__6305\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28052\
        );

    \I__6304\ : Sp12to4
    port map (
            O => \N__28055\,
            I => \N__28049\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__28052\,
            I => \N__28046\
        );

    \I__6302\ : Span12Mux_s10_h
    port map (
            O => \N__28049\,
            I => \N__28040\
        );

    \I__6301\ : Span4Mux_v
    port map (
            O => \N__28046\,
            I => \N__28037\
        );

    \I__6300\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28032\
        );

    \I__6299\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28032\
        );

    \I__6298\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28029\
        );

    \I__6297\ : Odrv12
    port map (
            O => \N__28040\,
            I => \c0.data_in_field_128\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__28037\,
            I => \c0.data_in_field_128\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__28032\,
            I => \c0.data_in_field_128\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__28029\,
            I => \c0.data_in_field_128\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__28013\
        );

    \I__6291\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28010\
        );

    \I__6290\ : Odrv12
    port map (
            O => \N__28013\,
            I => \c0.n2068\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__28010\,
            I => \c0.n2068\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27998\
        );

    \I__6286\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27995\
        );

    \I__6285\ : Span4Mux_h
    port map (
            O => \N__27998\,
            I => \N__27991\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27988\
        );

    \I__6283\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27983\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__27991\,
            I => \N__27980\
        );

    \I__6281\ : Span4Mux_h
    port map (
            O => \N__27988\,
            I => \N__27977\
        );

    \I__6280\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27974\
        );

    \I__6279\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27971\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27983\,
            I => \c0.data_in_field_46\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__27980\,
            I => \c0.data_in_field_46\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__27977\,
            I => \c0.data_in_field_46\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__27974\,
            I => \c0.data_in_field_46\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__27971\,
            I => \c0.data_in_field_46\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__27960\,
            I => \c0.n1965_cascade_\
        );

    \I__6272\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27954\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__27954\,
            I => \N__27948\
        );

    \I__6270\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27945\
        );

    \I__6269\ : InMux
    port map (
            O => \N__27952\,
            I => \N__27942\
        );

    \I__6268\ : InMux
    port map (
            O => \N__27951\,
            I => \N__27937\
        );

    \I__6267\ : Span4Mux_h
    port map (
            O => \N__27948\,
            I => \N__27934\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__27945\,
            I => \N__27931\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27928\
        );

    \I__6264\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27923\
        );

    \I__6263\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27923\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27916\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__27934\,
            I => \N__27916\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__27931\,
            I => \N__27916\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__27928\,
            I => \c0.data_in_field_91\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__27923\,
            I => \c0.data_in_field_91\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__27916\,
            I => \c0.data_in_field_91\
        );

    \I__6256\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27906\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__27906\,
            I => \N__27903\
        );

    \I__6254\ : Odrv4
    port map (
            O => \N__27903\,
            I => \c0.n24_adj_1930\
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__27900\,
            I => \N__27897\
        );

    \I__6252\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27893\
        );

    \I__6251\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27890\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27893\,
            I => \N__27886\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__27890\,
            I => \N__27883\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27889\,
            I => \N__27879\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__27886\,
            I => \N__27876\
        );

    \I__6246\ : Span12Mux_s10_h
    port map (
            O => \N__27883\,
            I => \N__27873\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27870\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__27879\,
            I => data_in_3_5
        );

    \I__6243\ : Odrv4
    port map (
            O => \N__27876\,
            I => data_in_3_5
        );

    \I__6242\ : Odrv12
    port map (
            O => \N__27873\,
            I => data_in_3_5
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__27870\,
            I => data_in_3_5
        );

    \I__6240\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27858\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27853\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27850\
        );

    \I__6237\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27847\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__27853\,
            I => \N__27844\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27840\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__27847\,
            I => \N__27837\
        );

    \I__6233\ : Sp12to4
    port map (
            O => \N__27844\,
            I => \N__27834\
        );

    \I__6232\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27831\
        );

    \I__6231\ : Span4Mux_h
    port map (
            O => \N__27840\,
            I => \N__27828\
        );

    \I__6230\ : Odrv4
    port map (
            O => \N__27837\,
            I => data_in_3_0
        );

    \I__6229\ : Odrv12
    port map (
            O => \N__27834\,
            I => data_in_3_0
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__27831\,
            I => data_in_3_0
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__27828\,
            I => data_in_3_0
        );

    \I__6226\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__27816\,
            I => \N__27811\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__27815\,
            I => \N__27808\
        );

    \I__6223\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27805\
        );

    \I__6222\ : Span4Mux_h
    port map (
            O => \N__27811\,
            I => \N__27802\
        );

    \I__6221\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27799\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__27805\,
            I => \N__27796\
        );

    \I__6219\ : Span4Mux_v
    port map (
            O => \N__27802\,
            I => \N__27792\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27787\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__27796\,
            I => \N__27787\
        );

    \I__6216\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27784\
        );

    \I__6215\ : Span4Mux_v
    port map (
            O => \N__27792\,
            I => \N__27781\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__27787\,
            I => \N__27778\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__27784\,
            I => data_in_2_6
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27781\,
            I => data_in_2_6
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__27778\,
            I => data_in_2_6
        );

    \I__6210\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__6208\ : Span4Mux_v
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__6207\ : Span4Mux_h
    port map (
            O => \N__27762\,
            I => \N__27759\
        );

    \I__6206\ : Odrv4
    port map (
            O => \N__27759\,
            I => \c0.n28_adj_1925\
        );

    \I__6205\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27750\
        );

    \I__6204\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27738\
        );

    \I__6203\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27738\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27735\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__27750\,
            I => \N__27732\
        );

    \I__6200\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27729\
        );

    \I__6199\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27726\
        );

    \I__6198\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27721\
        );

    \I__6197\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27721\
        );

    \I__6196\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27713\
        );

    \I__6195\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27710\
        );

    \I__6194\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27707\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27704\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27691\
        );

    \I__6191\ : Span4Mux_s2_h
    port map (
            O => \N__27732\,
            I => \N__27691\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__27729\,
            I => \N__27691\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27691\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__27721\,
            I => \N__27691\
        );

    \I__6187\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27688\
        );

    \I__6186\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27680\
        );

    \I__6185\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27677\
        );

    \I__6184\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27674\
        );

    \I__6183\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27671\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27668\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27658\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27658\
        );

    \I__6179\ : Span4Mux_v
    port map (
            O => \N__27704\,
            I => \N__27655\
        );

    \I__6178\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27652\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__27702\,
            I => \N__27649\
        );

    \I__6176\ : Span4Mux_v
    port map (
            O => \N__27691\,
            I => \N__27641\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__27688\,
            I => \N__27641\
        );

    \I__6174\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27636\
        );

    \I__6173\ : InMux
    port map (
            O => \N__27686\,
            I => \N__27636\
        );

    \I__6172\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27629\
        );

    \I__6171\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27624\
        );

    \I__6170\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27624\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27621\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27614\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27614\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27671\,
            I => \N__27614\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__27668\,
            I => \N__27609\
        );

    \I__6164\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27604\
        );

    \I__6163\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27601\
        );

    \I__6162\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27598\
        );

    \I__6161\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27595\
        );

    \I__6160\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27592\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__27658\,
            I => \N__27585\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__27655\,
            I => \N__27585\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27585\
        );

    \I__6156\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27582\
        );

    \I__6155\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27579\
        );

    \I__6154\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27574\
        );

    \I__6153\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27574\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__27641\,
            I => \N__27569\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27569\
        );

    \I__6150\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27565\
        );

    \I__6149\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27558\
        );

    \I__6148\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27558\
        );

    \I__6147\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27558\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27554\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27547\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__27621\,
            I => \N__27547\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27547\
        );

    \I__6142\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27543\
        );

    \I__6141\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27540\
        );

    \I__6140\ : Sp12to4
    port map (
            O => \N__27609\,
            I => \N__27537\
        );

    \I__6139\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27534\
        );

    \I__6138\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27531\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27528\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27517\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27517\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__27595\,
            I => \N__27517\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27517\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__27585\,
            I => \N__27517\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27514\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__27579\,
            I => \N__27507\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27507\
        );

    \I__6128\ : Span4Mux_v
    port map (
            O => \N__27569\,
            I => \N__27507\
        );

    \I__6127\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27504\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27501\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27498\
        );

    \I__6124\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27495\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__27554\,
            I => \N__27490\
        );

    \I__6122\ : Span4Mux_v
    port map (
            O => \N__27547\,
            I => \N__27490\
        );

    \I__6121\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27487\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__27543\,
            I => \N__27482\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27482\
        );

    \I__6118\ : Span12Mux_h
    port map (
            O => \N__27537\,
            I => \N__27477\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__27534\,
            I => \N__27477\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__27531\,
            I => \N__27470\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__27528\,
            I => \N__27470\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27470\
        );

    \I__6113\ : Span4Mux_v
    port map (
            O => \N__27514\,
            I => \N__27465\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__27507\,
            I => \N__27465\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__27504\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__27501\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__27498\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__27495\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__27490\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__27487\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6105\ : Odrv12
    port map (
            O => \N__27482\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6104\ : Odrv12
    port map (
            O => \N__27477\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__27470\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__27465\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__6101\ : InMux
    port map (
            O => \N__27444\,
            I => \N__27439\
        );

    \I__6100\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27436\
        );

    \I__6099\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27432\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27429\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27426\
        );

    \I__6096\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27423\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__27432\,
            I => \c0.data_in_field_24\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__27429\,
            I => \c0.data_in_field_24\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__27426\,
            I => \c0.data_in_field_24\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__27423\,
            I => \c0.data_in_field_24\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__6090\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__6088\ : Span12Mux_s1_h
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__6087\ : Odrv12
    port map (
            O => \N__27402\,
            I => \c0.n6039\
        );

    \I__6086\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27392\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__27395\,
            I => \N__27389\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__27392\,
            I => \N__27386\
        );

    \I__6082\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27383\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__27386\,
            I => \N__27380\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__27383\,
            I => \N__27376\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__27380\,
            I => \N__27373\
        );

    \I__6078\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27370\
        );

    \I__6077\ : Odrv12
    port map (
            O => \N__27376\,
            I => data_in_17_4
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__27373\,
            I => data_in_17_4
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__27370\,
            I => data_in_17_4
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__6073\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__27357\,
            I => \N__27353\
        );

    \I__6071\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27350\
        );

    \I__6070\ : Span4Mux_v
    port map (
            O => \N__27353\,
            I => \N__27347\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__27350\,
            I => \N__27344\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__27347\,
            I => \N__27340\
        );

    \I__6067\ : Span4Mux_h
    port map (
            O => \N__27344\,
            I => \N__27337\
        );

    \I__6066\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27334\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__27340\,
            I => data_in_5_4
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__27337\,
            I => data_in_5_4
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__27334\,
            I => data_in_5_4
        );

    \I__6062\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27323\
        );

    \I__6061\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27317\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27314\
        );

    \I__6058\ : Span4Mux_v
    port map (
            O => \N__27317\,
            I => \N__27311\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__27314\,
            I => \N__27306\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__27311\,
            I => \N__27306\
        );

    \I__6055\ : Span4Mux_h
    port map (
            O => \N__27306\,
            I => \N__27303\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__27303\,
            I => \c0.n5560\
        );

    \I__6053\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27296\
        );

    \I__6052\ : CascadeMux
    port map (
            O => \N__27299\,
            I => \N__27293\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27290\
        );

    \I__6050\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27287\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__27290\,
            I => \N__27281\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__27287\,
            I => \N__27278\
        );

    \I__6047\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27271\
        );

    \I__6046\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27271\
        );

    \I__6045\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27271\
        );

    \I__6044\ : Sp12to4
    port map (
            O => \N__27281\,
            I => \N__27268\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__27278\,
            I => \c0.data_in_field_106\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__27271\,
            I => \c0.data_in_field_106\
        );

    \I__6041\ : Odrv12
    port map (
            O => \N__27268\,
            I => \c0.data_in_field_106\
        );

    \I__6040\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27257\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__27260\,
            I => \N__27254\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__27257\,
            I => \N__27251\
        );

    \I__6037\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27248\
        );

    \I__6036\ : Span4Mux_v
    port map (
            O => \N__27251\,
            I => \N__27243\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27243\
        );

    \I__6034\ : Span4Mux_h
    port map (
            O => \N__27243\,
            I => \N__27238\
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__27242\,
            I => \N__27235\
        );

    \I__6032\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27231\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__27238\,
            I => \N__27228\
        );

    \I__6030\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27225\
        );

    \I__6029\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27222\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__27231\,
            I => \c0.data_in_field_2\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__27228\,
            I => \c0.data_in_field_2\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__27225\,
            I => \c0.data_in_field_2\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__27222\,
            I => \c0.data_in_field_2\
        );

    \I__6024\ : CascadeMux
    port map (
            O => \N__27213\,
            I => \c0.n5560_cascade_\
        );

    \I__6023\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__27198\,
            I => \c0.n34\
        );

    \I__6018\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__6016\ : Span4Mux_v
    port map (
            O => \N__27189\,
            I => \N__27185\
        );

    \I__6015\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27182\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__27185\,
            I => \N__27176\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__27176\
        );

    \I__6012\ : InMux
    port map (
            O => \N__27181\,
            I => \N__27173\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__27176\,
            I => data_in_5_7
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__27173\,
            I => data_in_5_7
        );

    \I__6009\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27161\
        );

    \I__6007\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27158\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__27161\,
            I => \N__27153\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__27158\,
            I => \N__27150\
        );

    \I__6004\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27145\
        );

    \I__6003\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27145\
        );

    \I__6002\ : Odrv4
    port map (
            O => \N__27153\,
            I => \c0.data_in_field_133\
        );

    \I__6001\ : Odrv12
    port map (
            O => \N__27150\,
            I => \c0.data_in_field_133\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__27145\,
            I => \c0.data_in_field_133\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27134\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__27137\,
            I => \N__27128\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27125\
        );

    \I__5996\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27120\
        );

    \I__5995\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27120\
        );

    \I__5994\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27115\
        );

    \I__5993\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27115\
        );

    \I__5992\ : Span4Mux_v
    port map (
            O => \N__27125\,
            I => \N__27112\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27109\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__27115\,
            I => \N__27104\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__27112\,
            I => \N__27104\
        );

    \I__5988\ : Odrv12
    port map (
            O => \N__27109\,
            I => \c0.data_in_field_21\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__27104\,
            I => \c0.data_in_field_21\
        );

    \I__5986\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27094\
        );

    \I__5985\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27091\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27088\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27085\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27081\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27078\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__27085\,
            I => \N__27075\
        );

    \I__5979\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27072\
        );

    \I__5978\ : Span4Mux_s3_h
    port map (
            O => \N__27081\,
            I => \N__27067\
        );

    \I__5977\ : Span4Mux_h
    port map (
            O => \N__27078\,
            I => \N__27064\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__27075\,
            I => \N__27061\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__27072\,
            I => \N__27058\
        );

    \I__5974\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27053\
        );

    \I__5973\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27053\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__27067\,
            I => \c0.data_in_field_143\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__27064\,
            I => \c0.data_in_field_143\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__27061\,
            I => \c0.data_in_field_143\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__27058\,
            I => \c0.data_in_field_143\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__27053\,
            I => \c0.data_in_field_143\
        );

    \I__5967\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27036\
        );

    \I__5965\ : Span4Mux_h
    port map (
            O => \N__27036\,
            I => \N__27033\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__27033\,
            I => \N__27029\
        );

    \I__5963\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27026\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__27029\,
            I => \c0.n5378\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__27026\,
            I => \c0.n5378\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__5959\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__27015\,
            I => \N__27011\
        );

    \I__5957\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27008\
        );

    \I__5956\ : Span4Mux_v
    port map (
            O => \N__27011\,
            I => \N__27004\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__27001\
        );

    \I__5954\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26998\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__27004\,
            I => data_in_11_5
        );

    \I__5952\ : Odrv4
    port map (
            O => \N__27001\,
            I => data_in_11_5
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__26998\,
            I => data_in_11_5
        );

    \I__5950\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26987\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__26990\,
            I => \N__26983\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__26987\,
            I => \N__26979\
        );

    \I__5947\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26974\
        );

    \I__5946\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26974\
        );

    \I__5945\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26971\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__26979\,
            I => \c0.data_in_field_55\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__26974\,
            I => \c0.data_in_field_55\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__26971\,
            I => \c0.data_in_field_55\
        );

    \I__5941\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26961\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__26961\,
            I => \N__26956\
        );

    \I__5939\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26953\
        );

    \I__5938\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26948\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__26956\,
            I => \N__26945\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26942\
        );

    \I__5935\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26937\
        );

    \I__5934\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26937\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26934\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__26945\,
            I => \c0.data_in_field_63\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__26942\,
            I => \c0.data_in_field_63\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__26937\,
            I => \c0.data_in_field_63\
        );

    \I__5929\ : Odrv12
    port map (
            O => \N__26934\,
            I => \c0.data_in_field_63\
        );

    \I__5928\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__5926\ : Span12Mux_s11_h
    port map (
            O => \N__26919\,
            I => \N__26914\
        );

    \I__5925\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26909\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26909\
        );

    \I__5923\ : Odrv12
    port map (
            O => \N__26914\,
            I => data_in_14_4
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__26909\,
            I => data_in_14_4
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__5920\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__26898\,
            I => \N__26894\
        );

    \I__5918\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26891\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__26894\,
            I => \N__26885\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26885\
        );

    \I__5915\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26882\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__26885\,
            I => \N__26879\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__26882\,
            I => \N__26874\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__26879\,
            I => \N__26871\
        );

    \I__5911\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26866\
        );

    \I__5910\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26866\
        );

    \I__5909\ : Odrv12
    port map (
            O => \N__26874\,
            I => \c0.data_in_field_48\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__26871\,
            I => \c0.data_in_field_48\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26866\,
            I => \c0.data_in_field_48\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \N__26855\
        );

    \I__5905\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26852\
        );

    \I__5904\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26849\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26845\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26842\
        );

    \I__5901\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26839\
        );

    \I__5900\ : Span4Mux_h
    port map (
            O => \N__26845\,
            I => \N__26836\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__26842\,
            I => \N__26833\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26830\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26825\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__26833\,
            I => \N__26822\
        );

    \I__5895\ : Span12Mux_s6_h
    port map (
            O => \N__26830\,
            I => \N__26819\
        );

    \I__5894\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26814\
        );

    \I__5893\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26814\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__26825\,
            I => \c0.data_in_field_32\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__26822\,
            I => \c0.data_in_field_32\
        );

    \I__5890\ : Odrv12
    port map (
            O => \N__26819\,
            I => \c0.data_in_field_32\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__26814\,
            I => \c0.data_in_field_32\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26802\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__26802\,
            I => \N__26796\
        );

    \I__5886\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26793\
        );

    \I__5885\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26790\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26786\
        );

    \I__5883\ : Span4Mux_h
    port map (
            O => \N__26796\,
            I => \N__26783\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__26793\,
            I => \N__26780\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__26790\,
            I => \N__26777\
        );

    \I__5880\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26774\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__26786\,
            I => \N__26771\
        );

    \I__5878\ : Span4Mux_h
    port map (
            O => \N__26783\,
            I => \N__26766\
        );

    \I__5877\ : Span4Mux_h
    port map (
            O => \N__26780\,
            I => \N__26766\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__26777\,
            I => \N__26763\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__26774\,
            I => \c0.data_in_field_40\
        );

    \I__5874\ : Odrv12
    port map (
            O => \N__26771\,
            I => \c0.data_in_field_40\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__26766\,
            I => \c0.data_in_field_40\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__26763\,
            I => \c0.data_in_field_40\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__26754\,
            I => \c0.n6033_cascade_\
        );

    \I__5870\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26748\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__5868\ : Span12Mux_v
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__5867\ : Odrv12
    port map (
            O => \N__26742\,
            I => \c0.n5791\
        );

    \I__5866\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26733\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__26733\,
            I => \c0.n1814\
        );

    \I__5863\ : CascadeMux
    port map (
            O => \N__26730\,
            I => \N__26727\
        );

    \I__5862\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26723\
        );

    \I__5861\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26720\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__26723\,
            I => \N__26717\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26714\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__26717\,
            I => \N__26711\
        );

    \I__5857\ : Span4Mux_h
    port map (
            O => \N__26714\,
            I => \N__26707\
        );

    \I__5856\ : Sp12to4
    port map (
            O => \N__26711\,
            I => \N__26704\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26701\
        );

    \I__5854\ : Sp12to4
    port map (
            O => \N__26707\,
            I => \N__26697\
        );

    \I__5853\ : Span12Mux_s11_h
    port map (
            O => \N__26704\,
            I => \N__26692\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__26701\,
            I => \N__26692\
        );

    \I__5851\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26689\
        );

    \I__5850\ : Span12Mux_v
    port map (
            O => \N__26697\,
            I => \N__26686\
        );

    \I__5849\ : Span12Mux_v
    port map (
            O => \N__26692\,
            I => \N__26683\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__26689\,
            I => data_in_19_1
        );

    \I__5847\ : Odrv12
    port map (
            O => \N__26686\,
            I => data_in_19_1
        );

    \I__5846\ : Odrv12
    port map (
            O => \N__26683\,
            I => data_in_19_1
        );

    \I__5845\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26672\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__26675\,
            I => \N__26669\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__26672\,
            I => \N__26666\
        );

    \I__5842\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26663\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__26666\,
            I => \N__26660\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__26663\,
            I => \N__26657\
        );

    \I__5839\ : Span4Mux_h
    port map (
            O => \N__26660\,
            I => \N__26654\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__26657\,
            I => \c0.n2143\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__26654\,
            I => \c0.n2143\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__26649\,
            I => \c0.n1814_cascade_\
        );

    \I__5835\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26639\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__26645\,
            I => \N__26636\
        );

    \I__5833\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26633\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26630\
        );

    \I__5831\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26627\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26624\
        );

    \I__5829\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26621\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__26633\,
            I => \N__26618\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__26630\,
            I => \N__26613\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__26627\,
            I => \N__26613\
        );

    \I__5825\ : Span12Mux_v
    port map (
            O => \N__26624\,
            I => \N__26608\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__26621\,
            I => \N__26605\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__26618\,
            I => \N__26600\
        );

    \I__5822\ : Span4Mux_v
    port map (
            O => \N__26613\,
            I => \N__26600\
        );

    \I__5821\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26595\
        );

    \I__5820\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26595\
        );

    \I__5819\ : Odrv12
    port map (
            O => \N__26608\,
            I => \c0.data_in_field_109\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__26605\,
            I => \c0.data_in_field_109\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__26600\,
            I => \c0.data_in_field_109\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__26595\,
            I => \c0.data_in_field_109\
        );

    \I__5815\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__26583\,
            I => \c0.n32_adj_1901\
        );

    \I__5813\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26576\
        );

    \I__5812\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26572\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__26576\,
            I => \N__26569\
        );

    \I__5810\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26566\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26561\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__26569\,
            I => \N__26561\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26558\
        );

    \I__5806\ : Sp12to4
    port map (
            O => \N__26561\,
            I => \N__26553\
        );

    \I__5805\ : Span12Mux_s11_h
    port map (
            O => \N__26558\,
            I => \N__26553\
        );

    \I__5804\ : Odrv12
    port map (
            O => \N__26553\,
            I => data_in_8_5
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__5802\ : InMux
    port map (
            O => \N__26547\,
            I => \N__26544\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__26541\,
            I => n318
        );

    \I__5799\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26534\
        );

    \I__5798\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26529\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__26534\,
            I => \N__26526\
        );

    \I__5796\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26523\
        );

    \I__5795\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26520\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__26529\,
            I => \r_Clock_Count_3\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__26526\,
            I => \r_Clock_Count_3\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__26523\,
            I => \r_Clock_Count_3\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__26520\,
            I => \r_Clock_Count_3\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__5789\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__26502\,
            I => n321
        );

    \I__5786\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__26496\,
            I => \N__26490\
        );

    \I__5784\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26485\
        );

    \I__5783\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26485\
        );

    \I__5782\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26482\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__26490\,
            I => \r_Clock_Count_0\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__26485\,
            I => \r_Clock_Count_0\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__26482\,
            I => \r_Clock_Count_0\
        );

    \I__5778\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26471\
        );

    \I__5777\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26468\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__26471\,
            I => \N__26465\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__26468\,
            I => data_out_18_5
        );

    \I__5774\ : Odrv12
    port map (
            O => \N__26465\,
            I => data_out_18_5
        );

    \I__5773\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26451\
        );

    \I__5772\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26451\
        );

    \I__5771\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26446\
        );

    \I__5770\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26446\
        );

    \I__5769\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26443\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__26451\,
            I => n782
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__26446\,
            I => n782
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__26443\,
            I => n782
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__26436\,
            I => \N__26433\
        );

    \I__5764\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26430\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__26430\,
            I => \N__26427\
        );

    \I__5762\ : Span4Mux_h
    port map (
            O => \N__26427\,
            I => \N__26424\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__26424\,
            I => n320
        );

    \I__5760\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__26418\,
            I => \N__26414\
        );

    \I__5758\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26409\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__26414\,
            I => \N__26406\
        );

    \I__5756\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26403\
        );

    \I__5755\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26400\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__26409\,
            I => \r_Clock_Count_1\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__26406\,
            I => \r_Clock_Count_1\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__26403\,
            I => \r_Clock_Count_1\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__26400\,
            I => \r_Clock_Count_1\
        );

    \I__5750\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26387\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__26390\,
            I => \N__26384\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26381\
        );

    \I__5747\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26378\
        );

    \I__5746\ : Odrv12
    port map (
            O => \N__26381\,
            I => rx_data_1
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__26378\,
            I => rx_data_1
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__5743\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__26367\,
            I => \N__26363\
        );

    \I__5741\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26360\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__26363\,
            I => \N__26357\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26354\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__26357\,
            I => \N__26350\
        );

    \I__5737\ : Span12Mux_h
    port map (
            O => \N__26354\,
            I => \N__26347\
        );

    \I__5736\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26344\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__26350\,
            I => data_in_14_3
        );

    \I__5734\ : Odrv12
    port map (
            O => \N__26347\,
            I => data_in_14_3
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__26344\,
            I => data_in_14_3
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__5731\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26330\
        );

    \I__5730\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26327\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__26330\,
            I => \N__26322\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26327\,
            I => \N__26322\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__26322\,
            I => \N__26318\
        );

    \I__5726\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26315\
        );

    \I__5725\ : Span4Mux_h
    port map (
            O => \N__26318\,
            I => \N__26312\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__26315\,
            I => data_in_13_3
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__26312\,
            I => data_in_13_3
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__26307\,
            I => \c0.n6309_cascade_\
        );

    \I__5721\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26298\
        );

    \I__5720\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26298\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__26298\,
            I => data_out_18_2
        );

    \I__5718\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26292\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__26292\,
            I => \c0.n1249\
        );

    \I__5716\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26286\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__26286\,
            I => \N__26283\
        );

    \I__5714\ : Odrv12
    port map (
            O => \N__26283\,
            I => \tx_data_4_N_keep\
        );

    \I__5713\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26277\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__26277\,
            I => \c0.tx.n3644\
        );

    \I__5711\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26271\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__26271\,
            I => n11_adj_1979
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__26268\,
            I => \n5818_cascade_\
        );

    \I__5708\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26262\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26259\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__26259\,
            I => n4155
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__26256\,
            I => \n4334_cascade_\
        );

    \I__5704\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__26250\,
            I => n1991
        );

    \I__5702\ : InMux
    port map (
            O => \N__26247\,
            I => \N__26243\
        );

    \I__5701\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26240\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__26243\,
            I => data_out_19_7
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__26240\,
            I => data_out_19_7
        );

    \I__5698\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__26232\,
            I => \c0.n17_adj_1950\
        );

    \I__5696\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__26226\,
            I => n4_adj_1982
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__26223\,
            I => \N__26220\
        );

    \I__5693\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26217\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__26217\,
            I => \c0.n17_adj_1908\
        );

    \I__5691\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26210\
        );

    \I__5690\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26207\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__26210\,
            I => data_out_18_7
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__26207\,
            I => data_out_18_7
        );

    \I__5687\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26195\
        );

    \I__5686\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26195\
        );

    \I__5685\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26192\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__26195\,
            I => \c0.n1508\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__26192\,
            I => \c0.n1508\
        );

    \I__5682\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26183\
        );

    \I__5681\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26180\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26177\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__26180\,
            I => data_out_19_2
        );

    \I__5678\ : Odrv4
    port map (
            O => \N__26177\,
            I => data_out_19_2
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__26172\,
            I => \c0.n1508_cascade_\
        );

    \I__5676\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26166\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__26166\,
            I => \c0.n5840\
        );

    \I__5674\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26159\
        );

    \I__5673\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26155\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__26159\,
            I => \N__26152\
        );

    \I__5671\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26149\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__26155\,
            I => \N__26146\
        );

    \I__5669\ : Span4Mux_v
    port map (
            O => \N__26152\,
            I => \N__26143\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__26149\,
            I => data_in_11_7
        );

    \I__5667\ : Odrv12
    port map (
            O => \N__26146\,
            I => data_in_11_7
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__26143\,
            I => data_in_11_7
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__26136\,
            I => \n5448_cascade_\
        );

    \I__5664\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26130\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26130\,
            I => \N__26127\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__26127\,
            I => n4_adj_1975
        );

    \I__5661\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26120\
        );

    \I__5660\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26117\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__26120\,
            I => data_out_19_4
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__26117\,
            I => data_out_19_4
        );

    \I__5657\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26106\
        );

    \I__5656\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26106\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__26106\,
            I => data_out_18_4
        );

    \I__5654\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26100\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__26100\,
            I => \N__26096\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26093\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__26096\,
            I => \N__26090\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__26093\,
            I => \c0.delay_counter_3\
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__26090\,
            I => \c0.delay_counter_3\
        );

    \I__5648\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__26082\,
            I => \N__26078\
        );

    \I__5646\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26075\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__26078\,
            I => \N__26072\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__26075\,
            I => \c0.delay_counter_6\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__26072\,
            I => \c0.delay_counter_6\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__5641\ : InMux
    port map (
            O => \N__26064\,
            I => \N__26060\
        );

    \I__5640\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26057\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__26060\,
            I => \N__26054\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__26057\,
            I => \c0.delay_counter_10\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__26054\,
            I => \c0.delay_counter_10\
        );

    \I__5636\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26046\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__26046\,
            I => \c0.n18_adj_1919\
        );

    \I__5634\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26040\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__26040\,
            I => \N__26036\
        );

    \I__5632\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26033\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__26036\,
            I => \N__26030\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__26033\,
            I => \c0.delay_counter_8\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__26030\,
            I => \c0.delay_counter_8\
        );

    \I__5628\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26022\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__26018\
        );

    \I__5626\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26015\
        );

    \I__5625\ : Span4Mux_v
    port map (
            O => \N__26018\,
            I => \N__26012\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__26015\,
            I => \c0.delay_counter_4\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__26012\,
            I => \c0.delay_counter_4\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__26007\,
            I => \c0.n20_adj_1922_cascade_\
        );

    \I__5621\ : InMux
    port map (
            O => \N__26004\,
            I => \N__26001\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__26001\,
            I => \N__25998\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__25998\,
            I => \c0.n16_adj_1921\
        );

    \I__5618\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25991\
        );

    \I__5617\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25988\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25985\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25979\
        );

    \I__5614\ : Span4Mux_v
    port map (
            O => \N__25985\,
            I => \N__25976\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__25984\,
            I => \N__25973\
        );

    \I__5612\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25970\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25967\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__25979\,
            I => \N__25962\
        );

    \I__5609\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25962\
        );

    \I__5608\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25959\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__25970\,
            I => \c0.data_in_field_77\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25967\,
            I => \c0.data_in_field_77\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__25962\,
            I => \c0.data_in_field_77\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__25959\,
            I => \c0.data_in_field_77\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__25950\,
            I => \c0.n6207_cascade_\
        );

    \I__5602\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25943\
        );

    \I__5601\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25940\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25937\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25940\,
            I => \N__25931\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__25937\,
            I => \N__25928\
        );

    \I__5597\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25921\
        );

    \I__5596\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25921\
        );

    \I__5595\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25921\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__25931\,
            I => \c0.data_in_field_69\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__25928\,
            I => \c0.data_in_field_69\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__25921\,
            I => \c0.data_in_field_69\
        );

    \I__5591\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25911\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__25911\,
            I => \c0.n5713\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__25908\,
            I => \N__25905\
        );

    \I__5588\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25902\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25898\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__25901\,
            I => \N__25895\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__25898\,
            I => \N__25890\
        );

    \I__5584\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25887\
        );

    \I__5583\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25882\
        );

    \I__5582\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25882\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__25890\,
            I => \N__25879\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__25887\,
            I => \N__25876\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__25882\,
            I => data_in_19_2
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__25879\,
            I => data_in_19_2
        );

    \I__5577\ : Odrv12
    port map (
            O => \N__25876\,
            I => data_in_19_2
        );

    \I__5576\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25865\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__25868\,
            I => \N__25862\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__25865\,
            I => \N__25858\
        );

    \I__5573\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25855\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25852\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__25858\,
            I => \N__25849\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__25855\,
            I => data_in_9_0
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__25852\,
            I => data_in_9_0
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__25849\,
            I => data_in_9_0
        );

    \I__5567\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__25839\,
            I => \N__25836\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__25836\,
            I => \N__25832\
        );

    \I__5564\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25829\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__25832\,
            I => \N__25825\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__25829\,
            I => \N__25822\
        );

    \I__5561\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25818\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__25825\,
            I => \N__25813\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__25822\,
            I => \N__25813\
        );

    \I__5558\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25810\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__25818\,
            I => \c0.data_in_field_42\
        );

    \I__5556\ : Odrv4
    port map (
            O => \N__25813\,
            I => \c0.data_in_field_42\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__25810\,
            I => \c0.data_in_field_42\
        );

    \I__5554\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__25800\,
            I => \N__25797\
        );

    \I__5552\ : Span4Mux_s2_h
    port map (
            O => \N__25797\,
            I => \N__25794\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__25794\,
            I => \N__25790\
        );

    \I__5550\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25784\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__5548\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25776\
        );

    \I__5547\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25776\
        );

    \I__5546\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25773\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__25784\,
            I => \c0.data_in_field_72\
        );

    \I__5544\ : Odrv4
    port map (
            O => \N__25781\,
            I => \c0.data_in_field_72\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__25776\,
            I => \c0.data_in_field_72\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__25773\,
            I => \c0.data_in_field_72\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25761\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25757\
        );

    \I__5539\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25753\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__25757\,
            I => \N__25750\
        );

    \I__5537\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25747\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25744\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__25750\,
            I => \N__25741\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__25747\,
            I => data_in_12_0
        );

    \I__5533\ : Odrv12
    port map (
            O => \N__25744\,
            I => data_in_12_0
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__25741\,
            I => data_in_12_0
        );

    \I__5531\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25728\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__25728\,
            I => \N__25724\
        );

    \I__5528\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25721\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__25724\,
            I => \N__25716\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__25721\,
            I => \N__25716\
        );

    \I__5525\ : Span4Mux_v
    port map (
            O => \N__25716\,
            I => \N__25711\
        );

    \I__5524\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25708\
        );

    \I__5523\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25705\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__25711\,
            I => \N__25702\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__25708\,
            I => data_in_18_2
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__25705\,
            I => data_in_18_2
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__25702\,
            I => data_in_18_2
        );

    \I__5518\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25692\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__25692\,
            I => \N__25688\
        );

    \I__5516\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25685\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__25688\,
            I => \N__25682\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25679\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__25682\,
            I => \N__25674\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__25679\,
            I => \N__25674\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__25674\,
            I => \N__25670\
        );

    \I__5510\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__25670\,
            I => data_in_17_2
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25667\,
            I => data_in_17_2
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__25662\,
            I => \N__25658\
        );

    \I__5506\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25655\
        );

    \I__5505\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25652\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__25655\,
            I => \N__25647\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__25652\,
            I => \N__25647\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__25644\,
            I => \N__25640\
        );

    \I__5500\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__25640\,
            I => \N__25634\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__25637\,
            I => data_in_6_2
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__25634\,
            I => data_in_6_2
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__25629\,
            I => \N__25625\
        );

    \I__5495\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25622\
        );

    \I__5494\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25619\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25616\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25612\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__25616\,
            I => \N__25609\
        );

    \I__5490\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25606\
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__25612\,
            I => data_in_5_2
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__25609\,
            I => data_in_5_2
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__25606\,
            I => data_in_5_2
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__5485\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25592\
        );

    \I__5484\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25584\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__25589\,
            I => \N__25584\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__25584\,
            I => \N__25580\
        );

    \I__5480\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25577\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__25580\,
            I => data_in_4_5
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__25577\,
            I => data_in_4_5
        );

    \I__5477\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25565\
        );

    \I__5475\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25562\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__25565\,
            I => \N__25559\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__25562\,
            I => \N__25556\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__25559\,
            I => \N__25550\
        );

    \I__5471\ : Span4Mux_v
    port map (
            O => \N__25556\,
            I => \N__25550\
        );

    \I__5470\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25547\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__25550\,
            I => \N__25544\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__25547\,
            I => \N__25539\
        );

    \I__5467\ : Sp12to4
    port map (
            O => \N__25544\,
            I => \N__25536\
        );

    \I__5466\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25531\
        );

    \I__5465\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25531\
        );

    \I__5464\ : Odrv12
    port map (
            O => \N__25539\,
            I => \c0.data_in_field_120\
        );

    \I__5463\ : Odrv12
    port map (
            O => \N__25536\,
            I => \c0.data_in_field_120\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__25531\,
            I => \c0.data_in_field_120\
        );

    \I__5461\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__25518\,
            I => \N__25514\
        );

    \I__5458\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25511\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25505\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__25508\,
            I => \c0.n2107\
        );

    \I__5454\ : Odrv12
    port map (
            O => \N__25505\,
            I => \c0.n2107\
        );

    \I__5453\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__25497\,
            I => \N__25493\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__25496\,
            I => \N__25490\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__5449\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25484\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__25487\,
            I => rx_data_2
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__25484\,
            I => rx_data_2
        );

    \I__5446\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__5444\ : Span4Mux_v
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__25467\,
            I => \c0.n6201\
        );

    \I__5441\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25459\
        );

    \I__5440\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25456\
        );

    \I__5439\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25451\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__25459\,
            I => \N__25448\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25445\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__25455\,
            I => \N__25442\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__25454\,
            I => \N__25438\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25435\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__25448\,
            I => \N__25430\
        );

    \I__5432\ : Span4Mux_h
    port map (
            O => \N__25445\,
            I => \N__25430\
        );

    \I__5431\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25427\
        );

    \I__5430\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25422\
        );

    \I__5429\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25422\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__25435\,
            I => \c0.data_in_field_101\
        );

    \I__5427\ : Odrv4
    port map (
            O => \N__25430\,
            I => \c0.data_in_field_101\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__25427\,
            I => \c0.data_in_field_101\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__25422\,
            I => \c0.data_in_field_101\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__5423\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25399\
        );

    \I__5422\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25396\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__25408\,
            I => \N__25393\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__25407\,
            I => \N__25387\
        );

    \I__5419\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25383\
        );

    \I__5418\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25376\
        );

    \I__5417\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25376\
        );

    \I__5416\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25373\
        );

    \I__5415\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25369\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25364\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__25396\,
            I => \N__25364\
        );

    \I__5412\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25361\
        );

    \I__5411\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25358\
        );

    \I__5410\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25355\
        );

    \I__5409\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25350\
        );

    \I__5408\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25350\
        );

    \I__5407\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25347\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__25383\,
            I => \N__25344\
        );

    \I__5405\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25339\
        );

    \I__5404\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25339\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__25376\,
            I => \N__25336\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25333\
        );

    \I__5401\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25330\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__25369\,
            I => \N__25327\
        );

    \I__5399\ : Span4Mux_h
    port map (
            O => \N__25364\,
            I => \N__25324\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__25361\,
            I => \N__25321\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25316\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__25355\,
            I => \N__25316\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25307\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25307\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__25344\,
            I => \N__25307\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25307\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25298\
        );

    \I__5390\ : Span4Mux_s3_h
    port map (
            O => \N__25333\,
            I => \N__25298\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__25330\,
            I => \N__25298\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__25327\,
            I => \N__25295\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__25324\,
            I => \N__25292\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__25321\,
            I => \N__25285\
        );

    \I__5385\ : Span4Mux_s1_h
    port map (
            O => \N__25316\,
            I => \N__25285\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__25307\,
            I => \N__25285\
        );

    \I__5383\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25282\
        );

    \I__5382\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25279\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__25298\,
            I => \N__25276\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__25295\,
            I => \N__25269\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__25292\,
            I => \N__25269\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__25285\,
            I => \N__25269\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__25282\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__25279\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__25276\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__5374\ : Odrv4
    port map (
            O => \N__25269\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__5373\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25253\
        );

    \I__5372\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25249\
        );

    \I__5371\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25244\
        );

    \I__5370\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25239\
        );

    \I__5369\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25239\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25235\
        );

    \I__5367\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25232\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__25249\,
            I => \N__25228\
        );

    \I__5365\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25225\
        );

    \I__5364\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25222\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25219\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25216\
        );

    \I__5361\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25213\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__25235\,
            I => \N__25210\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25207\
        );

    \I__5358\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25204\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__25228\,
            I => \N__25201\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__25225\,
            I => \N__25198\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25195\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__25219\,
            I => \N__25190\
        );

    \I__5353\ : Span4Mux_s2_h
    port map (
            O => \N__25216\,
            I => \N__25190\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__25213\,
            I => \N__25185\
        );

    \I__5351\ : Span4Mux_v
    port map (
            O => \N__25210\,
            I => \N__25185\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__25207\,
            I => \N__25182\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25173\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__25201\,
            I => \N__25173\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__25198\,
            I => \N__25173\
        );

    \I__5346\ : Span4Mux_s3_h
    port map (
            O => \N__25195\,
            I => \N__25173\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__25190\,
            I => \N__25170\
        );

    \I__5344\ : Odrv4
    port map (
            O => \N__25185\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__25182\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__25173\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__5341\ : Odrv4
    port map (
            O => \N__25170\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__5340\ : CascadeMux
    port map (
            O => \N__25161\,
            I => \c0.n5716_cascade_\
        );

    \I__5339\ : InMux
    port map (
            O => \N__25158\,
            I => \N__25155\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__25155\,
            I => \c0.n6195\
        );

    \I__5337\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25149\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__25149\,
            I => \N__25145\
        );

    \I__5335\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25141\
        );

    \I__5334\ : Span4Mux_v
    port map (
            O => \N__25145\,
            I => \N__25138\
        );

    \I__5333\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25135\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__25141\,
            I => \N__25131\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__25138\,
            I => \N__25126\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25126\
        );

    \I__5329\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25123\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__25131\,
            I => \N__25118\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__25126\,
            I => \N__25118\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__25123\,
            I => \c0.data_in_field_85\
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__25118\,
            I => \c0.data_in_field_85\
        );

    \I__5324\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25109\
        );

    \I__5323\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25106\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25101\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__25106\,
            I => \N__25098\
        );

    \I__5320\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25095\
        );

    \I__5319\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25091\
        );

    \I__5318\ : Span4Mux_h
    port map (
            O => \N__25101\,
            I => \N__25088\
        );

    \I__5317\ : Span12Mux_s3_h
    port map (
            O => \N__25098\,
            I => \N__25085\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25082\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25079\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__25091\,
            I => \c0.data_in_field_93\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__25088\,
            I => \c0.data_in_field_93\
        );

    \I__5312\ : Odrv12
    port map (
            O => \N__25085\,
            I => \c0.data_in_field_93\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__25082\,
            I => \c0.data_in_field_93\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25079\,
            I => \c0.data_in_field_93\
        );

    \I__5309\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__25065\,
            I => \c0.n37\
        );

    \I__5307\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__25055\
        );

    \I__5305\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25052\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__25055\,
            I => \N__25049\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25046\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__25049\,
            I => \N__25039\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__25046\,
            I => \N__25039\
        );

    \I__5300\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25036\
        );

    \I__5299\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25033\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__25039\,
            I => data_in_1_5
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__25036\,
            I => data_in_1_5
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__25033\,
            I => data_in_1_5
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__25026\,
            I => \N__25022\
        );

    \I__5294\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25019\
        );

    \I__5293\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25014\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25019\,
            I => \N__25011\
        );

    \I__5291\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25006\
        );

    \I__5290\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25006\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__25014\,
            I => \c0.data_in_field_13\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__25011\,
            I => \c0.data_in_field_13\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__25006\,
            I => \c0.data_in_field_13\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__5285\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__24993\,
            I => \c0.n6_adj_1939\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__24984\,
            I => \N__24979\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24974\
        );

    \I__5279\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24974\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__24979\,
            I => data_in_12_4
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__24974\,
            I => data_in_12_4
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__5275\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__24960\,
            I => \N__24955\
        );

    \I__5272\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24952\
        );

    \I__5271\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24949\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__24955\,
            I => data_in_11_4
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__24952\,
            I => data_in_11_4
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__24949\,
            I => data_in_11_4
        );

    \I__5267\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24939\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__24939\,
            I => \N__24936\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__24936\,
            I => \N__24933\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__24930\,
            I => \c0.n2089\
        );

    \I__5262\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__5260\ : Odrv12
    port map (
            O => \N__24921\,
            I => \c0.n2074\
        );

    \I__5259\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24915\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__24915\,
            I => \N__24911\
        );

    \I__5257\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24908\
        );

    \I__5256\ : Span12Mux_s6_h
    port map (
            O => \N__24911\,
            I => \N__24905\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24902\
        );

    \I__5254\ : Odrv12
    port map (
            O => \N__24905\,
            I => \c0.n5581\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__24902\,
            I => \c0.n5581\
        );

    \I__5252\ : InMux
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__24894\,
            I => \N__24891\
        );

    \I__5250\ : Span4Mux_v
    port map (
            O => \N__24891\,
            I => \N__24887\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24883\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__24887\,
            I => \N__24880\
        );

    \I__5247\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24877\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__24883\,
            I => \c0.data_in_field_44\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__24880\,
            I => \c0.data_in_field_44\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__24877\,
            I => \c0.data_in_field_44\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24865\
        );

    \I__5242\ : InMux
    port map (
            O => \N__24869\,
            I => \N__24862\
        );

    \I__5241\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24858\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24855\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__24862\,
            I => \N__24852\
        );

    \I__5238\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24849\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__24858\,
            I => \N__24846\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__24855\,
            I => \N__24842\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__24852\,
            I => \N__24839\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24836\
        );

    \I__5233\ : Span4Mux_v
    port map (
            O => \N__24846\,
            I => \N__24833\
        );

    \I__5232\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24829\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__24842\,
            I => \N__24826\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__24839\,
            I => \N__24819\
        );

    \I__5229\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24819\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__24833\,
            I => \N__24819\
        );

    \I__5227\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24816\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__24829\,
            I => \c0.data_in_field_100\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__24826\,
            I => \c0.data_in_field_100\
        );

    \I__5224\ : Odrv4
    port map (
            O => \N__24819\,
            I => \c0.data_in_field_100\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__24816\,
            I => \c0.data_in_field_100\
        );

    \I__5222\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24803\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24799\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24796\
        );

    \I__5219\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24793\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__24799\,
            I => \N__24789\
        );

    \I__5217\ : Span4Mux_h
    port map (
            O => \N__24796\,
            I => \N__24786\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__24793\,
            I => \N__24783\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24792\,
            I => \N__24778\
        );

    \I__5214\ : Span12Mux_s9_v
    port map (
            O => \N__24789\,
            I => \N__24775\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__24786\,
            I => \N__24772\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__24783\,
            I => \N__24769\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24766\
        );

    \I__5210\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24763\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24778\,
            I => \c0.data_in_field_50\
        );

    \I__5208\ : Odrv12
    port map (
            O => \N__24775\,
            I => \c0.data_in_field_50\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__24772\,
            I => \c0.data_in_field_50\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__24769\,
            I => \c0.data_in_field_50\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__24766\,
            I => \c0.data_in_field_50\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__24763\,
            I => \c0.data_in_field_50\
        );

    \I__5203\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24743\
        );

    \I__5201\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24740\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__24743\,
            I => \N__24737\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__24740\,
            I => \c0.n2053\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__24737\,
            I => \c0.n2053\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__5196\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__24717\,
            I => \c0.n2101\
        );

    \I__5191\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__24708\,
            I => \N__24704\
        );

    \I__5188\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24701\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__24704\,
            I => \N__24696\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24696\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__24696\,
            I => \c0.n2134\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__24693\,
            I => \c0.n31_adj_1900_cascade_\
        );

    \I__5183\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__24687\,
            I => \c0.n35\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__5180\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24677\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__24677\,
            I => \N__24671\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24667\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__24671\,
            I => \N__24664\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24661\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__24667\,
            I => \N__24658\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__24664\,
            I => data_in_0_2
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__24661\,
            I => data_in_0_2
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__24658\,
            I => data_in_0_2
        );

    \I__5170\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__24648\,
            I => \c0.n14\
        );

    \I__5168\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24642\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24642\,
            I => \c0.n5582\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__24639\,
            I => \N__24636\
        );

    \I__5165\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__5163\ : Odrv4
    port map (
            O => \N__24630\,
            I => \c0.n13_adj_1899\
        );

    \I__5162\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24624\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__24624\,
            I => \c0.n17_adj_1902\
        );

    \I__5160\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24615\
        );

    \I__5158\ : Odrv12
    port map (
            O => \N__24615\,
            I => \c0.n25_adj_1907\
        );

    \I__5157\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24609\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__24609\,
            I => \c0.n4_adj_1920\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24600\
        );

    \I__5154\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24597\
        );

    \I__5153\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24594\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24591\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__24600\,
            I => \N__24588\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__24597\,
            I => \N__24585\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24594\,
            I => \N__24582\
        );

    \I__5148\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24578\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__24588\,
            I => \N__24575\
        );

    \I__5146\ : Span12Mux_v
    port map (
            O => \N__24585\,
            I => \N__24572\
        );

    \I__5145\ : Span4Mux_h
    port map (
            O => \N__24582\,
            I => \N__24569\
        );

    \I__5144\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24566\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__24578\,
            I => \c0.data_in_field_122\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__24575\,
            I => \c0.data_in_field_122\
        );

    \I__5141\ : Odrv12
    port map (
            O => \N__24572\,
            I => \c0.data_in_field_122\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__24569\,
            I => \c0.data_in_field_122\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__24566\,
            I => \c0.data_in_field_122\
        );

    \I__5138\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__24552\,
            I => \N__24549\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__24546\,
            I => \c0.n5593\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__24543\,
            I => \N__24540\
        );

    \I__5133\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__24537\,
            I => \N__24533\
        );

    \I__5131\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24530\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__24533\,
            I => \N__24522\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24522\
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__24529\,
            I => \N__24518\
        );

    \I__5127\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24515\
        );

    \I__5126\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24512\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__24522\,
            I => \N__24509\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \N__24506\
        );

    \I__5123\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24503\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24500\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__24512\,
            I => \N__24497\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__24509\,
            I => \N__24494\
        );

    \I__5119\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24491\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__24503\,
            I => \c0.data_in_field_62\
        );

    \I__5117\ : Odrv12
    port map (
            O => \N__24500\,
            I => \c0.data_in_field_62\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__24497\,
            I => \c0.data_in_field_62\
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__24494\,
            I => \c0.data_in_field_62\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__24491\,
            I => \c0.data_in_field_62\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__24480\,
            I => \c0.n5593_cascade_\
        );

    \I__5112\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24474\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__24474\,
            I => \c0.n5430\
        );

    \I__5110\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__24468\,
            I => \c0.n33\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__24465\,
            I => \c0.n5430_cascade_\
        );

    \I__5107\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__5105\ : Odrv12
    port map (
            O => \N__24456\,
            I => \c0.n28_adj_1955\
        );

    \I__5104\ : InMux
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__24450\,
            I => \c0.n5384\
        );

    \I__5102\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24441\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__24438\,
            I => \N__24434\
        );

    \I__5098\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24431\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__24434\,
            I => \c0.n5476\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__24431\,
            I => \c0.n5476\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__24426\,
            I => \N__24423\
        );

    \I__5094\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__24420\,
            I => \N__24417\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__24417\,
            I => \N__24414\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__24414\,
            I => \c0.n5427\
        );

    \I__5090\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__24402\,
            I => \N__24398\
        );

    \I__5086\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24395\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__24398\,
            I => \c0.n5521\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__24395\,
            I => \c0.n5521\
        );

    \I__5083\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__24387\,
            I => \c0.n24_adj_1885\
        );

    \I__5081\ : InMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__24381\,
            I => \N__24377\
        );

    \I__5079\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__24377\,
            I => \N__24369\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24369\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__24369\,
            I => \c0.n1866\
        );

    \I__5075\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24362\
        );

    \I__5074\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24359\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24352\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__24356\,
            I => \N__24349\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__24355\,
            I => \N__24346\
        );

    \I__5069\ : Span4Mux_v
    port map (
            O => \N__24352\,
            I => \N__24339\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__24349\,
            I => \N__24339\
        );

    \I__5067\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24336\
        );

    \I__5066\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24331\
        );

    \I__5065\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24331\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__24339\,
            I => \c0.data_in_field_113\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__24336\,
            I => \c0.data_in_field_113\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__24331\,
            I => \c0.data_in_field_113\
        );

    \I__5061\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__24318\,
            I => \N__24313\
        );

    \I__5058\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24310\
        );

    \I__5057\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24306\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__24313\,
            I => \N__24303\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__24310\,
            I => \N__24300\
        );

    \I__5054\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24296\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__24306\,
            I => \N__24293\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__24303\,
            I => \N__24290\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__24300\,
            I => \N__24287\
        );

    \I__5050\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24284\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__24296\,
            I => \c0.data_in_field_57\
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__24293\,
            I => \c0.data_in_field_57\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__24290\,
            I => \c0.data_in_field_57\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__24287\,
            I => \c0.data_in_field_57\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__24284\,
            I => \c0.data_in_field_57\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__24273\,
            I => \c0.n10_cascade_\
        );

    \I__5043\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24267\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24264\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__24264\,
            I => \N__24260\
        );

    \I__5040\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24257\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__24260\,
            I => \N__24254\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__24254\,
            I => \c0.n5466\
        );

    \I__5036\ : Odrv12
    port map (
            O => \N__24251\,
            I => \c0.n5466\
        );

    \I__5035\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__24243\,
            I => \c0.n5519\
        );

    \I__5033\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24236\
        );

    \I__5032\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24233\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24230\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24227\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__24230\,
            I => \N__24223\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24220\
        );

    \I__5027\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24217\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__24223\,
            I => data_in_7_6
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__24220\,
            I => data_in_7_6
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__24217\,
            I => data_in_7_6
        );

    \I__5023\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24206\
        );

    \I__5022\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24203\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__24206\,
            I => \N__24199\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__24203\,
            I => \N__24196\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24193\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__24199\,
            I => \N__24190\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__24196\,
            I => \N__24187\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__24193\,
            I => data_in_6_6
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__24190\,
            I => data_in_6_6
        );

    \I__5014\ : Odrv4
    port map (
            O => \N__24187\,
            I => data_in_6_6
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__24180\,
            I => \N__24177\
        );

    \I__5012\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24173\
        );

    \I__5011\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24170\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24165\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24162\
        );

    \I__5008\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24159\
        );

    \I__5007\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24156\
        );

    \I__5006\ : Span12Mux_v
    port map (
            O => \N__24165\,
            I => \N__24153\
        );

    \I__5005\ : Odrv12
    port map (
            O => \N__24162\,
            I => data_in_18_0
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__24159\,
            I => data_in_18_0
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__24156\,
            I => data_in_18_0
        );

    \I__5002\ : Odrv12
    port map (
            O => \N__24153\,
            I => data_in_18_0
        );

    \I__5001\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__4999\ : Odrv12
    port map (
            O => \N__24138\,
            I => \c0.n5548\
        );

    \I__4998\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24131\
        );

    \I__4997\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24128\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__24131\,
            I => \N__24123\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24123\
        );

    \I__4994\ : Odrv12
    port map (
            O => \N__24123\,
            I => \c0.n5497\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__24120\,
            I => \N__24116\
        );

    \I__4992\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24113\
        );

    \I__4991\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24110\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__24113\,
            I => \N__24107\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24104\
        );

    \I__4988\ : Odrv12
    port map (
            O => \N__24107\,
            I => \c0.n5515\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__24104\,
            I => \c0.n5515\
        );

    \I__4986\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24093\
        );

    \I__4985\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24086\
        );

    \I__4984\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24086\
        );

    \I__4983\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24086\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__24093\,
            I => \r_Clock_Count_6\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__24086\,
            I => \r_Clock_Count_6\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__4979\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__24072\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__24072\,
            I => n317
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__24069\,
            I => \N__24063\
        );

    \I__4975\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24060\
        );

    \I__4974\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24055\
        );

    \I__4973\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24055\
        );

    \I__4972\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24052\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__24060\,
            I => \r_Clock_Count_4\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__24055\,
            I => \r_Clock_Count_4\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__24052\,
            I => \r_Clock_Count_4\
        );

    \I__4968\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__24042\,
            I => \c0.tx.n10_adj_1868\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__24039\,
            I => \N__24034\
        );

    \I__4965\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24030\
        );

    \I__4964\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24027\
        );

    \I__4963\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24024\
        );

    \I__4962\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24021\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__24030\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24027\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__24024\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__24021\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__4957\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24009\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__24009\,
            I => \c0.tx.n5627\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__24006\,
            I => \n11_adj_1979_cascade_\
        );

    \I__4954\ : InMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__24000\,
            I => \c0.tx.n5629\
        );

    \I__4952\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23993\
        );

    \I__4951\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23990\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__23993\,
            I => \c0.tx.n3120\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__23990\,
            I => \c0.tx.n3120\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \N__23981\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__23984\,
            I => \N__23974\
        );

    \I__4946\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23971\
        );

    \I__4945\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23968\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23963\
        );

    \I__4943\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23963\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23960\
        );

    \I__4941\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23957\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__23971\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__23968\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__23963\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__23960\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__23957\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__23946\,
            I => \c0.tx.n3120_cascade_\
        );

    \I__4934\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23940\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23937\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__23937\,
            I => n313
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__23934\,
            I => \n782_cascade_\
        );

    \I__4930\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23925\
        );

    \I__4929\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23922\
        );

    \I__4928\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23917\
        );

    \I__4927\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23917\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__23925\,
            I => \r_Clock_Count_8\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__23922\,
            I => \r_Clock_Count_8\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__23917\,
            I => \r_Clock_Count_8\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__4922\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23904\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23901\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__23901\,
            I => \N__23898\
        );

    \I__4919\ : Span4Mux_v
    port map (
            O => \N__23898\,
            I => \N__23894\
        );

    \I__4918\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23891\
        );

    \I__4917\ : Sp12to4
    port map (
            O => \N__23894\,
            I => \N__23885\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23885\
        );

    \I__4915\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23882\
        );

    \I__4914\ : Odrv12
    port map (
            O => \N__23885\,
            I => data_in_9_2
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__23882\,
            I => data_in_9_2
        );

    \I__4912\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__23874\,
            I => \c0.n5827\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__4909\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__23865\,
            I => \c0.n1253\
        );

    \I__4907\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__23850\,
            I => \tx_data_7_N_keep\
        );

    \I__4902\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23843\
        );

    \I__4901\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23840\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__23843\,
            I => data_out_18_0
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__23840\,
            I => data_out_18_0
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__23835\,
            I => \N__23832\
        );

    \I__4897\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23828\
        );

    \I__4896\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23825\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__23825\,
            I => data_out_19_0
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__23822\,
            I => data_out_19_0
        );

    \I__4892\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23814\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__23814\,
            I => \c0.n1198\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__23811\,
            I => \c0.n5810_cascade_\
        );

    \I__4889\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23804\
        );

    \I__4888\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23801\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__23804\,
            I => \c0.tx_data_0_N\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__23801\,
            I => \c0.tx_data_0_N\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__23796\,
            I => \c0.tx.n14_adj_1869_cascade_\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__23793\,
            I => \c0.tx.r_SM_Main_2_N_1767_1_cascade_\
        );

    \I__4883\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23787\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__23784\,
            I => \c0.tx.n5821\
        );

    \I__4880\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23775\
        );

    \I__4879\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23768\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23768\
        );

    \I__4877\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23768\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__23775\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__23768\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__23763\,
            I => \N__23760\
        );

    \I__4873\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23757\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__23754\,
            I => n315
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \c0.n17_adj_1913_cascade_\
        );

    \I__4869\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__23745\,
            I => \c0.tx.n5883\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__23742\,
            I => \c0.n1253_cascade_\
        );

    \I__4866\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23733\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__23733\,
            I => \c0.n5830\
        );

    \I__4863\ : CascadeMux
    port map (
            O => \N__23730\,
            I => \c0.n22_adj_1914_cascade_\
        );

    \I__4862\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__23724\,
            I => \tx_data_6_N_keep\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__23721\,
            I => \n5646_cascade_\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__23715\,
            I => n5645
        );

    \I__4857\ : IoInMux
    port map (
            O => \N__23712\,
            I => \N__23709\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__4855\ : Span4Mux_s0_v
    port map (
            O => \N__23706\,
            I => \N__23703\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__23703\,
            I => \N__23700\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__23700\,
            I => \N__23697\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__23694\,
            I => \LED_c\
        );

    \I__4850\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__23685\,
            I => \N__23681\
        );

    \I__4847\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23678\
        );

    \I__4846\ : Span4Mux_h
    port map (
            O => \N__23681\,
            I => \N__23672\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23669\
        );

    \I__4844\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23662\
        );

    \I__4843\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23662\
        );

    \I__4842\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23662\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__23672\,
            I => \c0.data_in_field_110\
        );

    \I__4840\ : Odrv12
    port map (
            O => \N__23669\,
            I => \c0.data_in_field_110\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__23662\,
            I => \c0.data_in_field_110\
        );

    \I__4838\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23651\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23648\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23643\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__23648\,
            I => \N__23643\
        );

    \I__4834\ : Span4Mux_v
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__23640\,
            I => \c0.n5533\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__4831\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23630\
        );

    \I__4830\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23627\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__23630\,
            I => data_out_18_6
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__23627\,
            I => data_out_18_6
        );

    \I__4827\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__23619\,
            I => \N__23616\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__23613\,
            I => \c0.n2077\
        );

    \I__4823\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23607\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__23607\,
            I => \N__23604\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__23601\,
            I => \c0.n5707\
        );

    \I__4819\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23595\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23592\
        );

    \I__4817\ : Odrv12
    port map (
            O => \N__23592\,
            I => \c0.n5710\
        );

    \I__4816\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23586\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__4814\ : Span4Mux_h
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__4813\ : Span4Mux_h
    port map (
            O => \N__23580\,
            I => \N__23577\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__23577\,
            I => \c0.n6198\
        );

    \I__4811\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23570\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23567\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__23570\,
            I => \c0.delay_counter_9\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__23567\,
            I => \c0.delay_counter_9\
        );

    \I__4807\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23558\
        );

    \I__4806\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__23558\,
            I => \c0.delay_counter_2\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__23555\,
            I => \c0.delay_counter_2\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__23550\,
            I => \N__23546\
        );

    \I__4802\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23543\
        );

    \I__4801\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23540\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__23543\,
            I => \c0.delay_counter_0\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__23540\,
            I => \c0.delay_counter_0\
        );

    \I__4798\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23531\
        );

    \I__4797\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__23531\,
            I => \c0.delay_counter_7\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__23528\,
            I => \c0.delay_counter_7\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__4793\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__23514\,
            I => \N__23511\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__23511\,
            I => \N__23506\
        );

    \I__4789\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23501\
        );

    \I__4788\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23501\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__23506\,
            I => data_in_5_0
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__23501\,
            I => data_in_5_0
        );

    \I__4785\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23489\
        );

    \I__4783\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23486\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__23489\,
            I => \N__23483\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23480\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__23483\,
            I => \N__23477\
        );

    \I__4779\ : Span4Mux_h
    port map (
            O => \N__23480\,
            I => \N__23474\
        );

    \I__4778\ : Sp12to4
    port map (
            O => \N__23477\,
            I => \N__23470\
        );

    \I__4777\ : Span4Mux_v
    port map (
            O => \N__23474\,
            I => \N__23467\
        );

    \I__4776\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23464\
        );

    \I__4775\ : Odrv12
    port map (
            O => \N__23470\,
            I => data_in_4_0
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__23467\,
            I => data_in_4_0
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__23464\,
            I => data_in_4_0
        );

    \I__4772\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23453\
        );

    \I__4771\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23446\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23443\
        );

    \I__4768\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23440\
        );

    \I__4767\ : Span4Mux_h
    port map (
            O => \N__23446\,
            I => \N__23437\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__23443\,
            I => \N__23434\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__23440\,
            I => data_in_8_4
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__23437\,
            I => data_in_8_4
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__23434\,
            I => data_in_8_4
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__4761\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__23415\,
            I => \N__23410\
        );

    \I__4757\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23405\
        );

    \I__4756\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23405\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__23410\,
            I => data_in_7_4
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__23405\,
            I => data_in_7_4
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__23400\,
            I => \N__23397\
        );

    \I__4752\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23393\
        );

    \I__4751\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23390\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23387\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23384\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__23387\,
            I => \N__23380\
        );

    \I__4747\ : Span12Mux_v
    port map (
            O => \N__23384\,
            I => \N__23377\
        );

    \I__4746\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23374\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__23380\,
            I => data_in_6_4
        );

    \I__4744\ : Odrv12
    port map (
            O => \N__23377\,
            I => data_in_6_4
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__23374\,
            I => data_in_6_4
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__4741\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23361\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__23361\,
            I => \N__23358\
        );

    \I__4739\ : Span4Mux_v
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__23355\,
            I => \N__23350\
        );

    \I__4737\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23345\
        );

    \I__4736\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23345\
        );

    \I__4735\ : Odrv4
    port map (
            O => \N__23350\,
            I => data_in_5_6
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__23345\,
            I => data_in_5_6
        );

    \I__4733\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23335\
        );

    \I__4732\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23332\
        );

    \I__4731\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23328\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__23335\,
            I => \N__23325\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23322\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23319\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__23328\,
            I => \c0.data_in_field_89\
        );

    \I__4726\ : Odrv12
    port map (
            O => \N__23325\,
            I => \c0.data_in_field_89\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__23322\,
            I => \c0.data_in_field_89\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__23319\,
            I => \c0.data_in_field_89\
        );

    \I__4723\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__23307\,
            I => \N__23303\
        );

    \I__4721\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23300\
        );

    \I__4720\ : Span12Mux_s9_h
    port map (
            O => \N__23303\,
            I => \N__23294\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23291\
        );

    \I__4718\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23284\
        );

    \I__4717\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23284\
        );

    \I__4716\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23284\
        );

    \I__4715\ : Odrv12
    port map (
            O => \N__23294\,
            I => \c0.data_in_field_90\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__23291\,
            I => \c0.data_in_field_90\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__23284\,
            I => \c0.data_in_field_90\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__4711\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__23268\,
            I => \N__23264\
        );

    \I__4708\ : InMux
    port map (
            O => \N__23267\,
            I => \N__23261\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__23264\,
            I => \N__23256\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23256\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__4703\ : Span4Mux_v
    port map (
            O => \N__23250\,
            I => \N__23246\
        );

    \I__4702\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23243\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__23246\,
            I => data_in_7_7
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__23243\,
            I => data_in_7_7
        );

    \I__4699\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23234\
        );

    \I__4698\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23231\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__23234\,
            I => \N__23228\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23222\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__4694\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23218\
        );

    \I__4693\ : Span4Mux_h
    port map (
            O => \N__23222\,
            I => \N__23215\
        );

    \I__4692\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23212\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__23218\,
            I => \c0.data_in_field_37\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__23215\,
            I => \c0.data_in_field_37\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__23212\,
            I => \c0.data_in_field_37\
        );

    \I__4688\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23202\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__23196\,
            I => \N__23192\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__4683\ : Span4Mux_h
    port map (
            O => \N__23192\,
            I => \N__23186\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__23189\,
            I => \c0.data_in_frame_18_0\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__23186\,
            I => \c0.data_in_frame_18_0\
        );

    \I__4680\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23177\
        );

    \I__4679\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23170\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23167\
        );

    \I__4676\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23164\
        );

    \I__4675\ : Odrv12
    port map (
            O => \N__23170\,
            I => data_in_4_1
        );

    \I__4674\ : Odrv4
    port map (
            O => \N__23167\,
            I => data_in_4_1
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__23164\,
            I => data_in_4_1
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__23157\,
            I => \N__23153\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__23156\,
            I => \N__23150\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23146\
        );

    \I__4669\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23143\
        );

    \I__4668\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23140\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__23146\,
            I => \N__23137\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23133\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__23140\,
            I => \N__23130\
        );

    \I__4664\ : Span4Mux_h
    port map (
            O => \N__23137\,
            I => \N__23127\
        );

    \I__4663\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23124\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__23133\,
            I => \N__23121\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__23130\,
            I => \N__23116\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__23127\,
            I => \N__23116\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__23124\,
            I => data_in_18_7
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__23121\,
            I => data_in_18_7
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__23116\,
            I => data_in_18_7
        );

    \I__4656\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23106\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__23106\,
            I => \N__23103\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__23103\,
            I => \N__23099\
        );

    \I__4653\ : InMux
    port map (
            O => \N__23102\,
            I => \N__23096\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__23099\,
            I => \N__23092\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__23096\,
            I => \N__23089\
        );

    \I__4650\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23086\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__23092\,
            I => data_in_17_7
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__23089\,
            I => data_in_17_7
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__23086\,
            I => data_in_17_7
        );

    \I__4646\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23076\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__4644\ : Odrv12
    port map (
            O => \N__23073\,
            I => \c0.n6_adj_1918\
        );

    \I__4643\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23066\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__23069\,
            I => \N__23063\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23059\
        );

    \I__4640\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23056\
        );

    \I__4639\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23053\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__23059\,
            I => \N__23048\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__23048\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__23053\,
            I => \N__23044\
        );

    \I__4635\ : Span4Mux_h
    port map (
            O => \N__23048\,
            I => \N__23041\
        );

    \I__4634\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23038\
        );

    \I__4633\ : Span12Mux_s9_h
    port map (
            O => \N__23044\,
            I => \N__23035\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__23041\,
            I => \N__23032\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__23038\,
            I => data_in_1_4
        );

    \I__4630\ : Odrv12
    port map (
            O => \N__23035\,
            I => data_in_1_4
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__23032\,
            I => data_in_1_4
        );

    \I__4628\ : InMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__23017\
        );

    \I__4626\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23014\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__23020\,
            I => \N__23010\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__23017\,
            I => \N__23007\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__23014\,
            I => \N__23004\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__23013\,
            I => \N__23000\
        );

    \I__4621\ : InMux
    port map (
            O => \N__23010\,
            I => \N__22997\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__23007\,
            I => \N__22994\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__23004\,
            I => \N__22991\
        );

    \I__4618\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22986\
        );

    \I__4617\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22986\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__22997\,
            I => \c0.data_in_field_18\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__22994\,
            I => \c0.data_in_field_18\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__22991\,
            I => \c0.data_in_field_18\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__22986\,
            I => \c0.data_in_field_18\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22974\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__22974\,
            I => \c0.n5372\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__22971\,
            I => \c0.n2043_cascade_\
        );

    \I__4609\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22963\
        );

    \I__4608\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22960\
        );

    \I__4607\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22956\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22953\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22950\
        );

    \I__4604\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22946\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__22956\,
            I => \N__22943\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__22953\,
            I => \N__22940\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__22950\,
            I => \N__22937\
        );

    \I__4600\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22934\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__22946\,
            I => \c0.data_in_field_107\
        );

    \I__4598\ : Odrv12
    port map (
            O => \N__22943\,
            I => \c0.data_in_field_107\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__22940\,
            I => \c0.data_in_field_107\
        );

    \I__4596\ : Odrv4
    port map (
            O => \N__22937\,
            I => \c0.data_in_field_107\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__22934\,
            I => \c0.data_in_field_107\
        );

    \I__4594\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22920\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__22920\,
            I => \N__22917\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__22917\,
            I => \N__22912\
        );

    \I__4591\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22909\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22906\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__22912\,
            I => \N__22903\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__22909\,
            I => data_in_13_6
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__22906\,
            I => data_in_13_6
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__22903\,
            I => data_in_13_6
        );

    \I__4585\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22892\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__22895\,
            I => \N__22889\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__22892\,
            I => \N__22886\
        );

    \I__4582\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22883\
        );

    \I__4581\ : Sp12to4
    port map (
            O => \N__22886\,
            I => \N__22878\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22878\
        );

    \I__4579\ : Span12Mux_s11_v
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__4578\ : Odrv12
    port map (
            O => \N__22875\,
            I => \c0.n5443\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__22863\,
            I => \c0.n47_adj_1897\
        );

    \I__4573\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__22851\,
            I => \c0.n48_adj_1895\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__22848\,
            I => \c0.n5567_cascade_\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__22842\,
            I => \c0.n49\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__4565\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__4563\ : Span4Mux_v
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__22827\,
            I => \c0.n6219\
        );

    \I__4561\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22820\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__22823\,
            I => \N__22817\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22814\
        );

    \I__4558\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22809\
        );

    \I__4557\ : Span4Mux_v
    port map (
            O => \N__22814\,
            I => \N__22806\
        );

    \I__4556\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22801\
        );

    \I__4555\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22801\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__22809\,
            I => \c0.data_in_field_5\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__22806\,
            I => \c0.data_in_field_5\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__22801\,
            I => \c0.data_in_field_5\
        );

    \I__4551\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22790\
        );

    \I__4550\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22787\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__22790\,
            I => \N__22784\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22781\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__22784\,
            I => \N__22778\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__22781\,
            I => \N__22773\
        );

    \I__4545\ : Span4Mux_h
    port map (
            O => \N__22778\,
            I => \N__22773\
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__22773\,
            I => \c0.n1979\
        );

    \I__4543\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__22767\,
            I => \N__22764\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__22764\,
            I => \N__22760\
        );

    \I__4540\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22757\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__22760\,
            I => \N__22752\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__22757\,
            I => \N__22752\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__22752\,
            I => \c0.n1958\
        );

    \I__4536\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__4534\ : Span4Mux_v
    port map (
            O => \N__22743\,
            I => \N__22739\
        );

    \I__4533\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22736\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__22739\,
            I => \N__22731\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__22736\,
            I => \N__22731\
        );

    \I__4530\ : Span4Mux_h
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__22728\,
            I => \c0.n2056\
        );

    \I__4528\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22722\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__22722\,
            I => \c0.n5506\
        );

    \I__4526\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__4524\ : Span4Mux_h
    port map (
            O => \N__22713\,
            I => \N__22709\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22706\
        );

    \I__4522\ : Span4Mux_h
    port map (
            O => \N__22709\,
            I => \N__22701\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__22706\,
            I => \N__22701\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__22701\,
            I => \c0.n5575\
        );

    \I__4519\ : CascadeMux
    port map (
            O => \N__22698\,
            I => \c0.n5506_cascade_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22692\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22688\
        );

    \I__4516\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22685\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__22688\,
            I => \N__22682\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22679\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__22682\,
            I => \c0.n5539\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__22679\,
            I => \c0.n5539\
        );

    \I__4511\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22670\
        );

    \I__4510\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22667\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__22670\,
            I => \N__22664\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22661\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__22664\,
            I => \N__22658\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__22661\,
            I => \N__22655\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__22658\,
            I => \c0.n1779\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__22655\,
            I => \c0.n1779\
        );

    \I__4503\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22646\
        );

    \I__4502\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22643\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22639\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22634\
        );

    \I__4499\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22631\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__22639\,
            I => \N__22628\
        );

    \I__4497\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22625\
        );

    \I__4496\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22622\
        );

    \I__4495\ : Span4Mux_h
    port map (
            O => \N__22634\,
            I => \N__22619\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__22631\,
            I => \c0.data_in_field_60\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__22628\,
            I => \c0.data_in_field_60\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__22625\,
            I => \c0.data_in_field_60\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__22622\,
            I => \c0.data_in_field_60\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__22619\,
            I => \c0.data_in_field_60\
        );

    \I__4489\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22605\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__22605\,
            I => \N__22601\
        );

    \I__4487\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22598\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__22601\,
            I => \c0.n5500\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__22598\,
            I => \c0.n5500\
        );

    \I__4484\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22586\
        );

    \I__4482\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22583\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__22586\,
            I => \N__22579\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22576\
        );

    \I__4479\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22571\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__22579\,
            I => \N__22566\
        );

    \I__4477\ : Span4Mux_h
    port map (
            O => \N__22576\,
            I => \N__22566\
        );

    \I__4476\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22563\
        );

    \I__4475\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22560\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__22571\,
            I => \c0.data_in_field_19\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__22566\,
            I => \c0.data_in_field_19\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__22563\,
            I => \c0.data_in_field_19\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__22560\,
            I => \c0.data_in_field_19\
        );

    \I__4470\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22548\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__4468\ : Span4Mux_s3_h
    port map (
            O => \N__22545\,
            I => \N__22541\
        );

    \I__4467\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22538\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__22541\,
            I => \N__22535\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__22535\,
            I => \N__22526\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__22532\,
            I => \N__22523\
        );

    \I__4462\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22520\
        );

    \I__4461\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22515\
        );

    \I__4460\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22515\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__22526\,
            I => \c0.data_in_field_139\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__22523\,
            I => \c0.data_in_field_139\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__22520\,
            I => \c0.data_in_field_139\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__22515\,
            I => \c0.data_in_field_139\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__4454\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22498\
        );

    \I__4453\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22495\
        );

    \I__4452\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22492\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__22498\,
            I => data_in_5_5
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__22495\,
            I => data_in_5_5
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__22492\,
            I => data_in_5_5
        );

    \I__4448\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22481\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__22484\,
            I => \N__22478\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22475\
        );

    \I__4445\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22472\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__22475\,
            I => \N__22469\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22464\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__22469\,
            I => \N__22464\
        );

    \I__4441\ : Span4Mux_h
    port map (
            O => \N__22464\,
            I => \N__22460\
        );

    \I__4440\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22457\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__22460\,
            I => data_in_6_1
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__22457\,
            I => data_in_6_1
        );

    \I__4437\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22446\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__22440\,
            I => \N__22435\
        );

    \I__4432\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22430\
        );

    \I__4431\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22430\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__22435\,
            I => data_in_5_1
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__22430\,
            I => data_in_5_1
        );

    \I__4428\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__4425\ : Sp12to4
    port map (
            O => \N__22416\,
            I => \N__22411\
        );

    \I__4424\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22406\
        );

    \I__4423\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22406\
        );

    \I__4422\ : Odrv12
    port map (
            O => \N__22411\,
            I => data_in_16_7
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__22406\,
            I => data_in_16_7
        );

    \I__4420\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22398\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__22398\,
            I => \c0.n25\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__4417\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__4415\ : Span4Mux_h
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__22383\,
            I => \c0.n23\
        );

    \I__4413\ : InMux
    port map (
            O => \N__22380\,
            I => \N__22377\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__22377\,
            I => \N__22374\
        );

    \I__4411\ : Sp12to4
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__4410\ : Span12Mux_v
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__4409\ : Odrv12
    port map (
            O => \N__22368\,
            I => \c0.n22_adj_1890\
        );

    \I__4408\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22360\
        );

    \I__4407\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22357\
        );

    \I__4406\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22354\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__22360\,
            I => \N__22351\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22347\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__22354\,
            I => \N__22342\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__22351\,
            I => \N__22339\
        );

    \I__4401\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22336\
        );

    \I__4400\ : Span4Mux_h
    port map (
            O => \N__22347\,
            I => \N__22333\
        );

    \I__4399\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22328\
        );

    \I__4398\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22328\
        );

    \I__4397\ : Odrv12
    port map (
            O => \N__22342\,
            I => \c0.data_in_field_61\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__22339\,
            I => \c0.data_in_field_61\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__22336\,
            I => \c0.data_in_field_61\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__22333\,
            I => \c0.data_in_field_61\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__22328\,
            I => \c0.data_in_field_61\
        );

    \I__4392\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22313\
        );

    \I__4391\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22310\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22304\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22304\
        );

    \I__4388\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22301\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__22304\,
            I => \N__22297\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__22301\,
            I => \N__22294\
        );

    \I__4385\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22291\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__22297\,
            I => \N__22288\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__22294\,
            I => \N__22285\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__22291\,
            I => data_in_3_1
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__22288\,
            I => data_in_3_1
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__22285\,
            I => data_in_3_1
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__22278\,
            I => \N__22275\
        );

    \I__4378\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22271\
        );

    \I__4377\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22268\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22265\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__22268\,
            I => \N__22261\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__22265\,
            I => \N__22258\
        );

    \I__4373\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22255\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__22261\,
            I => \N__22252\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__22258\,
            I => \N__22249\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__22255\,
            I => data_in_0_0
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__22252\,
            I => data_in_0_0
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__22249\,
            I => data_in_0_0
        );

    \I__4367\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__4365\ : Span4Mux_s3_h
    port map (
            O => \N__22236\,
            I => \N__22232\
        );

    \I__4364\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22229\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__22232\,
            I => \N__22223\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22223\
        );

    \I__4361\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22219\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__22223\,
            I => \N__22216\
        );

    \I__4359\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22213\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__22219\,
            I => \c0.data_in_field_0\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__22216\,
            I => \c0.data_in_field_0\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__22213\,
            I => \c0.data_in_field_0\
        );

    \I__4355\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22199\
        );

    \I__4353\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22196\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__22199\,
            I => \N__22189\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__22196\,
            I => \N__22189\
        );

    \I__4350\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22183\
        );

    \I__4349\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22183\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__22189\,
            I => \N__22180\
        );

    \I__4347\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22177\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__22183\,
            I => \c0.data_in_field_117\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__22180\,
            I => \c0.data_in_field_117\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__22177\,
            I => \c0.data_in_field_117\
        );

    \I__4343\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__22167\,
            I => \N__22163\
        );

    \I__4341\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22160\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__22163\,
            I => \c0.n1855\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__22160\,
            I => \c0.n1855\
        );

    \I__4338\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__4336\ : Span12Mux_v
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__4335\ : Odrv12
    port map (
            O => \N__22146\,
            I => \c0.n13\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__22143\,
            I => \c0.n12_adj_1898_cascade_\
        );

    \I__4333\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__22137\,
            I => \c0.tx.n5885\
        );

    \I__4331\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22130\
        );

    \I__4330\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22127\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__22130\,
            I => \c0.tx.n15\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__22127\,
            I => \c0.tx.n15\
        );

    \I__4327\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__22119\,
            I => \c0.tx.n5884\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22112\
        );

    \I__4324\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22109\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__22112\,
            I => \N__22105\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22102\
        );

    \I__4321\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22099\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__22105\,
            I => data_in_4_3
        );

    \I__4319\ : Odrv12
    port map (
            O => \N__22102\,
            I => data_in_4_3
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__22099\,
            I => data_in_4_3
        );

    \I__4317\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22088\
        );

    \I__4316\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22084\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__22088\,
            I => \N__22081\
        );

    \I__4314\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22078\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__22084\,
            I => \N__22074\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__22081\,
            I => \N__22069\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22069\
        );

    \I__4310\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22066\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__22074\,
            I => \N__22063\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__22069\,
            I => data_in_3_3
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__22066\,
            I => data_in_3_3
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__22063\,
            I => data_in_3_3
        );

    \I__4305\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22051\
        );

    \I__4304\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22048\
        );

    \I__4303\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22045\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__22051\,
            I => \N__22041\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__22048\,
            I => \N__22038\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__22045\,
            I => \N__22035\
        );

    \I__4299\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22032\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__22041\,
            I => \N__22027\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__22038\,
            I => \N__22027\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__22035\,
            I => data_in_2_2
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__22032\,
            I => data_in_2_2
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__22027\,
            I => data_in_2_2
        );

    \I__4293\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22016\
        );

    \I__4292\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22013\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22010\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__22007\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__22002\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__22007\,
            I => \N__21999\
        );

    \I__4287\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21996\
        );

    \I__4286\ : InMux
    port map (
            O => \N__22005\,
            I => \N__21993\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__22002\,
            I => data_in_1_2
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__21999\,
            I => data_in_1_2
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__21996\,
            I => data_in_1_2
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__21993\,
            I => data_in_1_2
        );

    \I__4281\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21979\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21976\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__21982\,
            I => \N__21971\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__21979\,
            I => \N__21968\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__21976\,
            I => \N__21965\
        );

    \I__4276\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21962\
        );

    \I__4275\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21959\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21956\
        );

    \I__4273\ : Span12Mux_s5_h
    port map (
            O => \N__21968\,
            I => \N__21953\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__21965\,
            I => \N__21950\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__21962\,
            I => \N__21945\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21945\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__21956\,
            I => \c0.data_in_field_80\
        );

    \I__4268\ : Odrv12
    port map (
            O => \N__21953\,
            I => \c0.data_in_field_80\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__21950\,
            I => \c0.data_in_field_80\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__21945\,
            I => \c0.data_in_field_80\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__21936\,
            I => \c0.n42_cascade_\
        );

    \I__4264\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21930\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__21918\,
            I => \c0.n48\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__21915\,
            I => \N__21911\
        );

    \I__4257\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21907\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21904\
        );

    \I__4255\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21901\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__21907\,
            I => \N__21896\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21896\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21892\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__21896\,
            I => \N__21889\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21886\
        );

    \I__4249\ : Span4Mux_h
    port map (
            O => \N__21892\,
            I => \N__21881\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__21889\,
            I => \N__21881\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__21886\,
            I => data_in_19_0
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__21881\,
            I => data_in_19_0
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__4244\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21869\
        );

    \I__4243\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21866\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21863\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21860\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__21863\,
            I => \N__21857\
        );

    \I__4239\ : Span4Mux_s3_h
    port map (
            O => \N__21860\,
            I => \N__21854\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__21857\,
            I => \N__21848\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__21854\,
            I => \N__21848\
        );

    \I__4236\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21845\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__21848\,
            I => data_in_15_7
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__21845\,
            I => data_in_15_7
        );

    \I__4233\ : InMux
    port map (
            O => \N__21840\,
            I => \bfn_9_27_0_\
        );

    \I__4232\ : InMux
    port map (
            O => \N__21837\,
            I => \c0.tx.n4764\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21834\,
            I => \c0.tx.n4765\
        );

    \I__4230\ : InMux
    port map (
            O => \N__21831\,
            I => \c0.tx.n4766\
        );

    \I__4229\ : InMux
    port map (
            O => \N__21828\,
            I => \c0.tx.n4767\
        );

    \I__4228\ : InMux
    port map (
            O => \N__21825\,
            I => \c0.tx.n4768\
        );

    \I__4227\ : InMux
    port map (
            O => \N__21822\,
            I => \c0.tx.n4769\
        );

    \I__4226\ : InMux
    port map (
            O => \N__21819\,
            I => \c0.tx.n4770\
        );

    \I__4225\ : InMux
    port map (
            O => \N__21816\,
            I => \bfn_9_28_0_\
        );

    \I__4224\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21805\
        );

    \I__4222\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21802\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21799\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__21805\,
            I => \N__21790\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__21802\,
            I => \N__21790\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21799\,
            I => \N__21790\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__21798\,
            I => \N__21787\
        );

    \I__4216\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21784\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__21790\,
            I => \N__21781\
        );

    \I__4214\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21778\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__21784\,
            I => \c0.data_in_field_4\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__21781\,
            I => \c0.data_in_field_4\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__21778\,
            I => \c0.data_in_field_4\
        );

    \I__4210\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21766\
        );

    \I__4209\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21762\
        );

    \I__4208\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21759\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21756\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__21765\,
            I => \N__21753\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21750\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__21759\,
            I => \N__21747\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__21756\,
            I => \N__21744\
        );

    \I__4202\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21740\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__21750\,
            I => \N__21737\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__21747\,
            I => \N__21734\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__21744\,
            I => \N__21731\
        );

    \I__4198\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21728\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__21740\,
            I => \c0.data_in_field_12\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__21737\,
            I => \c0.data_in_field_12\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__21734\,
            I => \c0.data_in_field_12\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__21731\,
            I => \c0.data_in_field_12\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__21728\,
            I => \c0.data_in_field_12\
        );

    \I__4192\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21714\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N__21711\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__21711\,
            I => \N__21708\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__21708\,
            I => \N__21705\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__21705\,
            I => \c0.n5722\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__21702\,
            I => \c0.tx.n3631_cascade_\
        );

    \I__4186\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21694\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__21698\,
            I => \N__21690\
        );

    \I__4184\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21687\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__21694\,
            I => \N__21684\
        );

    \I__4182\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21681\
        );

    \I__4181\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21677\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21674\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__21684\,
            I => \N__21669\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__21681\,
            I => \N__21669\
        );

    \I__4177\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21666\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__21677\,
            I => \c0.data_in_field_20\
        );

    \I__4175\ : Odrv12
    port map (
            O => \N__21674\,
            I => \c0.data_in_field_20\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__21669\,
            I => \c0.data_in_field_20\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__21666\,
            I => \c0.data_in_field_20\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__4171\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21651\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__21651\,
            I => \c0.n6189\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__21648\,
            I => \c0.tx.n5812_cascade_\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__21645\,
            I => \c0.tx.n14_cascade_\
        );

    \I__4167\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21639\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21635\
        );

    \I__4165\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21632\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__21635\,
            I => \N__21629\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21632\,
            I => \r_Tx_Data_7\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__21629\,
            I => \r_Tx_Data_7\
        );

    \I__4161\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21620\
        );

    \I__4160\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21617\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__21620\,
            I => \r_Tx_Data_6\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__21617\,
            I => \r_Tx_Data_6\
        );

    \I__4157\ : InMux
    port map (
            O => \N__21612\,
            I => \c0.n4759\
        );

    \I__4156\ : InMux
    port map (
            O => \N__21609\,
            I => \c0.n4760\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21606\,
            I => \bfn_9_24_0_\
        );

    \I__4154\ : InMux
    port map (
            O => \N__21603\,
            I => \c0.n4762\
        );

    \I__4153\ : InMux
    port map (
            O => \N__21600\,
            I => \c0.n4763\
        );

    \I__4152\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21593\
        );

    \I__4151\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21590\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__21593\,
            I => \c0.delay_counter_1\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__21590\,
            I => \c0.delay_counter_1\
        );

    \I__4148\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21581\
        );

    \I__4147\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21578\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__21581\,
            I => \c0.delay_counter_5\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__21578\,
            I => \c0.delay_counter_5\
        );

    \I__4144\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21569\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__21572\,
            I => \N__21565\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21562\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__21568\,
            I => \N__21559\
        );

    \I__4140\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21556\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__4138\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21550\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__21556\,
            I => \c0.data_in_field_116\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__21553\,
            I => \c0.data_in_field_116\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__21550\,
            I => \c0.data_in_field_116\
        );

    \I__4134\ : InMux
    port map (
            O => \N__21543\,
            I => \N__21540\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__21540\,
            I => \N__21534\
        );

    \I__4132\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21529\
        );

    \I__4131\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21529\
        );

    \I__4130\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21524\
        );

    \I__4129\ : Span4Mux_h
    port map (
            O => \N__21534\,
            I => \N__21521\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21518\
        );

    \I__4127\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21513\
        );

    \I__4126\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21513\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__21524\,
            I => \c0.data_in_field_124\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__21521\,
            I => \c0.data_in_field_124\
        );

    \I__4123\ : Odrv12
    port map (
            O => \N__21518\,
            I => \c0.data_in_field_124\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__21513\,
            I => \c0.data_in_field_124\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__21504\,
            I => \c0.n6171_cascade_\
        );

    \I__4120\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21498\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__21495\,
            I => \N__21492\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__21492\,
            I => \N__21489\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__21489\,
            I => \c0.n5731\
        );

    \I__4115\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21482\
        );

    \I__4114\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21479\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__21482\,
            I => \N__21475\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21472\
        );

    \I__4111\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21468\
        );

    \I__4110\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21465\
        );

    \I__4109\ : Span4Mux_v
    port map (
            O => \N__21472\,
            I => \N__21462\
        );

    \I__4108\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21459\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21456\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__21465\,
            I => data_in_3_2
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__21462\,
            I => data_in_3_2
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__21459\,
            I => data_in_3_2
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__21456\,
            I => data_in_3_2
        );

    \I__4102\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21444\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__4100\ : Span4Mux_h
    port map (
            O => \N__21441\,
            I => \N__21437\
        );

    \I__4099\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21434\
        );

    \I__4098\ : Span4Mux_h
    port map (
            O => \N__21437\,
            I => \N__21431\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21428\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__21431\,
            I => \c0.n1955\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__21428\,
            I => \c0.n1955\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__21423\,
            I => \N__21420\
        );

    \I__4093\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21414\
        );

    \I__4091\ : Span4Mux_v
    port map (
            O => \N__21414\,
            I => \N__21409\
        );

    \I__4090\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21404\
        );

    \I__4089\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21404\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__21409\,
            I => data_in_4_2
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__21404\,
            I => data_in_4_2
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__21399\,
            I => \N__21396\
        );

    \I__4085\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21392\
        );

    \I__4084\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21388\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21385\
        );

    \I__4082\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21382\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__21388\,
            I => \N__21378\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__21385\,
            I => \N__21375\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21372\
        );

    \I__4078\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21369\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__21378\,
            I => \N__21366\
        );

    \I__4076\ : Sp12to4
    port map (
            O => \N__21375\,
            I => \N__21361\
        );

    \I__4075\ : Span12Mux_v
    port map (
            O => \N__21372\,
            I => \N__21361\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__21369\,
            I => data_in_18_5
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__21366\,
            I => data_in_18_5
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__21361\,
            I => data_in_18_5
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__21354\,
            I => \N__21351\
        );

    \I__4070\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21344\
        );

    \I__4068\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21341\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__21344\,
            I => \N__21337\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21334\
        );

    \I__4065\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21331\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__21337\,
            I => data_in_17_5
        );

    \I__4063\ : Odrv12
    port map (
            O => \N__21334\,
            I => data_in_17_5
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__21331\,
            I => data_in_17_5
        );

    \I__4061\ : InMux
    port map (
            O => \N__21324\,
            I => \c0.n4754\
        );

    \I__4060\ : InMux
    port map (
            O => \N__21321\,
            I => \c0.n4755\
        );

    \I__4059\ : InMux
    port map (
            O => \N__21318\,
            I => \c0.n4756\
        );

    \I__4058\ : InMux
    port map (
            O => \N__21315\,
            I => \c0.n4757\
        );

    \I__4057\ : InMux
    port map (
            O => \N__21312\,
            I => \c0.n4758\
        );

    \I__4056\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21305\
        );

    \I__4055\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21302\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21299\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__21302\,
            I => \N__21296\
        );

    \I__4052\ : Span4Mux_v
    port map (
            O => \N__21299\,
            I => \N__21293\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__21296\,
            I => \N__21290\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__21293\,
            I => \N__21286\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__21290\,
            I => \N__21283\
        );

    \I__4048\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21280\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__21286\,
            I => data_in_15_5
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__21283\,
            I => data_in_15_5
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__21280\,
            I => data_in_15_5
        );

    \I__4044\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21270\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__21270\,
            I => \c0.n6414\
        );

    \I__4042\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21261\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__21261\,
            I => \c0.n5563\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__4038\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__21249\,
            I => \N__21245\
        );

    \I__4035\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21242\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__21245\,
            I => \N__21236\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__21242\,
            I => \N__21236\
        );

    \I__4032\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21233\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__21236\,
            I => data_in_11_1
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__21233\,
            I => data_in_11_1
        );

    \I__4029\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21224\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__21227\,
            I => \N__21221\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21218\
        );

    \I__4026\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21215\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__21218\,
            I => \N__21212\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21206\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__21212\,
            I => \N__21203\
        );

    \I__4022\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21200\
        );

    \I__4021\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21195\
        );

    \I__4020\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21195\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__21206\,
            I => \N__21192\
        );

    \I__4018\ : Odrv4
    port map (
            O => \N__21203\,
            I => \c0.data_in_field_45\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__21200\,
            I => \c0.data_in_field_45\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__21195\,
            I => \c0.data_in_field_45\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__21192\,
            I => \c0.data_in_field_45\
        );

    \I__4014\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__21180\,
            I => \N__21175\
        );

    \I__4012\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21172\
        );

    \I__4011\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21169\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__21175\,
            I => \N__21164\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21164\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21161\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__21164\,
            I => \c0.n2065\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__21161\,
            I => \c0.n2065\
        );

    \I__4005\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21153\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__21153\,
            I => \c0.n18\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__21150\,
            I => \c0.n2149_cascade_\
        );

    \I__4002\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__4000\ : Span12Mux_v
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__3999\ : Odrv12
    port map (
            O => \N__21138\,
            I => \c0.n21\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__3997\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__21129\,
            I => \N__21124\
        );

    \I__3995\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21121\
        );

    \I__3994\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21118\
        );

    \I__3993\ : Odrv12
    port map (
            O => \N__21124\,
            I => data_in_17_3
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__21121\,
            I => data_in_17_3
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__21118\,
            I => data_in_17_3
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__21111\,
            I => \N__21108\
        );

    \I__3989\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__21102\,
            I => \N__21096\
        );

    \I__3986\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21093\
        );

    \I__3985\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21088\
        );

    \I__3984\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21088\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__21096\,
            I => data_in_2_3
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__21093\,
            I => data_in_2_3
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__21088\,
            I => data_in_2_3
        );

    \I__3980\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21077\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__21080\,
            I => \N__21074\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21071\
        );

    \I__3977\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21067\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__21071\,
            I => \N__21064\
        );

    \I__3975\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21061\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__21067\,
            I => \N__21056\
        );

    \I__3973\ : Span4Mux_h
    port map (
            O => \N__21064\,
            I => \N__21056\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__21061\,
            I => data_in_6_7
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__21056\,
            I => data_in_6_7
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__3969\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__21045\,
            I => \N__21041\
        );

    \I__3967\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21038\
        );

    \I__3966\ : Span4Mux_v
    port map (
            O => \N__21041\,
            I => \N__21033\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__21038\,
            I => \N__21033\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__21033\,
            I => \N__21029\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__21032\,
            I => \N__21026\
        );

    \I__3962\ : Span4Mux_h
    port map (
            O => \N__21029\,
            I => \N__21023\
        );

    \I__3961\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21020\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__21023\,
            I => data_in_6_5
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__21020\,
            I => data_in_6_5
        );

    \I__3958\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21009\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__21009\,
            I => \N__21006\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__21006\,
            I => \c0.n25_adj_1948\
        );

    \I__3954\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20997\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20994\
        );

    \I__3952\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20991\
        );

    \I__3951\ : InMux
    port map (
            O => \N__21000\,
            I => \N__20988\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__20997\,
            I => \N__20985\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20982\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20979\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__20988\,
            I => \N__20968\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__20985\,
            I => \N__20968\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__20982\,
            I => \N__20968\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__20979\,
            I => \N__20968\
        );

    \I__3943\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20963\
        );

    \I__3942\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20963\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__20968\,
            I => \c0.data_in_field_94\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20963\,
            I => \c0.data_in_field_94\
        );

    \I__3939\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20955\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__20955\,
            I => \N__20952\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__20952\,
            I => \N__20947\
        );

    \I__3936\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20944\
        );

    \I__3935\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20940\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__20947\,
            I => \N__20935\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20935\
        );

    \I__3932\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20932\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__20940\,
            I => \c0.data_in_field_66\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__20935\,
            I => \c0.data_in_field_66\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__20932\,
            I => \c0.data_in_field_66\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__20925\,
            I => \N__20920\
        );

    \I__3927\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20917\
        );

    \I__3926\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20914\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20910\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20907\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20904\
        );

    \I__3922\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20901\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__20910\,
            I => \c0.data_in_field_79\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__20907\,
            I => \c0.data_in_field_79\
        );

    \I__3919\ : Odrv12
    port map (
            O => \N__20904\,
            I => \c0.data_in_field_79\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__20901\,
            I => \c0.data_in_field_79\
        );

    \I__3917\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20888\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20885\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__20885\,
            I => \N__20879\
        );

    \I__3913\ : Odrv12
    port map (
            O => \N__20882\,
            I => \c0.n5545\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__20879\,
            I => \c0.n5545\
        );

    \I__3911\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__3909\ : Span4Mux_h
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__3908\ : Span4Mux_h
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__20862\,
            I => \c0.n46\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__20859\,
            I => \N__20854\
        );

    \I__3905\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20851\
        );

    \I__3904\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20848\
        );

    \I__3903\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20844\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__20851\,
            I => \N__20839\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__20848\,
            I => \N__20836\
        );

    \I__3900\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20833\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__20844\,
            I => \N__20830\
        );

    \I__3898\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20825\
        );

    \I__3897\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20825\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__20839\,
            I => \N__20818\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__20836\,
            I => \N__20818\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20818\
        );

    \I__3893\ : Odrv12
    port map (
            O => \N__20830\,
            I => \c0.data_in_field_95\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__20825\,
            I => \c0.data_in_field_95\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__20818\,
            I => \c0.data_in_field_95\
        );

    \I__3890\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20806\
        );

    \I__3889\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20803\
        );

    \I__3888\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20799\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__20806\,
            I => \N__20796\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20793\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20790\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20787\
        );

    \I__3883\ : Span4Mux_s3_h
    port map (
            O => \N__20796\,
            I => \N__20784\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__20793\,
            I => \N__20781\
        );

    \I__3881\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20777\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__20787\,
            I => \N__20770\
        );

    \I__3879\ : Span4Mux_v
    port map (
            O => \N__20784\,
            I => \N__20770\
        );

    \I__3878\ : Span4Mux_v
    port map (
            O => \N__20781\,
            I => \N__20770\
        );

    \I__3877\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20767\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__20777\,
            I => \c0.data_in_field_96\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__20770\,
            I => \c0.data_in_field_96\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__20767\,
            I => \c0.data_in_field_96\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__20757\,
            I => \c0.n5590\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__20754\,
            I => \c0.n40_cascade_\
        );

    \I__3870\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__20745\,
            I => \c0.n45_adj_1892\
        );

    \I__3867\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20736\
        );

    \I__3866\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20733\
        );

    \I__3865\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20730\
        );

    \I__3864\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20727\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__20736\,
            I => \N__20724\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20721\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20718\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20715\
        );

    \I__3859\ : Span12Mux_v
    port map (
            O => \N__20724\,
            I => \N__20710\
        );

    \I__3858\ : Span12Mux_s8_h
    port map (
            O => \N__20721\,
            I => \N__20707\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__20718\,
            I => \N__20702\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__20715\,
            I => \N__20702\
        );

    \I__3855\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20697\
        );

    \I__3854\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20697\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__20710\,
            I => \c0.data_in_field_132\
        );

    \I__3852\ : Odrv12
    port map (
            O => \N__20707\,
            I => \c0.data_in_field_132\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__20702\,
            I => \c0.data_in_field_132\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__20697\,
            I => \c0.data_in_field_132\
        );

    \I__3849\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__20682\,
            I => \c0.n1969\
        );

    \I__3846\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__20676\,
            I => \N__20672\
        );

    \I__3844\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20669\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__20672\,
            I => \N__20664\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__20669\,
            I => \N__20664\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__20664\,
            I => \c0.n5403\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20654\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20650\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__20654\,
            I => \N__20647\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20643\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20640\
        );

    \I__3834\ : Span4Mux_v
    port map (
            O => \N__20647\,
            I => \N__20637\
        );

    \I__3833\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20634\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20631\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__20640\,
            I => \N__20626\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__20637\,
            I => \N__20626\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__20634\,
            I => data_in_19_4
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__20631\,
            I => data_in_19_4
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__20626\,
            I => data_in_19_4
        );

    \I__3826\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20616\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20610\
        );

    \I__3824\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20607\
        );

    \I__3823\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20604\
        );

    \I__3822\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20601\
        );

    \I__3821\ : Span12Mux_s6_h
    port map (
            O => \N__20610\,
            I => \N__20598\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20593\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20593\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__20601\,
            I => \c0.data_in_field_115\
        );

    \I__3817\ : Odrv12
    port map (
            O => \N__20598\,
            I => \c0.data_in_field_115\
        );

    \I__3816\ : Odrv12
    port map (
            O => \N__20593\,
            I => \c0.data_in_field_115\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__20586\,
            I => \c0.n1855_cascade_\
        );

    \I__3814\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__20577\,
            I => \N__20573\
        );

    \I__3811\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20570\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__20573\,
            I => \N__20567\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__20570\,
            I => \N__20564\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__20567\,
            I => \c0.n1917\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__20564\,
            I => \c0.n1917\
        );

    \I__3806\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20556\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__20556\,
            I => \N__20552\
        );

    \I__3804\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__20552\,
            I => \N__20544\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20544\
        );

    \I__3801\ : Span4Mux_h
    port map (
            O => \N__20544\,
            I => \N__20538\
        );

    \I__3800\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20533\
        );

    \I__3799\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__3798\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20530\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__20538\,
            I => \c0.data_in_field_34\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__20533\,
            I => \c0.data_in_field_34\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__20530\,
            I => \c0.data_in_field_34\
        );

    \I__3794\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__20520\,
            I => \N__20517\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__20517\,
            I => \N__20513\
        );

    \I__3791\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20510\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__20510\,
            I => \N__20504\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__20507\,
            I => \c0.n2092\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__20504\,
            I => \c0.n2092\
        );

    \I__3786\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20496\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20492\
        );

    \I__3784\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20489\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__20492\,
            I => \N__20484\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20484\
        );

    \I__3781\ : Span4Mux_h
    port map (
            O => \N__20484\,
            I => \N__20481\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__20481\,
            I => \c0.n5527\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__20478\,
            I => \c0.n5394_cascade_\
        );

    \I__3778\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20472\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20468\
        );

    \I__3776\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20465\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__20468\,
            I => \N__20462\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20459\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__20462\,
            I => \N__20456\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__20459\,
            I => \N__20453\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__20456\,
            I => \c0.n1926\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__20453\,
            I => \c0.n1926\
        );

    \I__3769\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20445\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20442\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__20433\,
            I => \c0.n19_adj_1889\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__3762\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20424\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__20424\,
            I => \N__20421\
        );

    \I__3760\ : Odrv12
    port map (
            O => \N__20421\,
            I => \c0.n22_adj_1886\
        );

    \I__3759\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20413\
        );

    \I__3758\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20408\
        );

    \I__3757\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20405\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20399\
        );

    \I__3755\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20396\
        );

    \I__3754\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20393\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__20408\,
            I => \N__20388\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20388\
        );

    \I__3751\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20385\
        );

    \I__3750\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20382\
        );

    \I__3749\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20379\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__20399\,
            I => \r_Bit_Index_0\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__20396\,
            I => \r_Bit_Index_0\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__20393\,
            I => \r_Bit_Index_0\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__20388\,
            I => \r_Bit_Index_0\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__20385\,
            I => \r_Bit_Index_0\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__20382\,
            I => \r_Bit_Index_0\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__20379\,
            I => \r_Bit_Index_0\
        );

    \I__3741\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20356\
        );

    \I__3740\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20353\
        );

    \I__3739\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20350\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__20361\,
            I => \N__20346\
        );

    \I__3737\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20341\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__20359\,
            I => \N__20338\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20335\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__20353\,
            I => \N__20330\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__20350\,
            I => \N__20330\
        );

    \I__3732\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20327\
        );

    \I__3731\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20320\
        );

    \I__3730\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20320\
        );

    \I__3729\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20320\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20317\
        );

    \I__3727\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20313\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__20335\,
            I => \N__20304\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__20330\,
            I => \N__20304\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20304\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__20320\,
            I => \N__20304\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__20317\,
            I => \N__20301\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20296\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__20313\,
            I => \N__20293\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__20304\,
            I => \N__20290\
        );

    \I__3718\ : Sp12to4
    port map (
            O => \N__20301\,
            I => \N__20287\
        );

    \I__3717\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20284\
        );

    \I__3716\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20279\
        );

    \I__3715\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20279\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__20293\,
            I => \N__20276\
        );

    \I__3713\ : Span4Mux_s2_h
    port map (
            O => \N__20290\,
            I => \N__20273\
        );

    \I__3712\ : Span12Mux_v
    port map (
            O => \N__20287\,
            I => \N__20270\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__20284\,
            I => \N__20265\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20265\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__20276\,
            I => \r_Rx_Data\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__20273\,
            I => \r_Rx_Data\
        );

    \I__3707\ : Odrv12
    port map (
            O => \N__20270\,
            I => \r_Rx_Data\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__20265\,
            I => \r_Rx_Data\
        );

    \I__3705\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__20253\,
            I => n1757
        );

    \I__3703\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20246\
        );

    \I__3702\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20243\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20240\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__3699\ : Span4Mux_v
    port map (
            O => \N__20240\,
            I => \N__20230\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__20237\,
            I => \N__20230\
        );

    \I__3697\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20227\
        );

    \I__3696\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20224\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__20230\,
            I => \N__20221\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__20227\,
            I => \N__20218\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__20224\,
            I => data_in_3_6
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__20221\,
            I => data_in_3_6
        );

    \I__3691\ : Odrv12
    port map (
            O => \N__20218\,
            I => data_in_3_6
        );

    \I__3690\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20205\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__20205\,
            I => \N__20202\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__20202\,
            I => \N__20197\
        );

    \I__3686\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20194\
        );

    \I__3685\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20191\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__20197\,
            I => data_in_0_5
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__20194\,
            I => data_in_0_5
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__20191\,
            I => data_in_0_5
        );

    \I__3681\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__20178\,
            I => \c0.n22_adj_1924\
        );

    \I__3678\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20168\
        );

    \I__3676\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20165\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__20168\,
            I => \N__20160\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20157\
        );

    \I__3673\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20154\
        );

    \I__3672\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20151\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__20160\,
            I => \N__20147\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__20157\,
            I => \N__20142\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__20154\,
            I => \N__20142\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__20151\,
            I => \N__20139\
        );

    \I__3667\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20136\
        );

    \I__3666\ : Span4Mux_v
    port map (
            O => \N__20147\,
            I => \N__20129\
        );

    \I__3665\ : Span4Mux_h
    port map (
            O => \N__20142\,
            I => \N__20129\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__20139\,
            I => \N__20129\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__20136\,
            I => \c0.data_in_field_141\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__20129\,
            I => \c0.data_in_field_141\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__20124\,
            I => \N__20119\
        );

    \I__3660\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20113\
        );

    \I__3659\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20113\
        );

    \I__3658\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20110\
        );

    \I__3657\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20107\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20102\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20102\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__20107\,
            I => data_in_18_4
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__20102\,
            I => data_in_18_4
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__20097\,
            I => \c0.tx.n40_cascade_\
        );

    \I__3651\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20089\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20084\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20084\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__20089\,
            I => \N__20081\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__20084\,
            I => \N__20078\
        );

    \I__3646\ : Odrv12
    port map (
            O => \N__20081\,
            I => n1760
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__20078\,
            I => n1760
        );

    \I__3644\ : CEMux
    port map (
            O => \N__20073\,
            I => \N__20070\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__20070\,
            I => \N__20067\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__20067\,
            I => \N__20063\
        );

    \I__3641\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20060\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__20063\,
            I => \c0.tx.n2247\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__20060\,
            I => \c0.tx.n2247\
        );

    \I__3638\ : SRMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__20052\,
            I => \c0.tx.n2356\
        );

    \I__3636\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20046\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20040\
        );

    \I__3634\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20037\
        );

    \I__3633\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20034\
        );

    \I__3632\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20029\
        );

    \I__3631\ : Span4Mux_h
    port map (
            O => \N__20040\,
            I => \N__20026\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20023\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20020\
        );

    \I__3628\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20015\
        );

    \I__3627\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20015\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__20029\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__20026\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__20023\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__20020\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__20015\,
            I => \c0.rx.r_Bit_Index_2\
        );

    \I__3621\ : InMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__20001\,
            I => \N__19994\
        );

    \I__3619\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19991\
        );

    \I__3618\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19986\
        );

    \I__3617\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19983\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19980\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__19994\,
            I => \N__19977\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19974\
        );

    \I__3613\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19969\
        );

    \I__3612\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19969\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__19986\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__19983\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__19980\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__19977\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__19974\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__19969\,
            I => \c0.rx.r_Bit_Index_1\
        );

    \I__3605\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19948\
        );

    \I__3603\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19945\
        );

    \I__3602\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19942\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__19948\,
            I => \N__19939\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19936\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19933\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__19939\,
            I => \c0.rx.n1706\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__19936\,
            I => \c0.rx.n1706\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__19933\,
            I => \c0.rx.n1706\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__19926\,
            I => \n1757_cascade_\
        );

    \I__3594\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19920\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__19917\,
            I => \N__19913\
        );

    \I__3591\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19910\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__19913\,
            I => rx_data_0
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__19910\,
            I => rx_data_0
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19902\
        );

    \I__3587\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19899\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19894\
        );

    \I__3585\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19889\
        );

    \I__3584\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19889\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__19894\,
            I => data_in_12_1
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__19889\,
            I => data_in_12_1
        );

    \I__3581\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19881\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__19881\,
            I => \N__19876\
        );

    \I__3579\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19873\
        );

    \I__3578\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19870\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__19876\,
            I => \N__19864\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19864\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19861\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19857\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__19864\,
            I => \N__19854\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__19861\,
            I => \N__19851\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19848\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__19857\,
            I => \c0.data_in_field_97\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__19854\,
            I => \c0.data_in_field_97\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__19851\,
            I => \c0.data_in_field_97\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__19848\,
            I => \c0.data_in_field_97\
        );

    \I__3566\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__3564\ : Span4Mux_v
    port map (
            O => \N__19833\,
            I => \N__19829\
        );

    \I__3563\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19826\
        );

    \I__3562\ : Span4Mux_h
    port map (
            O => \N__19829\,
            I => \N__19823\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__19826\,
            I => \c0.data_in_frame_19_5\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__19823\,
            I => \c0.data_in_frame_19_5\
        );

    \I__3559\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__19815\,
            I => \N__19811\
        );

    \I__3557\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19808\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__19811\,
            I => \N__19804\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19801\
        );

    \I__3554\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19798\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__19804\,
            I => data_in_14_6
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__19801\,
            I => data_in_14_6
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__19798\,
            I => data_in_14_6
        );

    \I__3550\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19786\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__19790\,
            I => \N__19783\
        );

    \I__3548\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19779\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19776\
        );

    \I__3546\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19773\
        );

    \I__3545\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19770\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__19779\,
            I => \N__19767\
        );

    \I__3543\ : Span4Mux_v
    port map (
            O => \N__19776\,
            I => \N__19764\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__19773\,
            I => \N__19761\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__19770\,
            I => data_in_19_7
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__19767\,
            I => data_in_19_7
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__19764\,
            I => data_in_19_7
        );

    \I__3538\ : Odrv12
    port map (
            O => \N__19761\,
            I => data_in_19_7
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19746\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__19746\,
            I => \N__19742\
        );

    \I__3534\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19739\
        );

    \I__3533\ : Span4Mux_s3_h
    port map (
            O => \N__19742\,
            I => \N__19736\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__19739\,
            I => \c0.data_in_frame_19_7\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__19736\,
            I => \c0.data_in_frame_19_7\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__19731\,
            I => \N__19726\
        );

    \I__3529\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19721\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19721\
        );

    \I__3527\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19718\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19715\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__19718\,
            I => \N__19711\
        );

    \I__3524\ : Span4Mux_h
    port map (
            O => \N__19715\,
            I => \N__19708\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19705\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__19711\,
            I => \N__19702\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__19708\,
            I => data_in_19_5
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19705\,
            I => data_in_19_5
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__19702\,
            I => data_in_19_5
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__19695\,
            I => \N__19692\
        );

    \I__3517\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19684\
        );

    \I__3515\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19681\
        );

    \I__3514\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19678\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__19684\,
            I => data_in_14_0
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__19681\,
            I => data_in_14_0
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__19678\,
            I => data_in_14_0
        );

    \I__3510\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19667\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19664\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19661\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19658\
        );

    \I__3506\ : Span12Mux_v
    port map (
            O => \N__19661\,
            I => \N__19654\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19651\
        );

    \I__3504\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19648\
        );

    \I__3503\ : Odrv12
    port map (
            O => \N__19654\,
            I => data_in_13_0
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__19651\,
            I => data_in_13_0
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__19648\,
            I => data_in_13_0
        );

    \I__3500\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19636\
        );

    \I__3499\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19633\
        );

    \I__3498\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19630\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__19636\,
            I => \N__19627\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__19633\,
            I => \N__19624\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__19630\,
            I => \N__19621\
        );

    \I__3494\ : Span4Mux_s2_h
    port map (
            O => \N__19627\,
            I => \N__19618\
        );

    \I__3493\ : Span12Mux_s6_h
    port map (
            O => \N__19624\,
            I => \N__19613\
        );

    \I__3492\ : Span4Mux_v
    port map (
            O => \N__19621\,
            I => \N__19610\
        );

    \I__3491\ : Span4Mux_h
    port map (
            O => \N__19618\,
            I => \N__19607\
        );

    \I__3490\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19602\
        );

    \I__3489\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19602\
        );

    \I__3488\ : Odrv12
    port map (
            O => \N__19613\,
            I => \c0.data_in_field_36\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__19610\,
            I => \c0.data_in_field_36\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__19607\,
            I => \c0.data_in_field_36\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__19602\,
            I => \c0.data_in_field_36\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19586\
        );

    \I__3482\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19583\
        );

    \I__3481\ : Span4Mux_s2_h
    port map (
            O => \N__19586\,
            I => \N__19579\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19576\
        );

    \I__3479\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19572\
        );

    \I__3478\ : Span4Mux_h
    port map (
            O => \N__19579\,
            I => \N__19567\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19567\
        );

    \I__3476\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19564\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__19572\,
            I => \c0.data_in_field_82\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__19567\,
            I => \c0.data_in_field_82\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__19564\,
            I => \c0.data_in_field_82\
        );

    \I__3472\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__19554\,
            I => \N__19550\
        );

    \I__3470\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19546\
        );

    \I__3469\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19543\
        );

    \I__3468\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19540\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__19546\,
            I => \c0.n1948\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__19543\,
            I => \c0.n1948\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__19540\,
            I => \c0.n1948\
        );

    \I__3464\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__19530\,
            I => \N__19526\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \N__19523\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__3460\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19516\
        );

    \I__3459\ : Span4Mux_h
    port map (
            O => \N__19520\,
            I => \N__19513\
        );

    \I__3458\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19510\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__19516\,
            I => data_in_15_1
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__19513\,
            I => data_in_15_1
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__19510\,
            I => data_in_15_1
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__3453\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19496\
        );

    \I__3452\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19493\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19490\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__19493\,
            I => \N__19487\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__19490\,
            I => \N__19481\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__19487\,
            I => \N__19481\
        );

    \I__3447\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19478\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__19481\,
            I => data_in_14_1
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__19478\,
            I => data_in_14_1
        );

    \I__3444\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__19470\,
            I => \N__19465\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__19469\,
            I => \N__19462\
        );

    \I__3441\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19458\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__19465\,
            I => \N__19455\
        );

    \I__3439\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19450\
        );

    \I__3438\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19450\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__19458\,
            I => \c0.data_in_field_127\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__19455\,
            I => \c0.data_in_field_127\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__19450\,
            I => \c0.data_in_field_127\
        );

    \I__3434\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19440\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N__19436\
        );

    \I__3432\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19433\
        );

    \I__3431\ : Sp12to4
    port map (
            O => \N__19436\,
            I => \N__19430\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__3429\ : Span12Mux_v
    port map (
            O => \N__19430\,
            I => \N__19424\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__19427\,
            I => \N__19421\
        );

    \I__3427\ : Odrv12
    port map (
            O => \N__19424\,
            I => n4
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__19421\,
            I => n4
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__3424\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19410\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__3422\ : Span4Mux_h
    port map (
            O => \N__19407\,
            I => \N__19402\
        );

    \I__3421\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19397\
        );

    \I__3420\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19397\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__19402\,
            I => data_in_13_1
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__19397\,
            I => data_in_13_1
        );

    \I__3417\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19389\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__19389\,
            I => \N__19385\
        );

    \I__3415\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19382\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__19385\,
            I => \N__19377\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19377\
        );

    \I__3412\ : Span4Mux_h
    port map (
            O => \N__19377\,
            I => \N__19373\
        );

    \I__3411\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19370\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__19373\,
            I => \N__19367\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__19370\,
            I => \c0.data_in_field_105\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__19367\,
            I => \c0.data_in_field_105\
        );

    \I__3407\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19359\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__19359\,
            I => \c0.n18_adj_1887\
        );

    \I__3405\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19353\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19350\
        );

    \I__3403\ : Span4Mux_s3_h
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__19344\,
            I => \c0.n20_adj_1888\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__19341\,
            I => \c0.tx2_transmit_N_1031_cascade_\
        );

    \I__3399\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19333\
        );

    \I__3398\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19328\
        );

    \I__3397\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19328\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__19333\,
            I => \c0.data_in_field_29\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__19328\,
            I => \c0.data_in_field_29\
        );

    \I__3394\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__3392\ : Odrv12
    port map (
            O => \N__19317\,
            I => \c0.n2030\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__19314\,
            I => \c0.n2030_cascade_\
        );

    \I__3390\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19308\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__19302\,
            I => \N__19298\
        );

    \I__3386\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19295\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__19298\,
            I => \N__19289\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19289\
        );

    \I__3383\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19286\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__19289\,
            I => data_in_15_2
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__19286\,
            I => data_in_15_2
        );

    \I__3380\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__19275\,
            I => \N__19270\
        );

    \I__3377\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19265\
        );

    \I__3376\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19265\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__19270\,
            I => \c0.data_in_field_22\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__19265\,
            I => \c0.data_in_field_22\
        );

    \I__3373\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19254\
        );

    \I__3371\ : Span4Mux_v
    port map (
            O => \N__19254\,
            I => \N__19251\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__19251\,
            I => \c0.n5436\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__19248\,
            I => \c0.n5436_cascade_\
        );

    \I__3368\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__19242\,
            I => \c0.n5509\
        );

    \I__3366\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19229\
        );

    \I__3364\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19226\
        );

    \I__3363\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19219\
        );

    \I__3362\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19219\
        );

    \I__3361\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19219\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__19229\,
            I => \c0.data_in_field_78\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__19226\,
            I => \c0.data_in_field_78\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__19219\,
            I => \c0.data_in_field_78\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__19212\,
            I => \c0.n5509_cascade_\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__19209\,
            I => \N__19203\
        );

    \I__3355\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19200\
        );

    \I__3354\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19197\
        );

    \I__3353\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19192\
        );

    \I__3352\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19192\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19185\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__19197\,
            I => \N__19185\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19182\
        );

    \I__3348\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19179\
        );

    \I__3347\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19176\
        );

    \I__3346\ : Span4Mux_v
    port map (
            O => \N__19185\,
            I => \N__19171\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__19182\,
            I => \N__19171\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__19179\,
            I => \c0.data_in_field_92\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__19176\,
            I => \c0.data_in_field_92\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__19171\,
            I => \c0.data_in_field_92\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__19164\,
            I => \N__19160\
        );

    \I__3340\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19156\
        );

    \I__3339\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19153\
        );

    \I__3338\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19150\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__19156\,
            I => \c0.data_in_field_52\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__19153\,
            I => \c0.data_in_field_52\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__19150\,
            I => \c0.data_in_field_52\
        );

    \I__3334\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__3332\ : Span4Mux_h
    port map (
            O => \N__19137\,
            I => \N__19133\
        );

    \I__3331\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19129\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__19133\,
            I => \N__19126\
        );

    \I__3329\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19123\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__19129\,
            I => \c0.data_in_field_103\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__19126\,
            I => \c0.data_in_field_103\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__19123\,
            I => \c0.data_in_field_103\
        );

    \I__3325\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19113\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__19113\,
            I => \c0.n2152\
        );

    \I__3323\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19102\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19098\
        );

    \I__3320\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19095\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__19102\,
            I => \N__19092\
        );

    \I__3318\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19089\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19084\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__19095\,
            I => \N__19084\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__19092\,
            I => \c0.data_in_field_43\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__19089\,
            I => \c0.data_in_field_43\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__19084\,
            I => \c0.data_in_field_43\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__19077\,
            I => \c0.n2152_cascade_\
        );

    \I__3311\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19071\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__19071\,
            I => \N__19067\
        );

    \I__3309\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19064\
        );

    \I__3308\ : Span4Mux_h
    port map (
            O => \N__19067\,
            I => \N__19061\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__19064\,
            I => \N__19058\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__19061\,
            I => \c0.n5397\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__19058\,
            I => \c0.n5397\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__3303\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__19044\,
            I => \N__19039\
        );

    \I__3300\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19036\
        );

    \I__3299\ : InMux
    port map (
            O => \N__19042\,
            I => \N__19033\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__19039\,
            I => data_in_11_6
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__19036\,
            I => data_in_11_6
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__19033\,
            I => data_in_11_6
        );

    \I__3295\ : InMux
    port map (
            O => \N__19026\,
            I => \N__19023\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__19023\,
            I => \N__19017\
        );

    \I__3293\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19014\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \N__19011\
        );

    \I__3291\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19008\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__19017\,
            I => \N__19005\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__19014\,
            I => \N__19002\
        );

    \I__3288\ : InMux
    port map (
            O => \N__19011\,
            I => \N__18999\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__19008\,
            I => \c0.data_in_field_75\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__19005\,
            I => \c0.data_in_field_75\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__19002\,
            I => \c0.data_in_field_75\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__18999\,
            I => \c0.data_in_field_75\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__18990\,
            I => \N__18987\
        );

    \I__3282\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__3280\ : Sp12to4
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__3279\ : Span12Mux_v
    port map (
            O => \N__18978\,
            I => \N__18973\
        );

    \I__3278\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18968\
        );

    \I__3277\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18968\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__18973\,
            I => data_in_17_6
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__18968\,
            I => data_in_17_6
        );

    \I__3274\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18959\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__18962\,
            I => \N__18955\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__18959\,
            I => \N__18952\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__18958\,
            I => \N__18949\
        );

    \I__3270\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18946\
        );

    \I__3269\ : Span4Mux_v
    port map (
            O => \N__18952\,
            I => \N__18941\
        );

    \I__3268\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18938\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__18946\,
            I => \N__18935\
        );

    \I__3266\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18930\
        );

    \I__3265\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18930\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__18941\,
            I => \c0.data_in_field_142\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__18938\,
            I => \c0.data_in_field_142\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__18935\,
            I => \c0.data_in_field_142\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__18930\,
            I => \c0.data_in_field_142\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__3259\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18915\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__18915\,
            I => \N__18911\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18906\
        );

    \I__3256\ : Span12Mux_s6_h
    port map (
            O => \N__18911\,
            I => \N__18903\
        );

    \I__3255\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18898\
        );

    \I__3254\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18898\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18895\
        );

    \I__3252\ : Odrv12
    port map (
            O => \N__18903\,
            I => \c0.data_in_field_33\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__18898\,
            I => \c0.data_in_field_33\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__18895\,
            I => \c0.data_in_field_33\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__18882\,
            I => \N__18878\
        );

    \I__3246\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18873\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__18878\,
            I => \N__18870\
        );

    \I__3244\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18867\
        );

    \I__3243\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18864\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__18873\,
            I => \c0.data_in_field_140\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__18870\,
            I => \c0.data_in_field_140\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__18867\,
            I => \c0.data_in_field_140\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__18864\,
            I => \c0.data_in_field_140\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18851\
        );

    \I__3237\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18848\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__18851\,
            I => \N__18845\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__18848\,
            I => \N__18842\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__18845\,
            I => \N__18836\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__18842\,
            I => \N__18836\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18833\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__18836\,
            I => data_in_12_7
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__18833\,
            I => data_in_12_7
        );

    \I__3229\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__18825\,
            I => \N__18820\
        );

    \I__3227\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18817\
        );

    \I__3226\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18814\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__18820\,
            I => \N__18809\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18804\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18804\
        );

    \I__3222\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18799\
        );

    \I__3221\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18799\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__18809\,
            I => \c0.data_in_field_126\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__18804\,
            I => \c0.data_in_field_126\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__18799\,
            I => \c0.data_in_field_126\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__18792\,
            I => \N__18786\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__18791\,
            I => \N__18783\
        );

    \I__3215\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18780\
        );

    \I__3214\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18777\
        );

    \I__3213\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18774\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18771\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__18780\,
            I => \N__18768\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18763\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__18774\,
            I => \N__18763\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__18771\,
            I => \N__18758\
        );

    \I__3207\ : Span4Mux_h
    port map (
            O => \N__18768\,
            I => \N__18758\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__18763\,
            I => \N__18755\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__18758\,
            I => \c0.data_in_field_118\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__18755\,
            I => \c0.data_in_field_118\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18744\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18744\,
            I => \N__18740\
        );

    \I__3200\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18737\
        );

    \I__3199\ : Span4Mux_s2_h
    port map (
            O => \N__18740\,
            I => \N__18733\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18730\
        );

    \I__3197\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18727\
        );

    \I__3196\ : Span4Mux_h
    port map (
            O => \N__18733\,
            I => \N__18719\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__18730\,
            I => \N__18719\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18719\
        );

    \I__3193\ : InMux
    port map (
            O => \N__18726\,
            I => \N__18715\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__18719\,
            I => \N__18712\
        );

    \I__3191\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18709\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__18715\,
            I => \c0.data_in_field_51\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__18712\,
            I => \c0.data_in_field_51\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__18709\,
            I => \c0.data_in_field_51\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__18702\,
            I => \N__18699\
        );

    \I__3186\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__18696\,
            I => \N__18691\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18686\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18686\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__18691\,
            I => data_in_16_5
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18686\,
            I => data_in_16_5
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__3179\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__18672\,
            I => \N__18667\
        );

    \I__3176\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18664\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18661\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__18667\,
            I => data_in_9_3
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__18664\,
            I => data_in_9_3
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__18661\,
            I => data_in_9_3
        );

    \I__3171\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18650\
        );

    \I__3170\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18647\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__18650\,
            I => \N__18641\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18641\
        );

    \I__3167\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18637\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__18641\,
            I => \N__18634\
        );

    \I__3165\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18631\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__18637\,
            I => \c0.data_in_field_3\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__18634\,
            I => \c0.data_in_field_3\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__18631\,
            I => \c0.data_in_field_3\
        );

    \I__3161\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18621\,
            I => \N__18617\
        );

    \I__3159\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18614\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__18617\,
            I => \c0.n2125\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__18614\,
            I => \c0.n2125\
        );

    \I__3156\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18606\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18602\
        );

    \I__3154\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18598\
        );

    \I__3153\ : Span4Mux_v
    port map (
            O => \N__18602\,
            I => \N__18595\
        );

    \I__3152\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18592\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__18598\,
            I => \c0.data_in_field_27\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__18595\,
            I => \c0.data_in_field_27\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__18592\,
            I => \c0.data_in_field_27\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__18582\,
            I => \c0.n5469\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__18579\,
            I => \N__18574\
        );

    \I__3145\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18569\
        );

    \I__3144\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18566\
        );

    \I__3143\ : InMux
    port map (
            O => \N__18574\,
            I => \N__18563\
        );

    \I__3142\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18560\
        );

    \I__3141\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18557\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18552\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18552\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18547\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18547\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__18557\,
            I => \c0.data_in_field_83\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__18552\,
            I => \c0.data_in_field_83\
        );

    \I__3134\ : Odrv12
    port map (
            O => \N__18547\,
            I => \c0.data_in_field_83\
        );

    \I__3133\ : InMux
    port map (
            O => \N__18540\,
            I => \N__18537\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__18537\,
            I => \N__18534\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__3130\ : Span4Mux_h
    port map (
            O => \N__18531\,
            I => \N__18528\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__18528\,
            I => \c0.n5454\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__18525\,
            I => \c0.n5469_cascade_\
        );

    \I__3127\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18519\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__18519\,
            I => \c0.n6_adj_1923\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__18516\,
            I => \c0.n5548_cascade_\
        );

    \I__3124\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18510\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__18510\,
            I => \N__18505\
        );

    \I__3122\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18500\
        );

    \I__3121\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18500\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__18505\,
            I => data_in_0_4
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__18500\,
            I => data_in_0_4
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__18495\,
            I => \N__18492\
        );

    \I__3117\ : InMux
    port map (
            O => \N__18492\,
            I => \N__18489\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__18489\,
            I => \N__18484\
        );

    \I__3115\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18479\
        );

    \I__3114\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18479\
        );

    \I__3113\ : Odrv12
    port map (
            O => \N__18484\,
            I => data_in_7_5
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__18479\,
            I => data_in_7_5
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__18474\,
            I => \c0.n1729_cascade_\
        );

    \I__3110\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18467\
        );

    \I__3109\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18461\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__18467\,
            I => \N__18458\
        );

    \I__3107\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18455\
        );

    \I__3106\ : InMux
    port map (
            O => \N__18465\,
            I => \N__18452\
        );

    \I__3105\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18449\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__18461\,
            I => \N__18446\
        );

    \I__3103\ : Span12Mux_v
    port map (
            O => \N__18458\,
            I => \N__18441\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__18455\,
            I => \N__18441\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__18452\,
            I => \c0.data_in_field_35\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__18449\,
            I => \c0.data_in_field_35\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__18446\,
            I => \c0.data_in_field_35\
        );

    \I__3098\ : Odrv12
    port map (
            O => \N__18441\,
            I => \c0.data_in_field_35\
        );

    \I__3097\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18427\
        );

    \I__3096\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18424\
        );

    \I__3095\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18420\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__18427\,
            I => \N__18417\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18414\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__18423\,
            I => \N__18411\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18408\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__18417\,
            I => \N__18403\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__18414\,
            I => \N__18403\
        );

    \I__3088\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18399\
        );

    \I__3087\ : Span4Mux_h
    port map (
            O => \N__18408\,
            I => \N__18396\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__18403\,
            I => \N__18393\
        );

    \I__3085\ : InMux
    port map (
            O => \N__18402\,
            I => \N__18390\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__18399\,
            I => \c0.data_in_field_9\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__18396\,
            I => \c0.data_in_field_9\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__18393\,
            I => \c0.data_in_field_9\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__18390\,
            I => \c0.data_in_field_9\
        );

    \I__3080\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18377\
        );

    \I__3079\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18374\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__3076\ : Span4Mux_s3_h
    port map (
            O => \N__18371\,
            I => \N__18365\
        );

    \I__3075\ : Span4Mux_v
    port map (
            O => \N__18368\,
            I => \N__18362\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__18365\,
            I => \N__18359\
        );

    \I__3073\ : Span4Mux_h
    port map (
            O => \N__18362\,
            I => \N__18354\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__18359\,
            I => \N__18351\
        );

    \I__3071\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18346\
        );

    \I__3070\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18346\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__18354\,
            I => \c0.data_in_field_54\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__18351\,
            I => \c0.data_in_field_54\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__18346\,
            I => \c0.data_in_field_54\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__18339\,
            I => \c0.n5369_cascade_\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__3064\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18325\
        );

    \I__3062\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18322\
        );

    \I__3061\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18319\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__18325\,
            I => data_in_0_3
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__18322\,
            I => data_in_0_3
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__18319\,
            I => data_in_0_3
        );

    \I__3057\ : InMux
    port map (
            O => \N__18312\,
            I => \N__18309\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__18309\,
            I => \c0.n26\
        );

    \I__3055\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__18303\,
            I => \c0.n27_adj_1928\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__18300\,
            I => \c0.n28_adj_1926_cascade_\
        );

    \I__3052\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__18294\,
            I => \c0.n25_adj_1929\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__18291\,
            I => \N__18287\
        );

    \I__3049\ : InMux
    port map (
            O => \N__18290\,
            I => \N__18283\
        );

    \I__3048\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18280\
        );

    \I__3047\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18276\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__18283\,
            I => \N__18273\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18270\
        );

    \I__3044\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18267\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18262\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__18273\,
            I => \N__18262\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__18270\,
            I => \N__18259\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__18267\,
            I => data_in_2_1
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__18262\,
            I => data_in_2_1
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__18259\,
            I => data_in_2_1
        );

    \I__3037\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18249\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18245\
        );

    \I__3035\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18242\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__18245\,
            I => \N__18237\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18237\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__18237\,
            I => \N__18232\
        );

    \I__3031\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18229\
        );

    \I__3030\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18226\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__18232\,
            I => data_in_1_0
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__18229\,
            I => data_in_1_0
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__18226\,
            I => data_in_1_0
        );

    \I__3026\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18216\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__18216\,
            I => \N__18213\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__18213\,
            I => \N__18208\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18203\
        );

    \I__3022\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18203\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__18208\,
            I => data_in_0_6
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__18203\,
            I => data_in_0_6
        );

    \I__3019\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18190\
        );

    \I__3017\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18187\
        );

    \I__3016\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18183\
        );

    \I__3015\ : Span4Mux_v
    port map (
            O => \N__18190\,
            I => \N__18180\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__18187\,
            I => \N__18177\
        );

    \I__3013\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18174\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18171\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__18180\,
            I => data_in_3_7
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__18177\,
            I => data_in_3_7
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__18174\,
            I => data_in_3_7
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__18171\,
            I => data_in_3_7
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__18162\,
            I => \N__18159\
        );

    \I__3006\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__18156\,
            I => \N__18153\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__18153\,
            I => \N__18147\
        );

    \I__3003\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18140\
        );

    \I__3002\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18140\
        );

    \I__3001\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18140\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__18147\,
            I => data_in_1_6
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__18140\,
            I => data_in_1_6
        );

    \I__2998\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18128\
        );

    \I__2997\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18128\
        );

    \I__2996\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18125\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__18128\,
            I => \N__18122\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__18125\,
            I => \N__18116\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__18122\,
            I => \N__18116\
        );

    \I__2992\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18113\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__18116\,
            I => \N__18110\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__18113\,
            I => data_in_1_7
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__18110\,
            I => data_in_1_7
        );

    \I__2988\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18101\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__18104\,
            I => \N__18097\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18094\
        );

    \I__2985\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18089\
        );

    \I__2984\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18089\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__18094\,
            I => data_in_0_7
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__18089\,
            I => data_in_0_7
        );

    \I__2981\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18081\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__18081\,
            I => \c0.n30_adj_1941\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18075\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__18075\,
            I => \c0.n4795\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__18072\,
            I => \N__18069\
        );

    \I__2976\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18066\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__18066\,
            I => \c0.n26_adj_1940\
        );

    \I__2974\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18060\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__18060\,
            I => \c0.rx.n5633\
        );

    \I__2972\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18053\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18050\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__18053\,
            I => \N__18047\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18044\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__18047\,
            I => n3636
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__18044\,
            I => n3636
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__2965\ : InMux
    port map (
            O => \N__18036\,
            I => \N__18032\
        );

    \I__2964\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18029\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__18032\,
            I => \c0.rx.n3850\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__18029\,
            I => \c0.rx.n3850\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__18019\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \N__18013\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18010\
        );

    \I__2958\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18007\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__18018\,
            I => \N__18000\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__17997\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__18016\,
            I => \N__17993\
        );

    \I__2954\ : InMux
    port map (
            O => \N__18013\,
            I => \N__17987\
        );

    \I__2953\ : InMux
    port map (
            O => \N__18010\,
            I => \N__17987\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__17984\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__18006\,
            I => \N__17980\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__18005\,
            I => \N__17977\
        );

    \I__2949\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17974\
        );

    \I__2948\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17967\
        );

    \I__2947\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17967\
        );

    \I__2946\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17967\
        );

    \I__2945\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17962\
        );

    \I__2944\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17962\
        );

    \I__2943\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17959\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__17987\,
            I => \N__17956\
        );

    \I__2941\ : Span4Mux_h
    port map (
            O => \N__17984\,
            I => \N__17953\
        );

    \I__2940\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17946\
        );

    \I__2939\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17946\
        );

    \I__2938\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17946\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__17974\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__17967\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__17962\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__17959\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__17956\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__17953\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__17946\,
            I => \r_SM_Main_1_adj_1990\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__17931\,
            I => \c0.rx.n3850_cascade_\
        );

    \I__2929\ : CEMux
    port map (
            O => \N__17928\,
            I => \N__17924\
        );

    \I__2928\ : CEMux
    port map (
            O => \N__17927\,
            I => \N__17921\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17915\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__17918\,
            I => \N__17911\
        );

    \I__2924\ : Span4Mux_v
    port map (
            O => \N__17915\,
            I => \N__17908\
        );

    \I__2923\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17905\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__17911\,
            I => \c0.rx.n2259\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__17908\,
            I => \c0.rx.n2259\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__17905\,
            I => \c0.rx.n2259\
        );

    \I__2919\ : SRMux
    port map (
            O => \N__17898\,
            I => \N__17894\
        );

    \I__2918\ : SRMux
    port map (
            O => \N__17897\,
            I => \N__17891\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17888\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17885\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__17888\,
            I => \N__17880\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__17885\,
            I => \N__17880\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__17880\,
            I => \c0.rx.n2367\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__17877\,
            I => \N__17874\
        );

    \I__2911\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17871\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17866\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \N__17862\
        );

    \I__2908\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17859\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__17866\,
            I => \N__17856\
        );

    \I__2906\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17851\
        );

    \I__2905\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17851\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17859\,
            I => data_in_2_5
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__17856\,
            I => data_in_2_5
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__17851\,
            I => data_in_2_5
        );

    \I__2901\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__2899\ : Span4Mux_v
    port map (
            O => \N__17838\,
            I => \N__17833\
        );

    \I__2898\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17828\
        );

    \I__2897\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17828\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__17833\,
            I => \N__17825\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__17828\,
            I => data_in_10_1
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__17825\,
            I => data_in_10_1
        );

    \I__2893\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17816\
        );

    \I__2892\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17813\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17810\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__17813\,
            I => \N__17805\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__17810\,
            I => \N__17805\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__17805\,
            I => \N__17801\
        );

    \I__2887\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17798\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__17801\,
            I => data_in_9_1
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__17798\,
            I => data_in_9_1
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \N__17790\
        );

    \I__2883\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17787\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__17787\,
            I => \N__17784\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__17784\,
            I => \N__17779\
        );

    \I__2880\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17774\
        );

    \I__2879\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17774\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__17779\,
            I => data_in_12_6
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__17774\,
            I => data_in_12_6
        );

    \I__2876\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17766\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17766\,
            I => \N__17763\
        );

    \I__2874\ : Span4Mux_v
    port map (
            O => \N__17763\,
            I => \N__17760\
        );

    \I__2873\ : Span4Mux_v
    port map (
            O => \N__17760\,
            I => \N__17756\
        );

    \I__2872\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__17756\,
            I => n1764
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__17753\,
            I => n1764
        );

    \I__2869\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17744\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17738\
        );

    \I__2866\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17735\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__17738\,
            I => rx_data_7
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__17735\,
            I => rx_data_7
        );

    \I__2863\ : InMux
    port map (
            O => \N__17730\,
            I => \N__17727\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__17727\,
            I => \N__17723\
        );

    \I__2861\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17720\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__17723\,
            I => \N__17717\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17714\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__17717\,
            I => \N__17709\
        );

    \I__2857\ : Span4Mux_h
    port map (
            O => \N__17714\,
            I => \N__17709\
        );

    \I__2856\ : Span4Mux_h
    port map (
            O => \N__17709\,
            I => \N__17705\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17702\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__17705\,
            I => data_in_15_6
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__17702\,
            I => data_in_15_6
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__17697\,
            I => \N__17692\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__17696\,
            I => \N__17685\
        );

    \I__2850\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17680\
        );

    \I__2849\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17675\
        );

    \I__2848\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17675\
        );

    \I__2847\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17670\
        );

    \I__2846\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17670\
        );

    \I__2845\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17667\
        );

    \I__2844\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17660\
        );

    \I__2843\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17660\
        );

    \I__2842\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17660\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__17680\,
            I => \N__17655\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__17675\,
            I => \N__17655\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__17670\,
            I => \r_SM_Main_0_adj_1991\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__17667\,
            I => \r_SM_Main_0_adj_1991\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__17660\,
            I => \r_SM_Main_0_adj_1991\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__17655\,
            I => \r_SM_Main_0_adj_1991\
        );

    \I__2835\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17642\
        );

    \I__2834\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17639\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__17642\,
            I => \N__17631\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17627\
        );

    \I__2831\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17622\
        );

    \I__2830\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17622\
        );

    \I__2829\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17615\
        );

    \I__2828\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17615\
        );

    \I__2827\ : InMux
    port map (
            O => \N__17634\,
            I => \N__17615\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__17631\,
            I => \N__17612\
        );

    \I__2825\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17609\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__17627\,
            I => \r_SM_Main_2_N_1824_2\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__17622\,
            I => \r_SM_Main_2_N_1824_2\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__17615\,
            I => \r_SM_Main_2_N_1824_2\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__17612\,
            I => \r_SM_Main_2_N_1824_2\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__17609\,
            I => \r_SM_Main_2_N_1824_2\
        );

    \I__2819\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17595\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__17595\,
            I => \c0.rx.n6291\
        );

    \I__2817\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17589\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__17589\,
            I => \N__17585\
        );

    \I__2815\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17582\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__17585\,
            I => \c0.n1889\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__17582\,
            I => \c0.n1889\
        );

    \I__2812\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17573\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \N__17570\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17567\
        );

    \I__2809\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17561\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__17567\,
            I => \N__17558\
        );

    \I__2807\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17551\
        );

    \I__2806\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17551\
        );

    \I__2805\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17551\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__17561\,
            I => \c0.data_in_field_76\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__17558\,
            I => \c0.data_in_field_76\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__17551\,
            I => \c0.data_in_field_76\
        );

    \I__2801\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17540\
        );

    \I__2800\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17537\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17534\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__17537\,
            I => \c0.data_in_frame_18_4\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__17534\,
            I => \c0.data_in_frame_18_4\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__17529\,
            I => \c0.n6243_cascade_\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__17526\,
            I => \c0.n5698_cascade_\
        );

    \I__2794\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17520\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__17520\,
            I => \N__17517\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__17517\,
            I => \c0.n6231\
        );

    \I__2791\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17511\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__17511\,
            I => \c0.n6237\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__17508\,
            I => \N__17505\
        );

    \I__2788\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17501\
        );

    \I__2787\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17496\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__17501\,
            I => \N__17493\
        );

    \I__2785\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17488\
        );

    \I__2784\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17488\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__17496\,
            I => \c0.data_in_field_102\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__17493\,
            I => \c0.data_in_field_102\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__17488\,
            I => \c0.data_in_field_102\
        );

    \I__2780\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__17478\,
            I => \c0.n5701\
        );

    \I__2778\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17471\
        );

    \I__2777\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17468\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__17471\,
            I => \N__17465\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__17468\,
            I => \N__17462\
        );

    \I__2774\ : Span4Mux_v
    port map (
            O => \N__17465\,
            I => \N__17458\
        );

    \I__2773\ : Span12Mux_v
    port map (
            O => \N__17462\,
            I => \N__17455\
        );

    \I__2772\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17452\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__17458\,
            I => data_in_10_6
        );

    \I__2770\ : Odrv12
    port map (
            O => \N__17455\,
            I => data_in_10_6
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__17452\,
            I => data_in_10_6
        );

    \I__2768\ : InMux
    port map (
            O => \N__17445\,
            I => \N__17442\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__17442\,
            I => \N__17436\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17432\
        );

    \I__2765\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17427\
        );

    \I__2764\ : InMux
    port map (
            O => \N__17439\,
            I => \N__17427\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__17436\,
            I => \N__17424\
        );

    \I__2762\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17421\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17418\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__17427\,
            I => \c0.data_in_field_86\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__17424\,
            I => \c0.data_in_field_86\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__17421\,
            I => \c0.data_in_field_86\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__17418\,
            I => \c0.data_in_field_86\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__17409\,
            I => \N__17406\
        );

    \I__2755\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__17403\,
            I => \c0.n5388\
        );

    \I__2753\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17397\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__17397\,
            I => \c0.n5418\
        );

    \I__2751\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17391\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__17391\,
            I => \N__17387\
        );

    \I__2749\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17384\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__17387\,
            I => \c0.n5491\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__17384\,
            I => \c0.n5491\
        );

    \I__2746\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17376\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__17376\,
            I => \c0.n44_adj_1894\
        );

    \I__2744\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17368\
        );

    \I__2743\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17365\
        );

    \I__2742\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17362\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__17368\,
            I => \c0.data_in_field_112\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__17365\,
            I => \c0.data_in_field_112\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__17362\,
            I => \c0.data_in_field_112\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__17355\,
            I => \N__17350\
        );

    \I__2737\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17347\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \N__17343\
        );

    \I__2735\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17340\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__17347\,
            I => \N__17337\
        );

    \I__2733\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17334\
        );

    \I__2732\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17331\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__17340\,
            I => \c0.data_in_field_30\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__17337\,
            I => \c0.data_in_field_30\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__17334\,
            I => \c0.data_in_field_30\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__17331\,
            I => \c0.data_in_field_30\
        );

    \I__2727\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17315\
        );

    \I__2725\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17312\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__17315\,
            I => \N__17304\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17304\
        );

    \I__2722\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17301\
        );

    \I__2721\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17296\
        );

    \I__2720\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17296\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__17304\,
            I => \c0.data_in_field_125\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__17301\,
            I => \c0.data_in_field_125\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__17296\,
            I => \c0.data_in_field_125\
        );

    \I__2716\ : InMux
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__17286\,
            I => \N__17280\
        );

    \I__2714\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17277\
        );

    \I__2713\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17274\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__17283\,
            I => \N__17270\
        );

    \I__2711\ : Span4Mux_s2_h
    port map (
            O => \N__17280\,
            I => \N__17265\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__17277\,
            I => \N__17265\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__17274\,
            I => \N__17262\
        );

    \I__2708\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17259\
        );

    \I__2707\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17256\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__17265\,
            I => \N__17253\
        );

    \I__2705\ : Span4Mux_h
    port map (
            O => \N__17262\,
            I => \N__17248\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17248\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__17256\,
            I => \c0.data_in_field_135\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__17253\,
            I => \c0.data_in_field_135\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__17248\,
            I => \c0.data_in_field_135\
        );

    \I__2700\ : InMux
    port map (
            O => \N__17241\,
            I => \N__17238\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__17238\,
            I => \N__17234\
        );

    \I__2698\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17231\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__17234\,
            I => \N__17228\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__17231\,
            I => \c0.n1908\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__17228\,
            I => \c0.n1908\
        );

    \I__2694\ : InMux
    port map (
            O => \N__17223\,
            I => \N__17220\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17220\,
            I => \N__17216\
        );

    \I__2692\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17213\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__17216\,
            I => \N__17204\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17204\
        );

    \I__2689\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17201\
        );

    \I__2688\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17198\
        );

    \I__2687\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17195\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__17209\,
            I => \N__17192\
        );

    \I__2685\ : Span4Mux_v
    port map (
            O => \N__17204\,
            I => \N__17187\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__17201\,
            I => \N__17187\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17182\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__17195\,
            I => \N__17182\
        );

    \I__2681\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17179\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__17187\,
            I => \N__17176\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__17182\,
            I => \N__17173\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__17179\,
            I => \c0.data_in_field_99\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__17176\,
            I => \c0.data_in_field_99\
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__17173\,
            I => \c0.data_in_field_99\
        );

    \I__2675\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17163\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__17163\,
            I => \N__17159\
        );

    \I__2673\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17156\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__17159\,
            I => \N__17150\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__17156\,
            I => \N__17147\
        );

    \I__2670\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17140\
        );

    \I__2669\ : InMux
    port map (
            O => \N__17154\,
            I => \N__17140\
        );

    \I__2668\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17140\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__17150\,
            I => \c0.data_in_field_65\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__17147\,
            I => \c0.data_in_field_65\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__17140\,
            I => \c0.data_in_field_65\
        );

    \I__2664\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17130\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__17130\,
            I => \N__17127\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__17127\,
            I => \N__17121\
        );

    \I__2661\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17118\
        );

    \I__2660\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17113\
        );

    \I__2659\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17113\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__17121\,
            I => \c0.data_in_field_129\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__17118\,
            I => \c0.data_in_field_129\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__17113\,
            I => \c0.data_in_field_129\
        );

    \I__2655\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17103\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__17103\,
            I => \N__17100\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__17100\,
            I => \N__17097\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__17097\,
            I => \c0.n5569\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__17094\,
            I => \c0.n5569_cascade_\
        );

    \I__2650\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17088\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__17088\,
            I => \N__17082\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__17087\,
            I => \N__17079\
        );

    \I__2647\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17076\
        );

    \I__2646\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17073\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__17082\,
            I => \N__17070\
        );

    \I__2644\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17067\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__17076\,
            I => \c0.data_in_field_114\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__17073\,
            I => \c0.data_in_field_114\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__17070\,
            I => \c0.data_in_field_114\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__17067\,
            I => \c0.data_in_field_114\
        );

    \I__2639\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17055\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__17055\,
            I => \N__17052\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__17052\,
            I => \N__17049\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__17049\,
            I => \c0.n20_adj_1882\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__17046\,
            I => \c0.n2062_cascade_\
        );

    \I__2634\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17040\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17037\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__17037\,
            I => \N__17034\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__17034\,
            I => \c0.n44\
        );

    \I__2630\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17028\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__17028\,
            I => \N__17023\
        );

    \I__2628\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17020\
        );

    \I__2627\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17017\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__17023\,
            I => \N__17014\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__17020\,
            I => \N__17011\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__17017\,
            I => \N__17007\
        );

    \I__2623\ : Span4Mux_s2_h
    port map (
            O => \N__17014\,
            I => \N__17002\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__17011\,
            I => \N__17002\
        );

    \I__2621\ : InMux
    port map (
            O => \N__17010\,
            I => \N__16999\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__17007\,
            I => \c0.data_in_field_134\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__17002\,
            I => \c0.data_in_field_134\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__16999\,
            I => \c0.data_in_field_134\
        );

    \I__2617\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16989\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16986\
        );

    \I__2615\ : Span4Mux_s3_h
    port map (
            O => \N__16986\,
            I => \N__16983\
        );

    \I__2614\ : Span4Mux_v
    port map (
            O => \N__16983\,
            I => \N__16979\
        );

    \I__2613\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16976\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__16979\,
            I => \c0.n5503\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__16976\,
            I => \c0.n5503\
        );

    \I__2610\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16968\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__16968\,
            I => \N__16964\
        );

    \I__2608\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16961\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__16964\,
            I => \N__16958\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__16961\,
            I => \N__16955\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__16958\,
            I => \c0.n2095\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__16955\,
            I => \c0.n2095\
        );

    \I__2603\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16947\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__16947\,
            I => \c0.n16_adj_1871\
        );

    \I__2601\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16940\
        );

    \I__2600\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16937\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__16940\,
            I => \N__16934\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__16937\,
            I => \N__16930\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__16934\,
            I => \N__16927\
        );

    \I__2596\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16924\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__16930\,
            I => \N__16921\
        );

    \I__2594\ : Span4Mux_s2_h
    port map (
            O => \N__16927\,
            I => \N__16918\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__16924\,
            I => data_in_11_3
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__16921\,
            I => data_in_11_3
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__16918\,
            I => data_in_11_3
        );

    \I__2590\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16908\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__16908\,
            I => \c0.n2021\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16901\
        );

    \I__2587\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16898\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__16901\,
            I => \N__16894\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__16898\,
            I => \N__16891\
        );

    \I__2584\ : InMux
    port map (
            O => \N__16897\,
            I => \N__16887\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__16894\,
            I => \N__16882\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__16891\,
            I => \N__16882\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16890\,
            I => \N__16879\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__16887\,
            I => \c0.data_in_field_10\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__16882\,
            I => \c0.data_in_field_10\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16879\,
            I => \c0.data_in_field_10\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__16872\,
            I => \c0.n2021_cascade_\
        );

    \I__2576\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16864\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16861\
        );

    \I__2574\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16857\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__16864\,
            I => \N__16854\
        );

    \I__2572\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16851\
        );

    \I__2571\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16848\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__16857\,
            I => \c0.data_in_field_41\
        );

    \I__2569\ : Odrv12
    port map (
            O => \N__16854\,
            I => \c0.data_in_field_41\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__16851\,
            I => \c0.data_in_field_41\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16848\,
            I => \c0.data_in_field_41\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__16839\,
            I => \c0.n2074_cascade_\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16830\
        );

    \I__2564\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16830\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__16830\,
            I => \c0.n2000\
        );

    \I__2562\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16823\
        );

    \I__2561\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16820\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16817\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16814\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__16817\,
            I => \N__16809\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__16814\,
            I => \N__16806\
        );

    \I__2556\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16801\
        );

    \I__2555\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16801\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__16809\,
            I => \c0.data_in_field_26\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__16806\,
            I => \c0.data_in_field_26\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__16801\,
            I => \c0.data_in_field_26\
        );

    \I__2551\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16791\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__2549\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16782\
        );

    \I__2548\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16779\
        );

    \I__2547\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16776\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__16785\,
            I => \N__16771\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16771\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__16779\,
            I => \N__16768\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__16776\,
            I => \N__16763\
        );

    \I__2542\ : Span4Mux_h
    port map (
            O => \N__16771\,
            I => \N__16760\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__16768\,
            I => \N__16757\
        );

    \I__2540\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16752\
        );

    \I__2539\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16752\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__16763\,
            I => \c0.data_in_field_64\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__16760\,
            I => \c0.data_in_field_64\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__16757\,
            I => \c0.data_in_field_64\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__16752\,
            I => \c0.data_in_field_64\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__16743\,
            I => \N__16740\
        );

    \I__2533\ : InMux
    port map (
            O => \N__16740\,
            I => \N__16737\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__16737\,
            I => \N__16733\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16730\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__16733\,
            I => \N__16726\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16730\,
            I => \N__16723\
        );

    \I__2528\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16720\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__16726\,
            I => data_in_8_2
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__16723\,
            I => data_in_8_2
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__16720\,
            I => data_in_8_2
        );

    \I__2524\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16709\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16709\,
            I => \N__16703\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16700\
        );

    \I__2520\ : Span4Mux_v
    port map (
            O => \N__16703\,
            I => \N__16695\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__16700\,
            I => \N__16695\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__16695\,
            I => \N__16691\
        );

    \I__2517\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16688\
        );

    \I__2516\ : Sp12to4
    port map (
            O => \N__16691\,
            I => \N__16685\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__16688\,
            I => data_in_5_3
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__16685\,
            I => data_in_5_3
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__16680\,
            I => \N__16677\
        );

    \I__2512\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16674\,
            I => \N__16671\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__16668\,
            I => \c0.n6183\
        );

    \I__2508\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16662\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__16662\,
            I => \c0.n20_adj_1958\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__16659\,
            I => \c0.n31_adj_1896_cascade_\
        );

    \I__2505\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16653\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__16653\,
            I => \c0.n41\
        );

    \I__2503\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16647\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__16647\,
            I => \N__16642\
        );

    \I__2501\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16638\
        );

    \I__2500\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16635\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__16642\,
            I => \N__16632\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16629\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__16638\,
            I => \N__16626\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__16635\,
            I => \c0.data_in_field_6\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__16632\,
            I => \c0.data_in_field_6\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16629\,
            I => \c0.data_in_field_6\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__16626\,
            I => \c0.data_in_field_6\
        );

    \I__2492\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16614\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__16614\,
            I => \c0.n10_adj_1915\
        );

    \I__2490\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16608\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__16608\,
            I => \N__16605\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__16605\,
            I => \c0.n1913\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__16602\,
            I => \N__16599\
        );

    \I__2486\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16595\
        );

    \I__2485\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16591\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__16595\,
            I => \N__16588\
        );

    \I__2483\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16584\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__16591\,
            I => \N__16581\
        );

    \I__2481\ : Span4Mux_h
    port map (
            O => \N__16588\,
            I => \N__16578\
        );

    \I__2480\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16575\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__16584\,
            I => \c0.data_in_field_7\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__16581\,
            I => \c0.data_in_field_7\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__16578\,
            I => \c0.data_in_field_7\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__16575\,
            I => \c0.data_in_field_7\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__16566\,
            I => \N__16562\
        );

    \I__2474\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16558\
        );

    \I__2473\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16555\
        );

    \I__2472\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16552\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__16558\,
            I => data_in_0_1
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__16555\,
            I => data_in_0_1
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__16552\,
            I => data_in_0_1
        );

    \I__2468\ : InMux
    port map (
            O => \N__16545\,
            I => \N__16542\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__2466\ : Sp12to4
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__16536\,
            I => \c0.n2104\
        );

    \I__2464\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16530\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__16530\,
            I => \c0.n1835\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__16527\,
            I => \c0.n2104_cascade_\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__16524\,
            I => \N__16521\
        );

    \I__2460\ : InMux
    port map (
            O => \N__16521\,
            I => \N__16518\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__16518\,
            I => \N__16515\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__16515\,
            I => \N__16512\
        );

    \I__2457\ : Span4Mux_s2_h
    port map (
            O => \N__16512\,
            I => \N__16507\
        );

    \I__2456\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16502\
        );

    \I__2455\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16502\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__16507\,
            I => data_in_8_1
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__16502\,
            I => data_in_8_1
        );

    \I__2452\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16491\
        );

    \I__2450\ : Span4Mux_h
    port map (
            O => \N__16491\,
            I => \N__16485\
        );

    \I__2449\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16478\
        );

    \I__2448\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16478\
        );

    \I__2447\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16478\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__16485\,
            I => data_in_1_3
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__16478\,
            I => data_in_1_3
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__16473\,
            I => \N__16470\
        );

    \I__2443\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16466\
        );

    \I__2442\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16463\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16459\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16456\
        );

    \I__2439\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16453\
        );

    \I__2438\ : Odrv12
    port map (
            O => \N__16459\,
            I => data_in_6_3
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__16456\,
            I => data_in_6_3
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__16453\,
            I => data_in_6_3
        );

    \I__2435\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16439\
        );

    \I__2434\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16439\
        );

    \I__2433\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16436\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__16439\,
            I => data_in_12_3
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__16436\,
            I => data_in_12_3
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__16431\,
            I => \N__16427\
        );

    \I__2429\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16423\
        );

    \I__2428\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16420\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16413\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16410\
        );

    \I__2424\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16407\
        );

    \I__2423\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16404\
        );

    \I__2422\ : Span4Mux_s1_h
    port map (
            O => \N__16413\,
            I => \N__16399\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__16410\,
            I => \N__16399\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__16407\,
            I => data_in_2_7
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__16404\,
            I => data_in_2_7
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__16399\,
            I => data_in_2_7
        );

    \I__2417\ : InMux
    port map (
            O => \N__16392\,
            I => \N__16388\
        );

    \I__2416\ : InMux
    port map (
            O => \N__16391\,
            I => \N__16385\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16382\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__16385\,
            I => \N__16378\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__16382\,
            I => \N__16375\
        );

    \I__2412\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16372\
        );

    \I__2411\ : Span4Mux_h
    port map (
            O => \N__16378\,
            I => \N__16368\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__16375\,
            I => \N__16363\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16363\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16358\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__16368\,
            I => \N__16355\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__16363\,
            I => \N__16352\
        );

    \I__2405\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16349\
        );

    \I__2404\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16346\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__16358\,
            I => \c0.data_in_field_131\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__16355\,
            I => \c0.data_in_field_131\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__16352\,
            I => \c0.data_in_field_131\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__16349\,
            I => \c0.data_in_field_131\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__16346\,
            I => \c0.data_in_field_131\
        );

    \I__2398\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16332\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__16332\,
            I => \N__16326\
        );

    \I__2396\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16323\
        );

    \I__2395\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16318\
        );

    \I__2394\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16318\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__16326\,
            I => data_in_1_1
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__16323\,
            I => data_in_1_1
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__16318\,
            I => data_in_1_1
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__16311\,
            I => \c0.rx.n6294_cascade_\
        );

    \I__2389\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16298\
        );

    \I__2388\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16298\
        );

    \I__2387\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16298\
        );

    \I__2386\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16290\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__16298\,
            I => \N__16287\
        );

    \I__2384\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16277\
        );

    \I__2383\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16277\
        );

    \I__2382\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16277\
        );

    \I__2381\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16277\
        );

    \I__2380\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16274\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__16290\,
            I => \N__16269\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__16287\,
            I => \N__16269\
        );

    \I__2377\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16266\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__16277\,
            I => \N__16263\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__16274\,
            I => \N__16260\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__16269\,
            I => \r_SM_Main_2_adj_1989\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__16266\,
            I => \r_SM_Main_2_adj_1989\
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__16263\,
            I => \r_SM_Main_2_adj_1989\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__16260\,
            I => \r_SM_Main_2_adj_1989\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__16251\,
            I => \c0.rx.n75_cascade_\
        );

    \I__2369\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16245\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__2367\ : Odrv12
    port map (
            O => \N__16242\,
            I => \c0.rx.n5815\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__16239\,
            I => \n4_adj_1980_cascade_\
        );

    \I__2365\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__2364\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16230\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__16230\,
            I => rx_data_4
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__16227\,
            I => \n2198_cascade_\
        );

    \I__2361\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16219\
        );

    \I__2360\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16216\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \N__16213\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__16219\,
            I => \N__16203\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__16216\,
            I => \N__16203\
        );

    \I__2356\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16194\
        );

    \I__2355\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16194\
        );

    \I__2354\ : InMux
    port map (
            O => \N__16211\,
            I => \N__16194\
        );

    \I__2353\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16194\
        );

    \I__2352\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16189\
        );

    \I__2351\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16189\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__16203\,
            I => \N__16184\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16184\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__16189\,
            I => \c0.rx.n359\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__16184\,
            I => \c0.rx.n359\
        );

    \I__2346\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16176\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__16176\,
            I => \c0.rx.n5859\
        );

    \I__2344\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16168\
        );

    \I__2343\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16165\
        );

    \I__2342\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16162\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__16168\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16165\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__16162\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__2338\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16152\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16149\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__16149\,
            I => \c0.rx.n5823\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__16146\,
            I => \N__16142\
        );

    \I__2334\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16139\
        );

    \I__2333\ : InMux
    port map (
            O => \N__16142\,
            I => \N__16135\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16132\
        );

    \I__2331\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16128\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16125\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__16132\,
            I => \N__16122\
        );

    \I__2328\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16119\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__16128\,
            I => data_in_18_6
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__16125\,
            I => data_in_18_6
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__16122\,
            I => data_in_18_6
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__16119\,
            I => data_in_18_6
        );

    \I__2323\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16106\
        );

    \I__2322\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16103\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__16106\,
            I => \N__16100\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__16103\,
            I => \c0.data_in_frame_18_6\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__16100\,
            I => \c0.data_in_frame_18_6\
        );

    \I__2318\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16091\
        );

    \I__2317\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16088\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__16091\,
            I => \N__16085\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__16088\,
            I => \c0.data_in_frame_18_7\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__16085\,
            I => \c0.data_in_frame_18_7\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__16080\,
            I => \N__16076\
        );

    \I__2312\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16073\
        );

    \I__2311\ : InMux
    port map (
            O => \N__16076\,
            I => \N__16070\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__16073\,
            I => \N__16067\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__16070\,
            I => \N__16063\
        );

    \I__2308\ : Span12Mux_v
    port map (
            O => \N__16067\,
            I => \N__16060\
        );

    \I__2307\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16057\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__16063\,
            I => data_in_7_1
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__16060\,
            I => data_in_7_1
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__16057\,
            I => data_in_7_1
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__16050\,
            I => \n1764_cascade_\
        );

    \I__2302\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16044\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__16044\,
            I => \N__16040\
        );

    \I__2300\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16037\
        );

    \I__2299\ : Odrv4
    port map (
            O => \N__16040\,
            I => rx_data_5
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__16037\,
            I => rx_data_5
        );

    \I__2297\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16029\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__16029\,
            I => \N__16025\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16022\
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__16025\,
            I => rx_data_6
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__16022\,
            I => rx_data_6
        );

    \I__2292\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16014\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__16014\,
            I => \c0.rx.n5822\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16011\,
            I => \N__16006\
        );

    \I__2289\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16003\
        );

    \I__2288\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16000\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__15997\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__16003\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__16000\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__15997\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__2283\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15987\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__15987\,
            I => n4_adj_1980
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__15984\,
            I => \N__15978\
        );

    \I__2280\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15975\
        );

    \I__2279\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15968\
        );

    \I__2278\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15968\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15968\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__15975\,
            I => data_in_19_6
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__15968\,
            I => data_in_19_6
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__15963\,
            I => \N__15959\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15956\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15953\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__15956\,
            I => \N__15950\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15953\,
            I => \c0.data_in_frame_19_0\
        );

    \I__2269\ : Odrv12
    port map (
            O => \N__15950\,
            I => \c0.data_in_frame_19_0\
        );

    \I__2268\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15940\
        );

    \I__2267\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15935\
        );

    \I__2266\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15935\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__15940\,
            I => \c0.data_in_field_17\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__15935\,
            I => \c0.data_in_field_17\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__15930\,
            I => \c0.n6093_cascade_\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15924\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15924\,
            I => \N__15921\
        );

    \I__2260\ : Span4Mux_h
    port map (
            O => \N__15921\,
            I => \N__15918\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__15918\,
            I => \c0.n5767\
        );

    \I__2258\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15911\
        );

    \I__2257\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15908\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__15911\,
            I => \N__15902\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__15908\,
            I => \N__15902\
        );

    \I__2254\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15899\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__15902\,
            I => data_in_16_2
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__15899\,
            I => data_in_16_2
        );

    \I__2251\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15891\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__15891\,
            I => \N__15888\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__15888\,
            I => \c0.n5512\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__15885\,
            I => \c0.n5512_cascade_\
        );

    \I__2247\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15879\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__15879\,
            I => \c0.n22\
        );

    \I__2245\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15873\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__15873\,
            I => \N__15869\
        );

    \I__2243\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15866\
        );

    \I__2242\ : Odrv12
    port map (
            O => \N__15869\,
            I => \c0.n2155\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__15866\,
            I => \c0.n2155\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__15861\,
            I => \c0.n2155_cascade_\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__15858\,
            I => \N__15855\
        );

    \I__2238\ : InMux
    port map (
            O => \N__15855\,
            I => \N__15852\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15849\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__15849\,
            I => \N__15846\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__15846\,
            I => \N__15843\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__15843\,
            I => \c0.n43\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15837\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__15837\,
            I => \N__15834\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__15834\,
            I => \N__15830\
        );

    \I__2230\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15827\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__15830\,
            I => \c0.n2026\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__15827\,
            I => \c0.n2026\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__15822\,
            I => \N__15819\
        );

    \I__2226\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15816\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__15816\,
            I => \N__15812\
        );

    \I__2224\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15809\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__15812\,
            I => \N__15805\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__15809\,
            I => \N__15802\
        );

    \I__2221\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15799\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__15805\,
            I => data_in_16_1
        );

    \I__2219\ : Odrv12
    port map (
            O => \N__15802\,
            I => data_in_16_1
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__15799\,
            I => data_in_16_1
        );

    \I__2217\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15786\
        );

    \I__2216\ : InMux
    port map (
            O => \N__15791\,
            I => \N__15786\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__15783\,
            I => \N__15780\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__15780\,
            I => \c0.n2080\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15774\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__15774\,
            I => \N__15770\
        );

    \I__2210\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15767\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__15770\,
            I => \c0.n2012\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__15767\,
            I => \c0.n2012\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__15762\,
            I => \N__15759\
        );

    \I__2206\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15755\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15752\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__15755\,
            I => \c0.n1973\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__15752\,
            I => \c0.n1973\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15743\
        );

    \I__2201\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15740\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__15743\,
            I => \N__15737\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__15740\,
            I => \N__15730\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__15737\,
            I => \N__15730\
        );

    \I__2197\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15727\
        );

    \I__2196\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15724\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__15730\,
            I => \N__15719\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__15727\,
            I => \N__15719\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__15724\,
            I => data_in_19_3
        );

    \I__2192\ : Odrv12
    port map (
            O => \N__15719\,
            I => data_in_19_3
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__15714\,
            I => \c0.n18_adj_1959_cascade_\
        );

    \I__2190\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__15708\,
            I => \N__15705\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__15705\,
            I => \c0.n16\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__15702\,
            I => \c0.n20_adj_1870_cascade_\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15696\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15696\,
            I => \c0.n5577\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__15693\,
            I => \c0.n2101_cascade_\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__15690\,
            I => \c0.n6_adj_1917_cascade_\
        );

    \I__2182\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15684\,
            I => \N__15680\
        );

    \I__2180\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15677\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__15680\,
            I => \N__15672\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__15677\,
            I => \N__15669\
        );

    \I__2177\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15664\
        );

    \I__2176\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15664\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__15672\,
            I => \c0.data_in_field_68\
        );

    \I__2174\ : Odrv12
    port map (
            O => \N__15669\,
            I => \c0.data_in_field_68\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__15664\,
            I => \c0.data_in_field_68\
        );

    \I__2172\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15654\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__15654\,
            I => \N__15650\
        );

    \I__2170\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15647\
        );

    \I__2169\ : Span4Mux_h
    port map (
            O => \N__15650\,
            I => \N__15644\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__15647\,
            I => \c0.n5557\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__15644\,
            I => \c0.n5557\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__15639\,
            I => \c0.n17_cascade_\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__15633\,
            I => \c0.n5574\
        );

    \I__2163\ : InMux
    port map (
            O => \N__15630\,
            I => \N__15627\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__15627\,
            I => \N__15624\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__15624\,
            I => \N__15620\
        );

    \I__2160\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15617\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__15620\,
            I => \c0.n5572\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__15617\,
            I => \c0.n5572\
        );

    \I__2157\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15608\
        );

    \I__2156\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15605\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__15608\,
            I => \N__15602\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__15605\,
            I => \N__15599\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__15602\,
            I => \N__15595\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__15599\,
            I => \N__15592\
        );

    \I__2151\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15589\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__15595\,
            I => data_in_8_7
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__15592\,
            I => data_in_8_7
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__15589\,
            I => data_in_8_7
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__15582\,
            I => \N__15579\
        );

    \I__2146\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15576\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__15576\,
            I => \N__15572\
        );

    \I__2144\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15569\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__15572\,
            I => \N__15565\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15562\
        );

    \I__2141\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15559\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__15565\,
            I => data_in_17_1
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__15562\,
            I => data_in_17_1
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__15559\,
            I => data_in_17_1
        );

    \I__2137\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15548\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__15551\,
            I => \N__15545\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__15548\,
            I => \N__15541\
        );

    \I__2134\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15536\
        );

    \I__2133\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15533\
        );

    \I__2132\ : Span12Mux_v
    port map (
            O => \N__15541\,
            I => \N__15530\
        );

    \I__2131\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15525\
        );

    \I__2130\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15525\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__15536\,
            I => \c0.data_in_field_138\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__15533\,
            I => \c0.data_in_field_138\
        );

    \I__2127\ : Odrv12
    port map (
            O => \N__15530\,
            I => \c0.data_in_field_138\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__15525\,
            I => \c0.data_in_field_138\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15513\
        );

    \I__2124\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15509\
        );

    \I__2123\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15505\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__15509\,
            I => \N__15502\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__15508\,
            I => \N__15499\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__15505\,
            I => \N__15494\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__15502\,
            I => \N__15494\
        );

    \I__2118\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15489\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__15494\,
            I => \N__15486\
        );

    \I__2116\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15481\
        );

    \I__2115\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15481\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__15489\,
            I => \c0.data_in_field_130\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__15486\,
            I => \c0.data_in_field_130\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__15481\,
            I => \c0.data_in_field_130\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__2110\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__15468\,
            I => \N__15465\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__15465\,
            I => \N__15462\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__15462\,
            I => \c0.n6213\
        );

    \I__2106\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15454\
        );

    \I__2105\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15451\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__15457\,
            I => \N__15448\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__15454\,
            I => \N__15445\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__15451\,
            I => \N__15442\
        );

    \I__2101\ : InMux
    port map (
            O => \N__15448\,
            I => \N__15437\
        );

    \I__2100\ : Span4Mux_s3_h
    port map (
            O => \N__15445\,
            I => \N__15434\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__15442\,
            I => \N__15431\
        );

    \I__2098\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15426\
        );

    \I__2097\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15426\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__15437\,
            I => \c0.data_in_field_73\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__15434\,
            I => \c0.data_in_field_73\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__15431\,
            I => \c0.data_in_field_73\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__15426\,
            I => \c0.data_in_field_73\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__15417\,
            I => \c0.n14_adj_1957_cascade_\
        );

    \I__2091\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15406\
        );

    \I__2090\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15406\
        );

    \I__2089\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15401\
        );

    \I__2088\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15401\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__15406\,
            I => \c0.data_in_field_53\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__15401\,
            I => \c0.data_in_field_53\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__15396\,
            I => \c0.n22_adj_1903_cascade_\
        );

    \I__2084\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15390\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__15390\,
            I => \c0.n18_adj_1904\
        );

    \I__2082\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15384\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__15384\,
            I => \c0.n20_adj_1905\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__15381\,
            I => \c0.n5589_cascade_\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__15378\,
            I => \N__15375\
        );

    \I__2078\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15372\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__15372\,
            I => \N__15369\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__15369\,
            I => \N__15366\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__15366\,
            I => \N__15363\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__15363\,
            I => \c0.n29\
        );

    \I__2073\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15354\
        );

    \I__2072\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15354\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__15354\,
            I => \c0.n5458\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \N__15348\
        );

    \I__2069\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15345\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__15345\,
            I => \N__15342\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__15342\,
            I => \N__15338\
        );

    \I__2066\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15335\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__15338\,
            I => \c0.n1994\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__15335\,
            I => \c0.n1994\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__15330\,
            I => \c0.n6009_cascade_\
        );

    \I__2062\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__15321\,
            I => \N__15318\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__15318\,
            I => \c0.n6012\
        );

    \I__2058\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15310\
        );

    \I__2057\ : InMux
    port map (
            O => \N__15314\,
            I => \N__15305\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15305\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__15310\,
            I => \c0.data_in_field_15\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__15305\,
            I => \c0.data_in_field_15\
        );

    \I__2053\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__15297\,
            I => \N__15294\
        );

    \I__2051\ : Span4Mux_s2_h
    port map (
            O => \N__15294\,
            I => \N__15291\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__15291\,
            I => \N__15286\
        );

    \I__2049\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15281\
        );

    \I__2048\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15281\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__15286\,
            I => \c0.data_in_field_8\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__15281\,
            I => \c0.data_in_field_8\
        );

    \I__2045\ : InMux
    port map (
            O => \N__15276\,
            I => \N__15273\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__15273\,
            I => \c0.n2039\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \c0.n2039_cascade_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15262\
        );

    \I__2041\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15258\
        );

    \I__2040\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15255\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__15262\,
            I => \N__15252\
        );

    \I__2038\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15249\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__15258\,
            I => \c0.data_in_field_23\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__15255\,
            I => \c0.data_in_field_23\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__15252\,
            I => \c0.data_in_field_23\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__15249\,
            I => \c0.data_in_field_23\
        );

    \I__2033\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15237\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__15237\,
            I => \c0.rx.n5857\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__15234\,
            I => \N__15230\
        );

    \I__2030\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15226\
        );

    \I__2029\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15223\
        );

    \I__2028\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15220\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__15226\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__15223\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__15220\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__2024\ : IoInMux
    port map (
            O => \N__15213\,
            I => \N__15210\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__15210\,
            I => tx_enable
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__15207\,
            I => \N__15204\
        );

    \I__2021\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15201\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__15201\,
            I => \N__15197\
        );

    \I__2019\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15194\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__15197\,
            I => \N__15190\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__15194\,
            I => \N__15187\
        );

    \I__2016\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15184\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__15190\,
            I => data_in_16_3
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__15187\,
            I => data_in_16_3
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__15184\,
            I => data_in_16_3
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__15177\,
            I => \N__15174\
        );

    \I__2011\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15168\
        );

    \I__2010\ : InMux
    port map (
            O => \N__15173\,
            I => \N__15168\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__15168\,
            I => rx_data_3
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__15165\,
            I => \N__15162\
        );

    \I__2007\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15158\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15161\,
            I => \N__15155\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__15158\,
            I => \N__15152\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__15155\,
            I => \N__15149\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__15152\,
            I => \N__15144\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__15149\,
            I => \N__15141\
        );

    \I__2001\ : InMux
    port map (
            O => \N__15148\,
            I => \N__15138\
        );

    \I__2000\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15135\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__15144\,
            I => \N__15132\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__15141\,
            I => data_in_18_1
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__15138\,
            I => data_in_18_1
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__15135\,
            I => data_in_18_1
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__15132\,
            I => data_in_18_1
        );

    \I__1994\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15111\
        );

    \I__1993\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15111\
        );

    \I__1992\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15111\
        );

    \I__1991\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15111\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__15111\,
            I => \N__15104\
        );

    \I__1989\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15095\
        );

    \I__1988\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15095\
        );

    \I__1987\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15095\
        );

    \I__1986\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15095\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__15104\,
            I => \c0.rx.n36\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__15095\,
            I => \c0.rx.n36\
        );

    \I__1983\ : InMux
    port map (
            O => \N__15090\,
            I => \c0.rx.n4778\
        );

    \I__1982\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15084\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__15084\,
            I => \c0.rx.n5361\
        );

    \I__1980\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15078\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__15078\,
            I => \c0.rx.n5858\
        );

    \I__1978\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15072\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__15072\,
            I => \c0.rx.n5854\
        );

    \I__1976\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15064\
        );

    \I__1975\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15061\
        );

    \I__1974\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15058\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__15064\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__15061\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__15058\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__1970\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15046\
        );

    \I__1969\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15041\
        );

    \I__1968\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15041\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__15046\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__15041\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__1965\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15031\
        );

    \I__1964\ : InMux
    port map (
            O => \N__15035\,
            I => \N__15028\
        );

    \I__1963\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15025\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__15031\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__15028\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__15025\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__15018\,
            I => \c0.rx.n8_cascade_\
        );

    \I__1958\ : InMux
    port map (
            O => \N__15015\,
            I => \N__15003\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15014\,
            I => \N__15003\
        );

    \I__1956\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15003\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15012\,
            I => \N__15003\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__15003\,
            I => \c0.rx.n1724\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__15000\,
            I => \c0.rx.n1724_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14988\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14985\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14995\,
            I => \N__14982\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14975\
        );

    \I__1948\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14975\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14975\
        );

    \I__1946\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14972\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__14988\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__14985\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__14982\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__14975\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14972\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__1940\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14958\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__14958\,
            I => \c0.rx.n5855\
        );

    \I__1938\ : InMux
    port map (
            O => \N__14955\,
            I => \N__14946\
        );

    \I__1937\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14943\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14938\
        );

    \I__1935\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14938\
        );

    \I__1934\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14931\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14931\
        );

    \I__1932\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14931\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__14946\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__14943\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__14938\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__14931\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__14922\,
            I => \N__14918\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14915\
        );

    \I__1925\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14911\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14908\
        );

    \I__1923\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14905\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__14911\,
            I => \c0.data_in_field_104\
        );

    \I__1921\ : Odrv12
    port map (
            O => \N__14908\,
            I => \c0.data_in_field_104\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__14905\,
            I => \c0.data_in_field_104\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__14898\,
            I => \c0.n6021_cascade_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14892\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14889\
        );

    \I__1916\ : Span4Mux_s3_h
    port map (
            O => \N__14889\,
            I => \N__14886\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__14886\,
            I => \c0.n5797\
        );

    \I__1914\ : InMux
    port map (
            O => \N__14883\,
            I => \bfn_4_27_0_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14877\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__14877\,
            I => \c0.rx.n5860\
        );

    \I__1911\ : InMux
    port map (
            O => \N__14874\,
            I => \c0.rx.n4772\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14871\,
            I => \c0.rx.n4773\
        );

    \I__1909\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14865\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__14865\,
            I => \c0.rx.n5856\
        );

    \I__1907\ : InMux
    port map (
            O => \N__14862\,
            I => \c0.rx.n4774\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14859\,
            I => \c0.rx.n4775\
        );

    \I__1905\ : InMux
    port map (
            O => \N__14856\,
            I => \c0.rx.n4776\
        );

    \I__1904\ : InMux
    port map (
            O => \N__14853\,
            I => \c0.rx.n4777\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__14850\,
            I => \c0.n6147_cascade_\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14844\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__14844\,
            I => \N__14841\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__14841\,
            I => \N__14838\
        );

    \I__1899\ : IoSpan4Mux
    port map (
            O => \N__14838\,
            I => \N__14835\
        );

    \I__1898\ : Span4Mux_s1_h
    port map (
            O => \N__14835\,
            I => \N__14832\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__14832\,
            I => \c0.n6150\
        );

    \I__1896\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14825\
        );

    \I__1895\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14822\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14819\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__14822\,
            I => \c0.data_in_frame_19_4\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__14819\,
            I => \c0.data_in_frame_19_4\
        );

    \I__1891\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14811\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__14808\,
            I => \N__14803\
        );

    \I__1888\ : InMux
    port map (
            O => \N__14807\,
            I => \N__14798\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14798\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__14803\,
            I => \c0.data_in_field_14\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14798\,
            I => \c0.data_in_field_14\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__14793\,
            I => \c0.n6255_cascade_\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__14790\,
            I => \N__14787\
        );

    \I__1882\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14784\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__14784\,
            I => \c0.n5692\
        );

    \I__1880\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14778\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__14778\,
            I => \N__14775\
        );

    \I__1878\ : Span4Mux_v
    port map (
            O => \N__14775\,
            I => \N__14770\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14765\
        );

    \I__1876\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14765\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__14770\,
            I => \c0.data_in_field_119\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__14765\,
            I => \c0.data_in_field_119\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__14760\,
            I => \c0.n6273_cascade_\
        );

    \I__1872\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14754\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__14754\,
            I => \N__14750\
        );

    \I__1870\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14746\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__14750\,
            I => \N__14743\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14740\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__14746\,
            I => \c0.data_in_field_111\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__14743\,
            I => \c0.data_in_field_111\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__14740\,
            I => \c0.data_in_field_111\
        );

    \I__1864\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14730\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__14730\,
            I => \c0.n5994\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__14727\,
            I => \c0.n5686_cascade_\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__14724\,
            I => \c0.n6261_cascade_\
        );

    \I__1860\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14718\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__14718\,
            I => \c0.n6264\
        );

    \I__1858\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14710\
        );

    \I__1857\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14707\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__14713\,
            I => \N__14704\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__14710\,
            I => \N__14701\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__14707\,
            I => \N__14698\
        );

    \I__1853\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14695\
        );

    \I__1852\ : Span4Mux_s3_h
    port map (
            O => \N__14701\,
            I => \N__14691\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__14698\,
            I => \N__14688\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14685\
        );

    \I__1849\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14682\
        );

    \I__1848\ : Sp12to4
    port map (
            O => \N__14691\,
            I => \N__14679\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__14688\,
            I => \N__14674\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__14685\,
            I => \N__14674\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__14682\,
            I => data_in_18_3
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__14679\,
            I => data_in_18_3
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__14674\,
            I => data_in_18_3
        );

    \I__1842\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14664\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__14664\,
            I => \N__14661\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__14661\,
            I => \c0.n5725\
        );

    \I__1839\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14655\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__14655\,
            I => \N__14652\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__14652\,
            I => \c0.n6165\
        );

    \I__1836\ : InMux
    port map (
            O => \N__14649\,
            I => \N__14646\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__14646\,
            I => \N__14643\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__14643\,
            I => \N__14640\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__14640\,
            I => \c0.n6168\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__14637\,
            I => \N__14634\
        );

    \I__1831\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14631\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__14631\,
            I => \c0.n20_adj_1878\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__1828\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14622\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__14622\,
            I => \N__14618\
        );

    \I__1826\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14615\
        );

    \I__1825\ : Span12Mux_s11_v
    port map (
            O => \N__14618\,
            I => \N__14611\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__14615\,
            I => \N__14608\
        );

    \I__1823\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14605\
        );

    \I__1822\ : Odrv12
    port map (
            O => \N__14611\,
            I => data_in_7_2
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__14608\,
            I => data_in_7_2
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__14605\,
            I => data_in_7_2
        );

    \I__1819\ : InMux
    port map (
            O => \N__14598\,
            I => \N__14595\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__14595\,
            I => \N__14591\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__14594\,
            I => \N__14587\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__14591\,
            I => \N__14583\
        );

    \I__1815\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14576\
        );

    \I__1814\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14576\
        );

    \I__1813\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14576\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__14583\,
            I => \c0.data_in_field_58\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__14576\,
            I => \c0.data_in_field_58\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__14571\,
            I => \N__14567\
        );

    \I__1809\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14564\
        );

    \I__1808\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14561\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__14564\,
            I => \c0.data_in_frame_19_6\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__14561\,
            I => \c0.data_in_frame_19_6\
        );

    \I__1805\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__14550\,
            I => \c0.n5578\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__14547\,
            I => \c0.n6177_cascade_\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__14544\,
            I => \c0.n5728_cascade_\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \c0.n16_adj_1873_cascade_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14535\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__14535\,
            I => \c0.n24\
        );

    \I__1797\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14526\
        );

    \I__1796\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14521\
        );

    \I__1795\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14521\
        );

    \I__1794\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14518\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__14526\,
            I => \c0.data_in_field_81\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__14521\,
            I => \c0.data_in_field_81\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__14518\,
            I => \c0.data_in_field_81\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__14511\,
            I => \N__14508\
        );

    \I__1789\ : InMux
    port map (
            O => \N__14508\,
            I => \N__14505\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14502\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__14502\,
            I => \N__14499\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__14499\,
            I => \c0.n5551\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__14496\,
            I => \c0.n5551_cascade_\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14490\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__14490\,
            I => \N__14487\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__14487\,
            I => \N__14483\
        );

    \I__1781\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14480\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__14483\,
            I => \c0.n1892\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__14480\,
            I => \c0.n1892\
        );

    \I__1778\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14472\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__14472\,
            I => \c0.n20\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__14469\,
            I => \c0.n19_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14461\
        );

    \I__1774\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14458\
        );

    \I__1773\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14455\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__14461\,
            I => data_in_10_3
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__14458\,
            I => data_in_10_3
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__14455\,
            I => data_in_10_3
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__14448\,
            I => \c0.n5412_cascade_\
        );

    \I__1768\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14442\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14439\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__14439\,
            I => \c0.n16_adj_1880\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__14436\,
            I => \c0.n22_adj_1881_cascade_\
        );

    \I__1764\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14430\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__14430\,
            I => \N__14427\
        );

    \I__1762\ : Span4Mux_s3_h
    port map (
            O => \N__14427\,
            I => \N__14424\
        );

    \I__1761\ : Sp12to4
    port map (
            O => \N__14424\,
            I => \N__14421\
        );

    \I__1760\ : Odrv12
    port map (
            O => \N__14421\,
            I => \c0.n24_adj_1884\
        );

    \I__1759\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14415\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__14415\,
            I => \N__14411\
        );

    \I__1757\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14406\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__14411\,
            I => \N__14403\
        );

    \I__1755\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14398\
        );

    \I__1754\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14398\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__14406\,
            I => \c0.data_in_field_11\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__14403\,
            I => \c0.data_in_field_11\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__14398\,
            I => \c0.data_in_field_11\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__14391\,
            I => \N__14387\
        );

    \I__1749\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14384\
        );

    \I__1748\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14380\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14377\
        );

    \I__1746\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14374\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__14380\,
            I => data_in_8_3
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__14377\,
            I => data_in_8_3
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__14374\,
            I => data_in_8_3
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__14367\,
            I => \N__14361\
        );

    \I__1741\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14358\
        );

    \I__1740\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14355\
        );

    \I__1739\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14352\
        );

    \I__1738\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14349\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__14358\,
            I => \c0.data_in_field_67\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__14355\,
            I => \c0.data_in_field_67\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__14352\,
            I => \c0.data_in_field_67\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__14349\,
            I => \c0.data_in_field_67\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__14340\,
            I => \c0.rx.n3589_cascade_\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__14337\,
            I => \c0.rx.n17_cascade_\
        );

    \I__1731\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14331\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__14331\,
            I => \c0.rx.n5817\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__14328\,
            I => \N__14325\
        );

    \I__1728\ : InMux
    port map (
            O => \N__14325\,
            I => \N__14322\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__14322\,
            I => \N__14317\
        );

    \I__1726\ : InMux
    port map (
            O => \N__14321\,
            I => \N__14314\
        );

    \I__1725\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14311\
        );

    \I__1724\ : Span4Mux_h
    port map (
            O => \N__14317\,
            I => \N__14308\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__14314\,
            I => data_in_15_3
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__14311\,
            I => data_in_15_3
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__14308\,
            I => data_in_15_3
        );

    \I__1720\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14298\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14294\
        );

    \I__1718\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14290\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__14294\,
            I => \N__14287\
        );

    \I__1716\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14284\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__14290\,
            I => \c0.data_in_field_59\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__14287\,
            I => \c0.data_in_field_59\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__14284\,
            I => \c0.data_in_field_59\
        );

    \I__1712\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14274\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__14274\,
            I => \N__14268\
        );

    \I__1710\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14263\
        );

    \I__1709\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14263\
        );

    \I__1708\ : InMux
    port map (
            O => \N__14271\,
            I => \N__14260\
        );

    \I__1707\ : Span4Mux_s3_h
    port map (
            O => \N__14268\,
            I => \N__14257\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14254\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__14260\,
            I => \c0.data_in_field_123\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__14257\,
            I => \c0.data_in_field_123\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__14254\,
            I => \c0.data_in_field_123\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__14247\,
            I => \N__14243\
        );

    \I__1701\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14239\
        );

    \I__1700\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14234\
        );

    \I__1699\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14234\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__14239\,
            I => data_in_7_3
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__14234\,
            I => data_in_7_3
        );

    \I__1696\ : InMux
    port map (
            O => \N__14229\,
            I => \c0.n4738\
        );

    \I__1695\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14222\
        );

    \I__1694\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14214\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__14222\,
            I => \N__14211\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \N__14208\
        );

    \I__1691\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14200\
        );

    \I__1690\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14200\
        );

    \I__1689\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14195\
        );

    \I__1688\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14195\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__14214\,
            I => \N__14190\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__14211\,
            I => \N__14190\
        );

    \I__1685\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14187\
        );

    \I__1684\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14182\
        );

    \I__1683\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14182\
        );

    \I__1682\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14179\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__14200\,
            I => \N__14174\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14174\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__14190\,
            I => \N__14171\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__14187\,
            I => \N__14168\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__14182\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__14179\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__14174\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__14171\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__14168\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__1672\ : CEMux
    port map (
            O => \N__14157\,
            I => \N__14154\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__14154\,
            I => \N__14151\
        );

    \I__1670\ : Odrv12
    port map (
            O => \N__14151\,
            I => \c0.n195\
        );

    \I__1669\ : SRMux
    port map (
            O => \N__14148\,
            I => \N__14145\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__14145\,
            I => \N__14142\
        );

    \I__1667\ : Span4Mux_h
    port map (
            O => \N__14142\,
            I => \N__14139\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__14139\,
            I => \c0.n2325\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__14136\,
            I => \N__14133\
        );

    \I__1664\ : InMux
    port map (
            O => \N__14133\,
            I => \N__14129\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \N__14120\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__14129\,
            I => \N__14116\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__14128\,
            I => \N__14108\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__14127\,
            I => \N__14105\
        );

    \I__1659\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14101\
        );

    \I__1658\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14092\
        );

    \I__1657\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14092\
        );

    \I__1656\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14092\
        );

    \I__1655\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14089\
        );

    \I__1654\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14086\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__14116\,
            I => \N__14083\
        );

    \I__1652\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14078\
        );

    \I__1651\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14078\
        );

    \I__1650\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14071\
        );

    \I__1649\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14071\
        );

    \I__1648\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14071\
        );

    \I__1647\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14064\
        );

    \I__1646\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14064\
        );

    \I__1645\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14064\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__14101\,
            I => \N__14061\
        );

    \I__1643\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14056\
        );

    \I__1642\ : InMux
    port map (
            O => \N__14099\,
            I => \N__14056\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__14092\,
            I => \N__14049\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__14089\,
            I => \N__14049\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__14086\,
            I => \N__14049\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__14083\,
            I => \N__14044\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14044\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__14071\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__14064\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__14061\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__14056\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__14049\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__14044\,
            I => \r_SM_Main_2_adj_1992\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14028\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__14028\,
            I => \c0.tx2.n14\
        );

    \I__1628\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14021\
        );

    \I__1627\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14018\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__14021\,
            I => \N__14013\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__14018\,
            I => \N__14008\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__14017\,
            I => \N__14003\
        );

    \I__1623\ : InMux
    port map (
            O => \N__14016\,
            I => \N__14000\
        );

    \I__1622\ : Span4Mux_s2_h
    port map (
            O => \N__14013\,
            I => \N__13997\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14012\,
            I => \N__13992\
        );

    \I__1620\ : InMux
    port map (
            O => \N__14011\,
            I => \N__13992\
        );

    \I__1619\ : Span4Mux_s2_h
    port map (
            O => \N__14008\,
            I => \N__13989\
        );

    \I__1618\ : InMux
    port map (
            O => \N__14007\,
            I => \N__13982\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13982\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13982\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__14000\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__13997\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13992\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__13989\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__13982\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__1610\ : CEMux
    port map (
            O => \N__13971\,
            I => \N__13968\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__13968\,
            I => \N__13965\
        );

    \I__1608\ : Span4Mux_s2_h
    port map (
            O => \N__13965\,
            I => \N__13960\
        );

    \I__1607\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13957\
        );

    \I__1606\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13954\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__13960\,
            I => n2208
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__13957\,
            I => n2208
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13954\,
            I => n2208
        );

    \I__1602\ : SRMux
    port map (
            O => \N__13947\,
            I => \N__13944\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__13944\,
            I => \N__13941\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__13941\,
            I => \N__13937\
        );

    \I__1599\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13934\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__13937\,
            I => n2339
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__13934\,
            I => n2339
        );

    \I__1596\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13922\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13922\
        );

    \I__1594\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13919\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13915\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__13919\,
            I => \N__13909\
        );

    \I__1591\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13906\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__13915\,
            I => \N__13903\
        );

    \I__1589\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13900\
        );

    \I__1588\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13895\
        );

    \I__1587\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13895\
        );

    \I__1586\ : Span4Mux_v
    port map (
            O => \N__13909\,
            I => \N__13890\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__13906\,
            I => \N__13890\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__13903\,
            I => \r_Bit_Index_0_adj_1995\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__13900\,
            I => \r_Bit_Index_0_adj_1995\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__13895\,
            I => \r_Bit_Index_0_adj_1995\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__13890\,
            I => \r_Bit_Index_0_adj_1995\
        );

    \I__1580\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13874\
        );

    \I__1579\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13871\
        );

    \I__1578\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13868\
        );

    \I__1577\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13863\
        );

    \I__1576\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13863\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__13874\,
            I => \c0.tx2.r_SM_Main_2_N_1767_1\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__13871\,
            I => \c0.tx2.r_SM_Main_2_N_1767_1\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__13868\,
            I => \c0.tx2.r_SM_Main_2_N_1767_1\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__13863\,
            I => \c0.tx2.r_SM_Main_2_N_1767_1\
        );

    \I__1571\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13851\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__13851\,
            I => \c0.tx2.n5847\
        );

    \I__1569\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13845\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__13845\,
            I => \c0.rx.n3589\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__13842\,
            I => \N__13839\
        );

    \I__1566\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13836\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__13836\,
            I => \N__13833\
        );

    \I__1564\ : Span4Mux_s2_h
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__13830\,
            I => \c0.n6081\
        );

    \I__1562\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__13824\,
            I => \N__13821\
        );

    \I__1560\ : Span4Mux_h
    port map (
            O => \N__13821\,
            I => \N__13818\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__13818\,
            I => \N__13815\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__13815\,
            I => \c0.n6084\
        );

    \I__1557\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13809\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__13809\,
            I => \c0.n5695\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__13806\,
            I => \c0.n6234_cascade_\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__13803\,
            I => \N__13799\
        );

    \I__1553\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13793\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13790\
        );

    \I__1551\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13784\
        );

    \I__1550\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13779\
        );

    \I__1549\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13779\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__13793\,
            I => \N__13774\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__13790\,
            I => \N__13774\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13767\
        );

    \I__1545\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13767\
        );

    \I__1544\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13767\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__13784\,
            I => \N__13761\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__13779\,
            I => \N__13761\
        );

    \I__1541\ : Span4Mux_h
    port map (
            O => \N__13774\,
            I => \N__13758\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__13767\,
            I => \N__13755\
        );

    \I__1539\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13752\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__13761\,
            I => \N__13749\
        );

    \I__1537\ : Sp12to4
    port map (
            O => \N__13758\,
            I => \N__13744\
        );

    \I__1536\ : Span12Mux_h
    port map (
            O => \N__13755\,
            I => \N__13744\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13752\,
            I => \c0.n1081\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__13749\,
            I => \c0.n1081\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__13744\,
            I => \c0.n1081\
        );

    \I__1532\ : CEMux
    port map (
            O => \N__13737\,
            I => \N__13733\
        );

    \I__1531\ : CEMux
    port map (
            O => \N__13736\,
            I => \N__13729\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13724\
        );

    \I__1529\ : CEMux
    port map (
            O => \N__13732\,
            I => \N__13721\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13718\
        );

    \I__1527\ : CEMux
    port map (
            O => \N__13728\,
            I => \N__13715\
        );

    \I__1526\ : CEMux
    port map (
            O => \N__13727\,
            I => \N__13712\
        );

    \I__1525\ : Span4Mux_h
    port map (
            O => \N__13724\,
            I => \N__13707\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13721\,
            I => \N__13707\
        );

    \I__1523\ : Span4Mux_s1_h
    port map (
            O => \N__13718\,
            I => \N__13702\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__13715\,
            I => \N__13702\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__13712\,
            I => \N__13699\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__13707\,
            I => \N__13696\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__13702\,
            I => \N__13693\
        );

    \I__1518\ : Sp12to4
    port map (
            O => \N__13699\,
            I => \N__13690\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__13696\,
            I => \N__13687\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__13693\,
            I => \c0.tx2.n1624\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__13690\,
            I => \c0.tx2.n1624\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__13687\,
            I => \c0.tx2.n1624\
        );

    \I__1513\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13677\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__13677\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__1511\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13671\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13671\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__13668\,
            I => \N__13665\
        );

    \I__1508\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13660\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__13664\,
            I => \N__13656\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13653\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13650\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__13659\,
            I => \N__13647\
        );

    \I__1503\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13641\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__13653\,
            I => \N__13638\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__13650\,
            I => \N__13635\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13647\,
            I => \N__13630\
        );

    \I__1499\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13630\
        );

    \I__1498\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13627\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13624\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__13641\,
            I => \N__13619\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__13638\,
            I => \N__13619\
        );

    \I__1494\ : Span4Mux_h
    port map (
            O => \N__13635\,
            I => \N__13616\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__13630\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__13627\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__13624\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__13619\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__13616\,
            I => \c0.tx2.r_Bit_Index_1\
        );

    \I__1488\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13602\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__13602\,
            I => \N__13599\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__13599\,
            I => \N__13596\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__13596\,
            I => \c0.tx2.n6003\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__13593\,
            I => \N__13588\
        );

    \I__1483\ : InMux
    port map (
            O => \N__13592\,
            I => \N__13583\
        );

    \I__1482\ : InMux
    port map (
            O => \N__13591\,
            I => \N__13583\
        );

    \I__1481\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13580\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13577\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13574\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__13577\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_909\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__13574\,
            I => \c0.FRAME_MATCHER_wait_for_transmission_N_909\
        );

    \I__1476\ : InMux
    port map (
            O => \N__13569\,
            I => \c0.n4735\
        );

    \I__1475\ : InMux
    port map (
            O => \N__13566\,
            I => \c0.n4736\
        );

    \I__1474\ : InMux
    port map (
            O => \N__13563\,
            I => \c0.n4737\
        );

    \I__1473\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13556\
        );

    \I__1472\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13553\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__13556\,
            I => \c0.data_in_frame_18_5\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__13553\,
            I => \c0.data_in_frame_18_5\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__13548\,
            I => \c0.n6225_cascade_\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__13545\,
            I => \c0.n6228_cascade_\
        );

    \I__1467\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13539\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__13539\,
            I => \N__13536\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__13536\,
            I => \N__13533\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__13533\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__13530\,
            I => \c0.n6267_cascade_\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__13527\,
            I => \c0.n6270_cascade_\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__13524\,
            I => \N__13521\
        );

    \I__1460\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13518\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__13518\,
            I => \N__13515\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__13515\,
            I => \N__13512\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__13512\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__13509\,
            I => \N__13506\
        );

    \I__1455\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13502\
        );

    \I__1454\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13499\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__13502\,
            I => \c0.data_in_frame_19_3\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__13499\,
            I => \c0.data_in_frame_19_3\
        );

    \I__1451\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13491\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__13491\,
            I => \N__13488\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__13488\,
            I => \c0.n22_adj_1876\
        );

    \I__1448\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13482\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13478\
        );

    \I__1446\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13474\
        );

    \I__1445\ : Span4Mux_s2_h
    port map (
            O => \N__13478\,
            I => \N__13471\
        );

    \I__1444\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13468\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__13474\,
            I => \c0.data_in_field_49\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__13471\,
            I => \c0.data_in_field_49\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__13468\,
            I => \c0.data_in_field_49\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__13461\,
            I => \c0.n5991_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__13458\,
            I => \N__13455\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__13455\,
            I => \N__13452\
        );

    \I__1437\ : Span4Mux_s2_h
    port map (
            O => \N__13452\,
            I => \N__13449\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__13449\,
            I => \c0.n6105\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__13446\,
            I => \c0.n5488_cascade_\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__13443\,
            I => \c0.n36_cascade_\
        );

    \I__1433\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13437\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__13437\,
            I => \c0.n45\
        );

    \I__1431\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13431\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__13431\,
            I => \c0.n12\
        );

    \I__1429\ : InMux
    port map (
            O => \N__13428\,
            I => \N__13425\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__13425\,
            I => \c0.n5488\
        );

    \I__1427\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13419\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__13419\,
            I => \c0.n5489\
        );

    \I__1425\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13413\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__13413\,
            I => \c0.n1886\
        );

    \I__1423\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13407\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__13407\,
            I => \c0.n1942\
        );

    \I__1421\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13401\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__13401\,
            I => \c0.n12_adj_1951\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__13398\,
            I => \N__13395\
        );

    \I__1418\ : InMux
    port map (
            O => \N__13395\,
            I => \N__13392\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__13392\,
            I => \N__13389\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__13389\,
            I => \N__13384\
        );

    \I__1415\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13381\
        );

    \I__1414\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13378\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__13384\,
            I => data_in_14_2
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__13381\,
            I => data_in_14_2
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__13378\,
            I => data_in_14_2
        );

    \I__1410\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13368\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13365\
        );

    \I__1408\ : Span4Mux_h
    port map (
            O => \N__13365\,
            I => \N__13362\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__13362\,
            I => \c0.n5536\
        );

    \I__1406\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13356\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__13356\,
            I => \c0.n5586\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__13353\,
            I => \c0.n5381_cascade_\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__13350\,
            I => \N__13347\
        );

    \I__1402\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13343\
        );

    \I__1401\ : InMux
    port map (
            O => \N__13346\,
            I => \N__13340\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__13343\,
            I => \N__13336\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__13340\,
            I => \N__13333\
        );

    \I__1398\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13330\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__13336\,
            I => data_in_13_7
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__13333\,
            I => data_in_13_7
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__13330\,
            I => data_in_13_7
        );

    \I__1394\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13320\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__13320\,
            I => \c0.n2009\
        );

    \I__1392\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13314\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__13308\,
            I => \N__13303\
        );

    \I__1388\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13300\
        );

    \I__1387\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13297\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__13303\,
            I => data_in_16_6
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__13300\,
            I => data_in_16_6
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__13297\,
            I => data_in_16_6
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__13290\,
            I => \c0.n1942_cascade_\
        );

    \I__1382\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13284\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__13284\,
            I => \c0.n18_adj_1938\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__13281\,
            I => \c0.n5578_cascade_\
        );

    \I__1379\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13275\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__13275\,
            I => \c0.n30\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__13272\,
            I => \c0.n6123_cascade_\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__13269\,
            I => \N__13266\
        );

    \I__1375\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13263\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__13263\,
            I => \c0.n5752\
        );

    \I__1373\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13256\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__13259\,
            I => \N__13253\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13249\
        );

    \I__1370\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13244\
        );

    \I__1369\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13244\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__13249\,
            I => data_in_14_7
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__13244\,
            I => data_in_14_7
        );

    \I__1366\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13236\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__13236\,
            I => \N__13233\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__13233\,
            I => \c0.n24_adj_1877\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__13230\,
            I => \N__13227\
        );

    \I__1362\ : InMux
    port map (
            O => \N__13227\,
            I => \N__13224\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__13224\,
            I => \N__13220\
        );

    \I__1360\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13217\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__13220\,
            I => \N__13214\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__13217\,
            I => \c0.data_in_frame_19_2\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__13214\,
            I => \c0.data_in_frame_19_2\
        );

    \I__1356\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13206\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__13206\,
            I => \c0.n5381\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__13203\,
            I => \c0.n6159_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13197\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__13197\,
            I => \N__13194\
        );

    \I__1351\ : Span4Mux_s2_h
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__13191\,
            I => \c0.n5737\
        );

    \I__1349\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__13185\,
            I => \c0.n5743\
        );

    \I__1347\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13179\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__13179\,
            I => \c0.n6141\
        );

    \I__1345\ : InMux
    port map (
            O => \N__13176\,
            I => \N__13171\
        );

    \I__1344\ : InMux
    port map (
            O => \N__13175\,
            I => \N__13166\
        );

    \I__1343\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13166\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__13171\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__13166\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13156\
        );

    \I__1339\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13151\
        );

    \I__1338\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13151\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__13156\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__13151\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1335\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13143\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__13143\,
            I => \c0.tx2.n316\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__13140\,
            I => \N__13137\
        );

    \I__1332\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13132\
        );

    \I__1331\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13129\
        );

    \I__1330\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13126\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13132\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__13129\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__13126\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1326\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13113\
        );

    \I__1325\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13110\
        );

    \I__1324\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13107\
        );

    \I__1323\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13104\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__13113\,
            I => \N__13101\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__13110\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__13107\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__13104\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__13101\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1317\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13089\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13086\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__13086\,
            I => \c0.tx2.n14_adj_1867\
        );

    \I__1314\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13080\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__13080\,
            I => \N__13077\
        );

    \I__1312\ : Odrv12
    port map (
            O => \N__13077\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \N__13071\
        );

    \I__1310\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13065\
        );

    \I__1309\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13062\
        );

    \I__1308\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13057\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13057\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__13065\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__13062\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__13057\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1303\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13042\
        );

    \I__1302\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13042\
        );

    \I__1301\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13037\
        );

    \I__1300\ : InMux
    port map (
            O => \N__13047\,
            I => \N__13037\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__13042\,
            I => \r_Clock_Count_8_adj_1994\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__13037\,
            I => \r_Clock_Count_8_adj_1994\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__13032\,
            I => \N__13027\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__13031\,
            I => \N__13023\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__13030\,
            I => \N__13020\
        );

    \I__1294\ : InMux
    port map (
            O => \N__13027\,
            I => \N__13017\
        );

    \I__1293\ : InMux
    port map (
            O => \N__13026\,
            I => \N__13014\
        );

    \I__1292\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13009\
        );

    \I__1291\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13009\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__13017\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13014\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__13009\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1287\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12998\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12995\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12998\,
            I => \c0.tx2.n31\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__12995\,
            I => \c0.tx2.n31\
        );

    \I__1283\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12987\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12984\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__12984\,
            I => \c0.tx2.n9\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__12981\,
            I => \c0.tx2.n5631_cascade_\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12974\
        );

    \I__1278\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12971\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__12974\,
            I => \c0.tx2.n78\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__12971\,
            I => \c0.tx2.n78\
        );

    \I__1275\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12953\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12953\
        );

    \I__1273\ : InMux
    port map (
            O => \N__12964\,
            I => \N__12950\
        );

    \I__1272\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12947\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12938\
        );

    \I__1270\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12938\
        );

    \I__1269\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12938\
        );

    \I__1268\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12938\
        );

    \I__1267\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12935\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__12953\,
            I => \N__12930\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N__12930\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__12947\,
            I => n4544
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__12938\,
            I => n4544
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__12935\,
            I => n4544
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__12930\,
            I => n4544
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__12921\,
            I => \N__12917\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__12920\,
            I => \N__12913\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12909\
        );

    \I__1257\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12906\
        );

    \I__1256\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12901\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12901\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12909\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__12906\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__12901\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__12894\,
            I => \N__12888\
        );

    \I__1250\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12885\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__12892\,
            I => \N__12878\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12873\
        );

    \I__1247\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12870\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__12885\,
            I => \N__12867\
        );

    \I__1245\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12858\
        );

    \I__1244\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12858\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12858\
        );

    \I__1242\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12858\
        );

    \I__1241\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12853\
        );

    \I__1240\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12853\
        );

    \I__1239\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12850\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__12873\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__12870\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__12867\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__12858\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__12853\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__12850\,
            I => \r_SM_Main_1_adj_1993\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__12837\,
            I => \c0.tx2.r_SM_Main_2_N_1767_1_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12831\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__12831\,
            I => \c0.tx2.n315\
        );

    \I__1229\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12825\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__12825\,
            I => \c0.tx2.n5824\
        );

    \I__1227\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12819\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__12819\,
            I => \c0.tx2.n5816\
        );

    \I__1225\ : InMux
    port map (
            O => \N__12816\,
            I => \N__12813\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12810\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__12810\,
            I => \c0.tx2.n314\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__12807\,
            I => \N__12804\
        );

    \I__1221\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12801\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__12801\,
            I => \c0.tx2.n319\
        );

    \I__1219\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12793\
        );

    \I__1218\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12788\
        );

    \I__1217\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12788\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__12793\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__12788\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1214\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12778\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12775\
        );

    \I__1212\ : InMux
    port map (
            O => \N__12781\,
            I => \N__12772\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__12778\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__12775\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__12772\,
            I => \c0.tx2.r_Bit_Index_2\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__12765\,
            I => \N__12761\
        );

    \I__1207\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12758\
        );

    \I__1206\ : InMux
    port map (
            O => \N__12761\,
            I => \N__12755\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__12758\,
            I => \c0.tx2.n1136\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__12755\,
            I => \c0.tx2.n1136\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__12750\,
            I => \n4_adj_1973_cascade_\
        );

    \I__1202\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12742\
        );

    \I__1201\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12737\
        );

    \I__1200\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12737\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__12742\,
            I => tx2_active
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__12737\,
            I => tx2_active
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__12732\,
            I => \N__12726\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__12731\,
            I => \N__12723\
        );

    \I__1195\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12717\
        );

    \I__1194\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12717\
        );

    \I__1193\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12710\
        );

    \I__1192\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12710\
        );

    \I__1191\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12710\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__12717\,
            I => \c0.r_SM_Main_2_N_1770_0\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__12710\,
            I => \c0.r_SM_Main_2_N_1770_0\
        );

    \I__1188\ : IoInMux
    port map (
            O => \N__12705\,
            I => \N__12701\
        );

    \I__1187\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12698\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__12701\,
            I => \N__12695\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__12698\,
            I => \N__12692\
        );

    \I__1184\ : Span4Mux_s1_h
    port map (
            O => \N__12695\,
            I => \N__12688\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__12692\,
            I => \N__12685\
        );

    \I__1182\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12682\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__12688\,
            I => tx2_o
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__12685\,
            I => tx2_o
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__12682\,
            I => tx2_o
        );

    \I__1178\ : IoInMux
    port map (
            O => \N__12675\,
            I => \N__12672\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__12672\,
            I => \N__12669\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__12669\,
            I => tx2_enable
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__12666\,
            I => \N__12663\
        );

    \I__1174\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12657\
        );

    \I__1172\ : Odrv12
    port map (
            O => \N__12657\,
            I => \c0.n6117\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__12654\,
            I => \c0.n5536_cascade_\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__12651\,
            I => \c0.n5570_cascade_\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12645\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__12645\,
            I => \c0.n27_adj_1910\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__12642\,
            I => \c0.n3689_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12636\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__12636\,
            I => \c0.tx2.n12\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__12630\,
            I => \c0.n3689\
        );

    \I__1162\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__12624\,
            I => \N__12619\
        );

    \I__1160\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12614\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12614\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__12619\,
            I => \c0.n3703\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__12614\,
            I => \c0.n3703\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \c0.n6282_cascade_\
        );

    \I__1155\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12603\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__12603\,
            I => \N__12600\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__12600\,
            I => \N__12597\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__12597\,
            I => \c0.n6132\
        );

    \I__1151\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12591\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__12591\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__12588\,
            I => \N__12585\
        );

    \I__1148\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12582\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__12582\,
            I => \c0.n6069\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__12579\,
            I => \c0.n6249_cascade_\
        );

    \I__1145\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12573\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12570\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__12570\,
            I => \c0.n28\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__12567\,
            I => \c0.n3703_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12561\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__12561\,
            I => \c0.n47\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__12558\,
            I => \c0.n52_cascade_\
        );

    \I__1138\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12552\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__12552\,
            I => \c0.n31\
        );

    \I__1136\ : InMux
    port map (
            O => \N__12549\,
            I => \N__12546\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__12543\,
            I => \c0.n32\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \c0.n24_adj_1879_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__12531\,
            I => \c0.n6102\
        );

    \I__1129\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12525\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__12525\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__1127\ : InMux
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__12519\,
            I => \N__12516\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__12516\,
            I => \c0.tx2.n6045\
        );

    \I__1124\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12510\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__12510\,
            I => \N__12506\
        );

    \I__1122\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12503\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__12506\,
            I => \N__12500\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__12503\,
            I => \c0.data_in_frame_18_2\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__12500\,
            I => \c0.data_in_frame_18_2\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__12495\,
            I => \c0.n6297_cascade_\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__1116\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12486\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__12486\,
            I => \c0.n6300\
        );

    \I__1114\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12480\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12476\
        );

    \I__1112\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12473\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__12476\,
            I => \N__12470\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__12473\,
            I => \c0.data_in_frame_18_3\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__12470\,
            I => \c0.data_in_frame_18_3\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__12465\,
            I => \c0.n6279_cascade_\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__12462\,
            I => \c0.n6075_cascade_\
        );

    \I__1106\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12456\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__12456\,
            I => \c0.n5773\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__12453\,
            I => \c0.n5454_cascade_\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__12450\,
            I => \c0.n27_cascade_\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__12447\,
            I => \N__12444\
        );

    \I__1101\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12441\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__12441\,
            I => \c0.n6063\
        );

    \I__1099\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12435\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__12435\,
            I => \c0.n5776\
        );

    \I__1097\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12429\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__12429\,
            I => \c0.n6099\
        );

    \I__1095\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12423\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__12423\,
            I => \N__12420\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__12420\,
            I => \N__12417\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__12417\,
            I => \c0.tx2.n6006\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__12414\,
            I => \c0.n5375_cascade_\
        );

    \I__1090\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12408\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__12408\,
            I => \N__12405\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__12405\,
            I => \c0.n5755\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__12402\,
            I => \c0.n6135_cascade_\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__12399\,
            I => \c0.n5746_cascade_\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__12396\,
            I => \c0.n6153_cascade_\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__12393\,
            I => \c0.n5740_cascade_\
        );

    \I__1083\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12387\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__12387\,
            I => \c0.n6129\
        );

    \I__1081\ : InMux
    port map (
            O => \N__12384\,
            I => \c0.tx2.n4779\
        );

    \I__1080\ : InMux
    port map (
            O => \N__12381\,
            I => \c0.tx2.n4780\
        );

    \I__1079\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__12375\,
            I => \c0.tx2.n318\
        );

    \I__1077\ : InMux
    port map (
            O => \N__12372\,
            I => \c0.tx2.n4781\
        );

    \I__1076\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__12366\,
            I => \c0.tx2.n317\
        );

    \I__1074\ : InMux
    port map (
            O => \N__12363\,
            I => \c0.tx2.n4782\
        );

    \I__1073\ : InMux
    port map (
            O => \N__12360\,
            I => \c0.tx2.n4783\
        );

    \I__1072\ : InMux
    port map (
            O => \N__12357\,
            I => \c0.tx2.n4784\
        );

    \I__1071\ : InMux
    port map (
            O => \N__12354\,
            I => \c0.tx2.n4785\
        );

    \I__1070\ : InMux
    port map (
            O => \N__12351\,
            I => \bfn_1_30_0_\
        );

    \I__1069\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12345\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__12345\,
            I => n313_adj_1997
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__12342\,
            I => \c0.tx2.o_Tx_Serial_N_1798_cascade_\
        );

    \I__1066\ : InMux
    port map (
            O => \N__12339\,
            I => \bfn_1_29_0_\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__12336\,
            I => \c0.n6027_cascade_\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__12333\,
            I => \c0.n5794_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12327\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__12327\,
            I => \c0.n6015\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \c0.n6072_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__12318\,
            I => \c0.n6018\
        );

    \I__1058\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__12312\,
            I => \N__12309\
        );

    \I__1056\ : Span4Mux_v
    port map (
            O => \N__12309\,
            I => \N__12306\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__12306\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__1053\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12297\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__12297\,
            I => \N__12294\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__12294\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__12291\,
            I => \c0.tx2.n6048_cascade_\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__12288\,
            I => \c0.n6057_cascade_\
        );

    \I__1048\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12282\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__12282\,
            I => \c0.n6306\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__12279\,
            I => \c0.n6060_cascade_\
        );

    \I__1045\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12273\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__12273\,
            I => \c0.n6087\
        );

    \I__1043\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12267\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__12267\,
            I => \N__12264\
        );

    \I__1041\ : Odrv12
    port map (
            O => \N__12264\,
            I => \c0.n5770\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__12261\,
            I => \c0.n5788_cascade_\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__12258\,
            I => \c0.n6111_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__12255\,
            I => \c0.n5758_cascade_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12249\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__12249\,
            I => \c0.n5761\
        );

    \I__1035\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12242\
        );

    \I__1034\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12239\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__12242\,
            I => \N__12236\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__12239\,
            I => \c0.data_in_frame_18_1\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__12236\,
            I => \c0.data_in_frame_18_1\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__12231\,
            I => \N__12228\
        );

    \I__1029\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12224\
        );

    \I__1028\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12221\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__12224\,
            I => \N__12218\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__12221\,
            I => \c0.data_in_frame_19_1\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__12218\,
            I => \c0.data_in_frame_19_1\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__12213\,
            I => \c0.n6303_cascade_\
        );

    \I__1023\ : IoInMux
    port map (
            O => \N__12210\,
            I => \N__12207\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__1021\ : IoSpan4Mux
    port map (
            O => \N__12204\,
            I => \N__12201\
        );

    \I__1020\ : IoSpan4Mux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__1019\ : IoSpan4Mux
    port map (
            O => \N__12198\,
            I => \N__12195\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__12195\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n4786\,
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n4771\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n4761\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n4746\,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4717,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4725,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n4733,
            carryinitout => \bfn_14_28_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12210\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35977\,
            in1 => \N__18121\,
            in2 => \_gnd_net_\,
            in3 => \N__16430\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i146_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__12245\,
            in1 => \N__15161\,
            in2 => \N__33217\,
            in3 => \N__32111\,
            lcout => \c0.data_in_frame_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i154_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__32144\,
            in2 => \N__26730\,
            in3 => \N__33083\,
            lcout => \c0.data_in_frame_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5749_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27756\,
            in1 => \N__19593\,
            in2 => \N__30175\,
            in3 => \N__23310\,
            lcout => OPEN,
            ltout => \c0.n6111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6111_bdd_4_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30105\,
            in1 => \N__31014\,
            in2 => \N__12258\,
            in3 => \N__20958\,
            lcout => OPEN,
            ltout => \c0.n5758_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5759_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__25257\,
            in1 => \N__25382\,
            in2 => \N__12255\,
            in3 => \N__12252\,
            lcout => \c0.n6099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1047_2_lut_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25256\,
            lcout => \c0.n1081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6105_bdd_4_lut_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__13458\,
            in1 => \N__28310\,
            in2 => \N__27299\,
            in3 => \N__30101\,
            lcout => \c0.n5761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__12246\,
            in1 => \N__30110\,
            in2 => \N__12231\,
            in3 => \N__27719\,
            lcout => OPEN,
            ltout => \c0.n6303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6303_bdd_4_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30111\,
            in1 => \N__30896\,
            in2 => \N__12213\,
            in3 => \N__17133\,
            lcout => \c0.n6306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5734_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__25260\,
            in1 => \N__12459\,
            in2 => \N__25407\,
            in3 => \N__12438\,
            lcout => OPEN,
            ltout => \c0.n6057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6057_bdd_4_lut_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__15927\,
            in1 => \N__25390\,
            in2 => \N__12288\,
            in3 => \N__12270\,
            lcout => OPEN,
            ltout => \c0.n6060_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__12285\,
            in1 => \N__14226\,
            in2 => \N__12279\,
            in3 => \N__13766\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37469\,
            ce => \N__13736\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5729_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27716\,
            in1 => \N__24316\,
            in2 => \N__30176\,
            in3 => \N__13485\,
            lcout => \c0.n6087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6081_bdd_4_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30109\,
            in1 => \N__27098\,
            in2 => \N__13842\,
            in3 => \N__17289\,
            lcout => \c0.n6084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15657\,
            in1 => \N__29433\,
            in2 => \N__14511\,
            in3 => \N__24918\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6087_bdd_4_lut_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__29949\,
            in1 => \N__16869\,
            in2 => \N__18921\,
            in3 => \N__12276\,
            lcout => \c0.n5770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6039_bdd_4_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29947\,
            in1 => \N__22242\,
            in2 => \N__27414\,
            in3 => \N__15300\,
            lcout => OPEN,
            ltout => \c0.n5788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6015_bdd_4_lut_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__25392\,
            in1 => \N__26751\,
            in2 => \N__12261\,
            in3 => \N__12330\,
            lcout => \c0.n6018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5680_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27717\,
            in1 => \N__28356\,
            in2 => \N__30070\,
            in3 => \N__21984\,
            lcout => OPEN,
            ltout => \c0.n6027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6027_bdd_4_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__25803\,
            in2 => \N__12336\,
            in3 => \N__16794\,
            lcout => OPEN,
            ltout => \c0.n5794_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5699_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__25391\,
            in1 => \N__25247\,
            in2 => \N__12333\,
            in3 => \N__14895\,
            lcout => \c0.n6015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6069_bdd_4_lut_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29999\,
            in1 => \N__28065\,
            in2 => \N__12588\,
            in3 => \N__30573\,
            lcout => OPEN,
            ltout => \c0.n6072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14225\,
            in1 => \N__13798\,
            in2 => \N__12324\,
            in3 => \N__12321\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37485\,
            ce => \N__13728\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i123_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35682\,
            in1 => \N__19294\,
            in2 => \_gnd_net_\,
            in3 => \N__15914\,
            lcout => data_in_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i107_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35683\,
            in1 => \N__13388\,
            in2 => \_gnd_net_\,
            in3 => \N__28367\,
            lcout => data_in_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n6045_bdd_4_lut_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__12315\,
            in1 => \N__13645\,
            in2 => \N__12303\,
            in3 => \N__12522\,
            lcout => OPEN,
            ltout => \c0.tx2.n6048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i367224_i1_3_lut_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12781\,
            in2 => \N__12291\,
            in3 => \N__12426\,
            lcout => OPEN,
            ltout => \c0.tx2.o_Tx_Serial_N_1798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i26_3_lut_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14024\,
            in2 => \N__12342\,
            in3 => \N__12893\,
            lcout => \c0.tx2.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__13929\,
            in1 => \_gnd_net_\,
            in2 => \N__13659\,
            in3 => \N__12783\,
            lcout => \c0.tx2.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => \N__13971\,
            sr => \N__13947\
        );

    \c0.tx2.r_Bit_Index_i1_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13646\,
            in2 => \_gnd_net_\,
            in3 => \N__13928\,
            lcout => \c0.tx2.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37509\,
            ce => \N__13971\,
            sr => \N__13947\
        );

    \c0.data_in_0___i143_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35509\,
            in1 => \N__18976\,
            in2 => \_gnd_net_\,
            in3 => \N__16145\,
            lcout => data_in_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i135_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18977\,
            in1 => \N__35510\,
            in2 => \_gnd_net_\,
            in3 => \N__13306\,
            lcout => data_in_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i3_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__12965\,
            in1 => \N__12378\,
            in2 => \N__14128\,
            in3 => \N__13118\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i4_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__12369\,
            in1 => \N__14104\,
            in2 => \N__12921\,
            in3 => \N__12966\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14025\,
            in1 => \N__12891\,
            in2 => \N__14127\,
            in3 => \N__13881\,
            lcout => \r_SM_Main_2_adj_1992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i127_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35500\,
            in1 => \N__13307\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => data_in_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_2_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12964\,
            in1 => \N__13176\,
            in2 => \_gnd_net_\,
            in3 => \N__12339\,
            lcout => \c0.tx2.n5824\,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => \c0.tx2.n4779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_3_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12958\,
            in1 => \N__13161\,
            in2 => \_gnd_net_\,
            in3 => \N__12384\,
            lcout => \c0.tx2.n5816\,
            ltout => OPEN,
            carryin => \c0.tx2.n4779\,
            carryout => \c0.tx2.n4780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_4_lut_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12798\,
            in2 => \_gnd_net_\,
            in3 => \N__12381\,
            lcout => \c0.tx2.n319\,
            ltout => OPEN,
            carryin => \c0.tx2.n4780\,
            carryout => \c0.tx2.n4781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_5_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13117\,
            in2 => \_gnd_net_\,
            in3 => \N__12372\,
            lcout => \c0.tx2.n318\,
            ltout => OPEN,
            carryin => \c0.tx2.n4781\,
            carryout => \c0.tx2.n4782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_6_lut_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12916\,
            in2 => \_gnd_net_\,
            in3 => \N__12363\,
            lcout => \c0.tx2.n317\,
            ltout => OPEN,
            carryin => \c0.tx2.n4782\,
            carryout => \c0.tx2.n4783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_7_lut_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13136\,
            in2 => \_gnd_net_\,
            in3 => \N__12360\,
            lcout => \c0.tx2.n316\,
            ltout => OPEN,
            carryin => \c0.tx2.n4783\,
            carryout => \c0.tx2.n4784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_8_lut_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13026\,
            in2 => \_gnd_net_\,
            in3 => \N__12357\,
            lcout => \c0.tx2.n315\,
            ltout => OPEN,
            carryin => \c0.tx2.n4784\,
            carryout => \c0.tx2.n4785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_9_lut_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13070\,
            in2 => \_gnd_net_\,
            in3 => \N__12354\,
            lcout => \c0.tx2.n314\,
            ltout => OPEN,
            carryin => \c0.tx2.n4785\,
            carryout => \c0.tx2.n4786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_10_lut_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13049\,
            in2 => \_gnd_net_\,
            in3 => \N__12351\,
            lcout => n313_adj_1997,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i8_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__13050\,
            in1 => \N__12348\,
            in2 => \N__14132\,
            in3 => \N__12963\,
            lcout => \r_Clock_Count_8_adj_1994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i124_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35976\,
            in1 => \N__14320\,
            in2 => \_gnd_net_\,
            in3 => \N__15200\,
            lcout => data_in_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i116_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35975\,
            in1 => \N__26353\,
            in2 => \_gnd_net_\,
            in3 => \N__14321\,
            lcout => data_in_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5769_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27748\,
            in1 => \N__20619\,
            in2 => \N__30185\,
            in3 => \N__14277\,
            lcout => OPEN,
            ltout => \c0.n6135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6135_bdd_4_lut_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__17223\,
            in1 => \N__30132\,
            in2 => \N__12402\,
            in3 => \N__22966\,
            lcout => OPEN,
            ltout => \c0.n5746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5789_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__13188\,
            in1 => \N__25406\,
            in2 => \N__12399\,
            in3 => \N__25258\,
            lcout => \c0.n6129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5784_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__14301\,
            in1 => \N__27747\,
            in2 => \N__18750\,
            in3 => \N__30144\,
            lcout => OPEN,
            ltout => \c0.n6153_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6153_bdd_4_lut_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30145\,
            in1 => \N__19110\,
            in2 => \N__12396\,
            in3 => \N__18471\,
            lcout => OPEN,
            ltout => \c0.n5740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6129_bdd_4_lut_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__13200\,
            in1 => \N__25403\,
            in2 => \N__12393\,
            in3 => \N__12390\,
            lcout => \c0.n6132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i132_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35974\,
            in1 => \N__21128\,
            in2 => \_gnd_net_\,
            in3 => \N__15193\,
            lcout => data_in_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5709_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27746\,
            in1 => \N__24365\,
            in2 => \N__30193\,
            in3 => \N__28196\,
            lcout => \c0.n6063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i148_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__12479\,
            in2 => \N__33273\,
            in3 => \N__14714\,
            lcout => \c0.data_in_frame_18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6063_bdd_4_lut_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__19392\,
            in1 => \N__29943\,
            in2 => \N__12447\,
            in3 => \N__19884\,
            lcout => \c0.n5776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i54_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__18488\,
            in1 => \_gnd_net_\,
            in2 => \N__21032\,
            in3 => \N__35942\,
            lcout => data_in_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6099_bdd_4_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__25386\,
            in1 => \N__12411\,
            in2 => \N__13269\,
            in3 => \N__12432\,
            lcout => \c0.n6102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i62_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35941\,
            in1 => \N__26575\,
            in2 => \_gnd_net_\,
            in3 => \N__18487\,
            lcout => data_in_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n6003_bdd_4_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__13542\,
            in1 => \N__13663\,
            in2 => \N__13524\,
            in3 => \N__13605\,
            lcout => \c0.tx2.n6006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_916_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17219\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24605\,
            lcout => OPEN,
            ltout => \c0.n5375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13239\,
            in1 => \N__13209\,
            in2 => \N__12414\,
            in3 => \N__13278\,
            lcout => \c0.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6117_bdd_4_lut_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30146\,
            in1 => \N__25842\,
            in2 => \N__12666\,
            in3 => \N__20559\,
            lcout => \c0.n5755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i147_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__12509\,
            in1 => \N__33250\,
            in2 => \N__32235\,
            in3 => \N__25734\,
            lcout => \c0.data_in_frame_18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i80_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__31341\,
            in1 => \N__32143\,
            in2 => \N__20925\,
            in3 => \N__33251\,
            lcout => \c0.data_in_field_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5719_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27718\,
            in1 => \N__23340\,
            in2 => \N__30069\,
            in3 => \N__14532\,
            lcout => OPEN,
            ltout => \c0.n6075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6075_bdd_4_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30053\,
            in1 => \N__17166\,
            in2 => \N__12462\,
            in3 => \N__15459\,
            lcout => \c0.n5773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_866_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20913\,
            in2 => \_gnd_net_\,
            in3 => \N__13477\,
            lcout => \c0.n5454\,
            ltout => \c0.n5454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_851_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16789\,
            in1 => \N__26959\,
            in2 => \N__12453\,
            in3 => \N__25112\,
            lcout => \c0.n1892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_932_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19641\,
            in2 => \_gnd_net_\,
            in3 => \N__21001\,
            lcout => \c0.n2009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_811_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21447\,
            in1 => \N__29514\,
            in2 => \N__14713\,
            in3 => \N__15512\,
            lcout => OPEN,
            ltout => \c0.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__30614\,
            in2 => \N__12450\,
            in3 => \N__17284\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i25_4_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17043\,
            in1 => \N__20874\,
            in2 => \N__15858\,
            in3 => \N__13440\,
            lcout => OPEN,
            ltout => \c0.n52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_812_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__12564\,
            in1 => \N__21933\,
            in2 => \N__12558\,
            in3 => \N__13422\,
            lcout => OPEN,
            ltout => \c0.n24_adj_1879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_839_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__12555\,
            in1 => \N__12549\,
            in2 => \N__12540\,
            in3 => \N__13359\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14217\,
            in1 => \N__13796\,
            in2 => \N__12492\,
            in3 => \N__12537\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37491\,
            ce => \N__13727\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__12594\,
            in1 => \N__12528\,
            in2 => \N__13664\,
            in3 => \N__13927\,
            lcout => \c0.tx2.n6045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5903_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__12513\,
            in1 => \N__29823\,
            in2 => \N__13230\,
            in3 => \N__27635\,
            lcout => OPEN,
            ltout => \c0.n6297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6297_bdd_4_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29824\,
            in1 => \N__15493\,
            in2 => \N__12495\,
            in3 => \N__15540\,
            lcout => \c0.n6300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5898_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__12483\,
            in1 => \N__29825\,
            in2 => \N__27702\,
            in3 => \N__13505\,
            lcout => OPEN,
            ltout => \c0.n6279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6279_bdd_4_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29826\,
            in1 => \N__16392\,
            in2 => \N__12465\,
            in3 => \N__22551\,
            lcout => OPEN,
            ltout => \c0.n6282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14218\,
            in1 => \N__13797\,
            in2 => \N__12609\,
            in3 => \N__12606\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37491\,
            ce => \N__13727\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_940_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15492\,
            in2 => \_gnd_net_\,
            in3 => \N__15539\,
            lcout => \c0.n2056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i131_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32474\,
            in1 => \N__32234\,
            in2 => \N__15508\,
            in3 => \N__15915\,
            lcout => \c0.data_in_field_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5714_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__27684\,
            in2 => \N__30148\,
            in3 => \N__15962\,
            lcout => \c0.n6069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5864_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__27683\,
            in1 => \N__30055\,
            in2 => \N__24543\,
            in3 => \N__18380\,
            lcout => OPEN,
            ltout => \c0.n6249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6249_bdd_4_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30054\,
            in1 => \N__30615\,
            in2 => \N__12579\,
            in3 => \N__28005\,
            lcout => \c0.n5695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i115_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35501\,
            in1 => \N__13387\,
            in2 => \_gnd_net_\,
            in3 => \N__19301\,
            lcout => data_in_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i64_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15611\,
            in1 => \N__35502\,
            in2 => \_gnd_net_\,
            in3 => \N__23249\,
            lcout => data_in_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3459_4_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32233\,
            in1 => \N__12648\,
            in2 => \N__15378\,
            in3 => \N__12576\,
            lcout => \c0.n3703\,
            ltout => \c0.n3703_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5628_2_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__32372\,
            in1 => \_gnd_net_\,
            in2 => \N__12567\,
            in3 => \_gnd_net_\,
            lcout => \c0.n2325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5754_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27546\,
            in1 => \N__14598\,
            in2 => \N__29924\,
            in3 => \N__24806\,
            lcout => \c0.n6117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_846_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29562\,
            in2 => \_gnd_net_\,
            in3 => \N__18381\,
            lcout => \c0.n5536\,
            ltout => \c0.n5536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_827_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17058\,
            in1 => \N__14433\,
            in2 => \N__12654\,
            in3 => \N__16992\,
            lcout => OPEN,
            ltout => \c0.n5570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_840_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101111"
        )
    port map (
            in0 => \N__19356\,
            in1 => \N__20448\,
            in2 => \N__12651\,
            in3 => \N__22380\,
            lcout => \c0.n27_adj_1910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i489_3_lut_4_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__12746\,
            in1 => \N__12730\,
            in2 => \N__32437\,
            in3 => \N__12622\,
            lcout => \c0.n195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3445_2_lut_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12729\,
            lcout => \c0.n3689\,
            ltout => \c0.n3689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000110011"
        )
    port map (
            in0 => \N__13591\,
            in1 => \N__12627\,
            in2 => \N__12642\,
            in3 => \N__32379\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__14126\,
            in1 => \N__12691\,
            in2 => \_gnd_net_\,
            in3 => \N__12639\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_1801_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001001111"
        )
    port map (
            in0 => \N__12633\,
            in1 => \N__13592\,
            in2 => \N__32438\,
            in3 => \N__12623\,
            lcout => \c0.r_SM_Main_2_N_1770_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i895_2_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12782\,
            in2 => \_gnd_net_\,
            in3 => \N__13644\,
            lcout => \c0.tx2.n1136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i28_4_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__12764\,
            in1 => \N__12722\,
            in2 => \N__12894\,
            in3 => \N__13854\,
            lcout => \c0.tx2.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2088_4_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__12882\,
            in1 => \N__13914\,
            in2 => \N__12765\,
            in3 => \N__13963\,
            lcout => n2339,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5614_4_lut_4_lut_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__12883\,
            in1 => \N__14011\,
            in2 => \N__12731\,
            in3 => \N__13879\,
            lcout => OPEN,
            ltout => \n4_adj_1973_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__14100\,
            in1 => \N__12747\,
            in2 => \N__12750\,
            in3 => \N__12884\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12881\,
            in1 => \N__14099\,
            in2 => \N__12732\,
            in3 => \N__14012\,
            lcout => \c0.tx2.n1624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12704\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__17695\,
            in2 => \N__18023\,
            in3 => \N__17645\,
            lcout => \r_SM_Main_2_adj_1989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__14115\,
            in1 => \N__14007\,
            in2 => \N__12892\,
            in3 => \N__13880\,
            lcout => \r_SM_Main_1_adj_1993\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i3_4_lut_adj_799_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__12876\,
            in1 => \N__12912\,
            in2 => \N__14017\,
            in3 => \N__13116\,
            lcout => \c0.tx2.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7_4_lut_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12977\,
            in1 => \N__13092\,
            in2 => \N__12920\,
            in3 => \N__13001\,
            lcout => \c0.tx2.r_SM_Main_2_N_1767_1\,
            ltout => \c0.tx2.r_SM_Main_2_N_1767_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_4_lut_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__14006\,
            in1 => \N__12877\,
            in2 => \N__12837\,
            in3 => \N__14114\,
            lcout => n2208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_793_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__13848\,
            in1 => \N__16286\,
            in2 => \N__18022\,
            in3 => \N__20300\,
            lcout => \c0.rx.n359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i6_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__12834\,
            in1 => \N__12961\,
            in2 => \N__13032\,
            in3 => \N__14125\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13175\,
            in1 => \N__12828\,
            in2 => \_gnd_net_\,
            in3 => \N__14111\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i1_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12822\,
            in1 => \N__14123\,
            in2 => \_gnd_net_\,
            in3 => \N__13160\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i7_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__12960\,
            in1 => \N__12816\,
            in2 => \N__13074\,
            in3 => \N__14113\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i2_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__12797\,
            in1 => \N__12962\,
            in2 => \N__12807\,
            in3 => \N__14124\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i85_2_lut_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12796\,
            in2 => \_gnd_net_\,
            in3 => \N__13135\,
            lcout => \c0.tx2.n78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13174\,
            in2 => \_gnd_net_\,
            in3 => \N__13159\,
            lcout => \c0.tx2.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i5_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__12959\,
            in1 => \N__13146\,
            in2 => \N__13140\,
            in3 => \N__14112\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i6_4_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__13119\,
            in2 => \N__13030\,
            in3 => \N__13047\,
            lcout => \c0.tx2.n14_adj_1867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13083\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5285_4_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13069\,
            in1 => \N__13048\,
            in2 => \N__13031\,
            in3 => \N__13002\,
            lcout => OPEN,
            ltout => \c0.tx2.n5631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_adj_800_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__14119\,
            in1 => \N__12990\,
            in2 => \N__12981\,
            in3 => \N__12978\,
            lcout => n4544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i44_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35943\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__16694\,
            lcout => data_in_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i60_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32063\,
            in1 => \N__33138\,
            in2 => \N__14247\,
            in3 => \N__14297\,
            lcout => \c0.data_in_field_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i60_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35944\,
            in1 => \N__14242\,
            in2 => \_gnd_net_\,
            in3 => \N__14390\,
            lcout => data_in_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5794_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27749\,
            in1 => \N__18609\,
            in2 => \N__30208\,
            in3 => \N__22593\,
            lcout => OPEN,
            ltout => \c0.n6159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6159_bdd_4_lut_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30186\,
            in1 => \N__18654\,
            in2 => \N__13203\,
            in3 => \N__14414\,
            lcout => \c0.n5737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6141_bdd_4_lut_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__13182\,
            in1 => \N__19026\,
            in2 => \N__30207\,
            in3 => \N__14365\,
            lcout => \c0.n5743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5774_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27608\,
            in1 => \N__18572\,
            in2 => \N__30059\,
            in3 => \N__27957\,
            lcout => \c0.n6141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_850_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18466\,
            in1 => \N__14773\,
            in2 => \_gnd_net_\,
            in3 => \N__14364\,
            lcout => \c0.n2095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16416\,
            in1 => \N__18194\,
            in2 => \_gnd_net_\,
            in3 => \N__35939\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i120_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21872\,
            in1 => \_gnd_net_\,
            in2 => \N__36023\,
            in3 => \N__13252\,
            lcout => data_in_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i120_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__14774\,
            in1 => \N__33026\,
            in2 => \N__13259\,
            in3 => \N__31850\,
            lcout => \c0.data_in_field_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i104_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35935\,
            in1 => \N__13346\,
            in2 => \_gnd_net_\,
            in3 => \N__18841\,
            lcout => data_in_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i68_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35933\,
            in1 => \N__18671\,
            in2 => \_gnd_net_\,
            in3 => \N__14383\,
            lcout => data_in_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5764_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27753\,
            in1 => \N__23025\,
            in2 => \N__30060\,
            in3 => \N__16827\,
            lcout => OPEN,
            ltout => \c0.n6123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6123_bdd_4_lut_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30147\,
            in1 => \N__27261\,
            in2 => \N__13272\,
            in3 => \N__16905\,
            lcout => \c0.n5752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i112_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35932\,
            in1 => \N__13260\,
            in2 => \_gnd_net_\,
            in3 => \N__13339\,
            lcout => data_in_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_adj_983_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28195\,
            in1 => \N__24119\,
            in2 => \_gnd_net_\,
            in3 => \N__22968\,
            lcout => \c0.n24_adj_1877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i84_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16944\,
            in1 => \N__35934\,
            in2 => \_gnd_net_\,
            in3 => \N__14464\,
            lcout => data_in_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i140_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35681\,
            in1 => \N__21127\,
            in2 => \_gnd_net_\,
            in3 => \N__14715\,
            lcout => data_in_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i155_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32071\,
            in1 => \N__13223\,
            in2 => \N__25908\,
            in3 => \N__32978\,
            lcout => \c0.data_in_frame_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_854_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20614\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27097\,
            lcout => \c0.n5381\,
            ltout => \c0.n5381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__15777\,
            in2 => \N__13353\,
            in3 => \N__16381\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_902_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__24870\,
            in2 => \N__28311\,
            in3 => \N__26799\,
            lcout => \c0.n18_adj_1938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i112_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32977\,
            in1 => \N__32072\,
            in2 => \N__13350\,
            in3 => \N__14753\,
            lcout => \c0.data_in_field_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20171\,
            in1 => \N__13323\,
            in2 => \N__24355\,
            in3 => \N__27042\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i82_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32064\,
            in1 => \N__17844\,
            in2 => \N__32778\,
            in3 => \N__14531\,
            lcout => \c0.data_in_field_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i135_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__17031\,
            in1 => \N__13317\,
            in2 => \N__32217\,
            in3 => \N__32598\,
            lcout => \c0.data_in_field_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i96_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__20843\,
            in1 => \N__26163\,
            in2 => \N__32779\,
            in3 => \N__32076\,
            lcout => \c0.data_in_field_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_921_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20842\,
            in1 => \N__20811\,
            in2 => \_gnd_net_\,
            in3 => \N__14530\,
            lcout => \c0.n1942\,
            ltout => \c0.n1942_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_920_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25148\,
            in1 => \N__18577\,
            in2 => \N__13290\,
            in3 => \N__19879\,
            lcout => \c0.n5578\,
            ltout => \c0.n5578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_984_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13287\,
            in1 => \N__17106\,
            in2 => \N__13281\,
            in3 => \N__20892\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_972_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23238\,
            in1 => \N__25517\,
            in2 => \N__15351\,
            in3 => \N__13404\,
            lcout => \c0.n5488\,
            ltout => \c0.n5488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_2_lut_3_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14418\,
            in2 => \N__13446\,
            in3 => \N__16391\,
            lcout => OPEN,
            ltout => \c0.n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__15840\,
            in2 => \N__13443\,
            in3 => \N__21769\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_810_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13434\,
            in1 => \N__13416\,
            in2 => \N__15165\,
            in3 => \N__13428\,
            lcout => \c0.n5489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_909_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18578\,
            in2 => \_gnd_net_\,
            in3 => \N__19880\,
            lcout => \c0.n1886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_970_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13410\,
            in1 => \N__16967\,
            in2 => \N__15762\,
            in3 => \N__14486\,
            lcout => \c0.n12_adj_1951\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i115_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32982\,
            in1 => \N__32067\,
            in2 => \N__13398\,
            in3 => \N__17086\,
            lcout => \c0.data_in_field_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13371\,
            in1 => \N__15630\,
            in2 => \N__14637\,
            in3 => \N__14538\,
            lcout => \c0.n5586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i156_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__32065\,
            in1 => \N__15747\,
            in2 => \N__13509\,
            in3 => \N__32985\,
            lcout => \c0.data_in_frame_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i72_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36024\,
            in1 => \N__31337\,
            in2 => \_gnd_net_\,
            in3 => \N__15598\,
            lcout => data_in_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16904\,
            in1 => \N__18431\,
            in2 => \_gnd_net_\,
            in3 => \N__18743\,
            lcout => \c0.n22_adj_1876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i139_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32983\,
            in1 => \N__32068\,
            in2 => \N__15551\,
            in3 => \N__25695\,
            lcout => \c0.data_in_field_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i50_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32066\,
            in1 => \N__32984\,
            in2 => \N__22484\,
            in3 => \N__13481\,
            lcout => \c0.data_in_field_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5652_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__28130\,
            in1 => \N__27647\,
            in2 => \N__20859\,
            in3 => \N__29802\,
            lcout => OPEN,
            ltout => \c0.n5991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5991_bdd_4_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29803\,
            in1 => \N__30779\,
            in2 => \N__13461\,
            in3 => \N__20924\,
            lcout => \c0.n5994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i119_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__32756\,
            in1 => \N__19818\,
            in2 => \N__18791\,
            in3 => \N__32070\,
            lcout => \c0.data_in_field_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5744_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27646\,
            in1 => \N__17085\,
            in2 => \N__29938\,
            in3 => \N__24606\,
            lcout => \c0.n6105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i79_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36043\,
            in1 => \N__31183\,
            in2 => \_gnd_net_\,
            in3 => \N__17474\,
            lcout => data_in_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i96_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26158\,
            in1 => \N__36044\,
            in2 => \_gnd_net_\,
            in3 => \N__18854\,
            lcout => data_in_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i150_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32069\,
            in1 => \N__13560\,
            in2 => \N__21399\,
            in3 => \N__32757\,
            lcout => \c0.data_in_frame_18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5849_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27633\,
            in1 => \N__19839\,
            in2 => \N__30126\,
            in3 => \N__13559\,
            lcout => OPEN,
            ltout => \c0.n6225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6225_bdd_4_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__30025\,
            in2 => \N__13548\,
            in3 => \N__27168\,
            lcout => OPEN,
            ltout => \c0.n6228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14220\,
            in1 => \N__13789\,
            in2 => \N__13545\,
            in3 => \N__23589\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => \N__13737\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5879_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27634\,
            in1 => \N__17544\,
            in2 => \N__30127\,
            in3 => \N__14829\,
            lcout => OPEN,
            ltout => \c0.n6267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6267_bdd_4_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__29827\,
            in1 => \N__20742\,
            in2 => \N__13530\,
            in3 => \N__18888\,
            lcout => OPEN,
            ltout => \c0.n6270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__14219\,
            in1 => \N__13788\,
            in2 => \N__13527\,
            in3 => \N__14649\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37510\,
            ce => \N__13737\,
            sr => \_gnd_net_\
        );

    \c0.i5622_4_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__13787\,
            in1 => \N__30018\,
            in2 => \N__14221\,
            in3 => \N__27632\,
            lcout => \c0.FRAME_MATCHER_wait_for_transmission_N_909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5724_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__16095\,
            in1 => \N__29782\,
            in2 => \N__19752\,
            in3 => \N__27557\,
            lcout => \c0.n6081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__13827\,
            in1 => \N__14207\,
            in2 => \N__13803\,
            in3 => \N__14721\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => \N__13732\,
            sr => \_gnd_net_\
        );

    \c0.n6231_bdd_4_lut_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__13812\,
            in1 => \N__25306\,
            in2 => \N__14790\,
            in3 => \N__17523\,
            lcout => OPEN,
            ltout => \c0.n6234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__14847\,
            in1 => \N__14206\,
            in2 => \N__13806\,
            in3 => \N__13802\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37522\,
            ce => \N__13732\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_5690_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__13680\,
            in1 => \N__13674\,
            in2 => \N__13668\,
            in3 => \N__13918\,
            lcout => \c0.tx2.n6003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_525_526__i1_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27568\,
            in2 => \N__13593\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \c0.n4735\,
            clk => \N__37534\,
            ce => \N__14157\,
            sr => \N__14148\
        );

    \c0.byte_transmit_counter2_525_526__i2_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29792\,
            in2 => \_gnd_net_\,
            in3 => \N__13569\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n4735\,
            carryout => \c0.n4736\,
            clk => \N__37534\,
            ce => \N__14157\,
            sr => \N__14148\
        );

    \c0.byte_transmit_counter2_525_526__i3_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25238\,
            in2 => \_gnd_net_\,
            in3 => \N__13566\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \c0.n4736\,
            carryout => \c0.n4737\,
            clk => \N__37534\,
            ce => \N__14157\,
            sr => \N__14148\
        );

    \c0.byte_transmit_counter2_525_526__i4_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25305\,
            in2 => \_gnd_net_\,
            in3 => \N__13563\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \c0.n4737\,
            carryout => \c0.n4738\,
            clk => \N__37534\,
            ce => \N__14157\,
            sr => \N__14148\
        );

    \c0.byte_transmit_counter2_525_526__i5_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14205\,
            in2 => \_gnd_net_\,
            in3 => \N__14229\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37534\,
            ce => \N__14157\,
            sr => \N__14148\
        );

    \c0.tx2.r_SM_Main_i0_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__14016\,
            in1 => \N__13878\,
            in2 => \N__14136\,
            in3 => \N__14031\,
            lcout => \c0.tx2.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__13913\,
            in1 => \N__13964\,
            in2 => \_gnd_net_\,
            in3 => \N__13940\,
            lcout => \r_Bit_Index_0_adj_1995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16208\,
            in1 => \N__14997\,
            in2 => \_gnd_net_\,
            in3 => \N__14880\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5567_2_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13912\,
            in2 => \_gnd_net_\,
            in3 => \N__13877\,
            lcout => \c0.tx2.n5847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16209\,
            in1 => \N__14868\,
            in2 => \_gnd_net_\,
            in3 => \N__15069\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i16_4_lut_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111111"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__17630\,
            in2 => \N__18024\,
            in3 => \N__14334\,
            lcout => \c0.rx.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5570_2_lut_3_lut_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15014\,
            in1 => \N__14994\,
            in2 => \_gnd_net_\,
            in3 => \N__14955\,
            lcout => \c0.rx.n5823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_adj_794_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14993\,
            in1 => \N__14953\,
            in2 => \N__17697\,
            in3 => \N__15015\,
            lcout => \c0.rx.n3589\,
            ltout => \c0.rx.n3589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5560_2_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14340\,
            in3 => \N__20299\,
            lcout => \c0.rx.n5815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__14992\,
            in1 => \N__14952\,
            in2 => \N__20316\,
            in3 => \N__15012\,
            lcout => OPEN,
            ltout => \c0.rx.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5574_4_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__15013\,
            in1 => \N__17691\,
            in2 => \N__14337\,
            in3 => \N__15087\,
            lcout => \c0.rx.n5817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i59_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35641\,
            in1 => \N__14614\,
            in2 => \_gnd_net_\,
            in3 => \N__16736\,
            lcout => data_in_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i124_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33077\,
            in1 => \N__32125\,
            in2 => \N__14328\,
            in3 => \N__14271\,
            lcout => \c0.data_in_field_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i51_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36070\,
            in1 => \N__14621\,
            in2 => \_gnd_net_\,
            in3 => \N__25643\,
            lcout => data_in_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_939_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14273\,
            in1 => \N__14293\,
            in2 => \_gnd_net_\,
            in3 => \N__18653\,
            lcout => \c0.n1979\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_980_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14272\,
            in1 => \N__14409\,
            in2 => \N__14367\,
            in3 => \N__16361\,
            lcout => \c0.n1926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i52_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14246\,
            in1 => \N__36071\,
            in2 => \_gnd_net_\,
            in3 => \N__16462\,
            lcout => data_in_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i12_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__16497\,
            in1 => \N__32124\,
            in2 => \N__33219\,
            in3 => \N__14410\,
            lcout => \c0.data_in_field_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i105_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__33174\,
            in1 => \N__31847\,
            in2 => \N__14922\,
            in3 => \N__19671\,
            lcout => \c0.data_in_field_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i24_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31845\,
            in1 => \N__33175\,
            in2 => \N__16426\,
            in3 => \N__15266\,
            lcout => \c0.data_in_field_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6183_bdd_4_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30172\,
            in1 => \N__24897\,
            in2 => \N__16680\,
            in3 => \N__19640\,
            lcout => \c0.n5725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i138_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36069\,
            in1 => \N__15568\,
            in2 => \_gnd_net_\,
            in3 => \N__15148\,
            lcout => data_in_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i76_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35962\,
            in1 => \N__18670\,
            in2 => \_gnd_net_\,
            in3 => \N__14465\,
            lcout => data_in_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i16_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__18133\,
            in1 => \N__31848\,
            in2 => \N__33245\,
            in3 => \N__15315\,
            lcout => \c0.data_in_field_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i68_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31846\,
            in1 => \N__33176\,
            in2 => \N__14391\,
            in3 => \N__14366\,
            lcout => \c0.data_in_field_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i66_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35940\,
            in1 => \N__17820\,
            in2 => \_gnd_net_\,
            in3 => \N__16510\,
            lcout => data_in_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i122_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36064\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__15815\,
            lcout => data_in_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_883_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14914\,
            in2 => \_gnd_net_\,
            in3 => \N__16641\,
            lcout => \c0.n2143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i26_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__22316\,
            in1 => \N__32211\,
            in2 => \N__30828\,
            in3 => \N__33081\,
            lcout => \c0.data_in_field_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_adj_815_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17212\,
            in2 => \_gnd_net_\,
            in3 => \N__16790\,
            lcout => \c0.n16_adj_1880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i84_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__14466\,
            in1 => \N__32212\,
            in2 => \N__18579\,
            in3 => \N__33082\,
            lcout => \c0.data_in_field_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__36068\,
            in2 => \_gnd_net_\,
            in3 => \N__18279\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i58_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16511\,
            in1 => \_gnd_net_\,
            in2 => \N__36075\,
            in3 => \N__16066\,
            lcout => data_in_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_915_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27327\,
            lcout => OPEN,
            ltout => \c0.n5412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_816_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15276\,
            in1 => \N__28188\,
            in2 => \N__14448\,
            in3 => \N__18430\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1881_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_818_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14445\,
            in1 => \N__24807\,
            in2 => \N__14436\,
            in3 => \N__25524\,
            lcout => \c0.n24_adj_1884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_872_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29607\,
            in1 => \N__14749\,
            in2 => \_gnd_net_\,
            in3 => \N__14529\,
            lcout => \c0.n2134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i107_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__27286\,
            in1 => \N__32868\,
            in2 => \N__28395\,
            in3 => \N__32227\,
            lcout => \c0.data_in_field_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_879_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17010\,
            in1 => \N__27284\,
            in2 => \_gnd_net_\,
            in3 => \N__14806\,
            lcout => \c0.n5554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i15_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__14807\,
            in1 => \N__32869\,
            in2 => \N__18162\,
            in3 => \N__32228\,
            lcout => \c0.data_in_field_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i130_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36072\,
            in1 => \N__15575\,
            in2 => \_gnd_net_\,
            in3 => \N__15808\,
            lcout => data_in_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_960_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24536\,
            in1 => \N__22364\,
            in2 => \_gnd_net_\,
            in3 => \N__29608\,
            lcout => \c0.n5551\,
            ltout => \c0.n5551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1007_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24344\,
            in2 => \N__14496\,
            in3 => \N__24299\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i48_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__32860\,
            in1 => \N__29612\,
            in2 => \N__32284\,
            in3 => \N__27195\,
            lcout => \c0.data_in_field_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22793\,
            in1 => \N__20523\,
            in2 => \N__19731\,
            in3 => \N__14493\,
            lcout => OPEN,
            ltout => \c0.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_836_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011111111"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__21147\,
            in2 => \N__14469\,
            in3 => \N__15699\,
            lcout => \c0.n20_adj_1905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i114_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__24345\,
            in1 => \N__32861\,
            in2 => \N__19503\,
            in3 => \N__32226\,
            lcout => \c0.data_in_field_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14556\,
            in1 => \N__25463\,
            in2 => \_gnd_net_\,
            in3 => \N__28131\,
            lcout => \c0.n18_adj_1904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5804_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__19206\,
            in1 => \N__27667\,
            in2 => \N__30171\,
            in3 => \N__29558\,
            lcout => OPEN,
            ltout => \c0.n6177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6177_bdd_4_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__15687\,
            in1 => \N__17577\,
            in2 => \N__14547\,
            in3 => \N__30089\,
            lcout => OPEN,
            ltout => \c0.n5728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5814_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__25372\,
            in1 => \N__25248\,
            in2 => \N__14544\,
            in3 => \N__21501\,
            lcout => \c0.n6165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_946_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17285\,
            in1 => \N__25995\,
            in2 => \N__19209\,
            in3 => \N__17241\,
            lcout => \c0.n1973\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i58_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32240\,
            in1 => \N__32643\,
            in2 => \N__16080\,
            in3 => \N__24309\,
            lcout => \c0.data_in_field_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16131\,
            in2 => \_gnd_net_\,
            in3 => \N__15544\,
            lcout => OPEN,
            ltout => \c0.n16_adj_1873_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15441\,
            in1 => \N__15882\,
            in2 => \N__14541\,
            in3 => \N__17445\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6165_bdd_4_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__21717\,
            in1 => \N__14667\,
            in2 => \N__25408\,
            in3 => \N__14658\,
            lcout => \c0.n6168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15440\,
            in1 => \N__30518\,
            in2 => \N__30882\,
            in3 => \N__15872\,
            lcout => \c0.n2012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i159_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__32201\,
            in1 => \N__14570\,
            in2 => \N__32988\,
            in3 => \N__15983\,
            lcout => \c0.data_in_frame_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i74_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__17819\,
            in1 => \N__32202\,
            in2 => \N__15457\,
            in3 => \N__32777\,
            lcout => \c0.data_in_field_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6213_bdd_4_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__29939\,
            in1 => \N__21228\,
            in2 => \N__15474\,
            in3 => \N__23237\,
            lcout => \c0.n5710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i86_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32705\,
            in1 => \N__32219\,
            in2 => \N__28857\,
            in3 => \N__25134\,
            lcout => \c0.data_in_field_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28239\,
            in1 => \N__28349\,
            in2 => \N__14594\,
            in3 => \N__16826\,
            lcout => \c0.n20_adj_1878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i59_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32704\,
            in1 => \N__32218\,
            in2 => \N__14628\,
            in3 => \N__14590\,
            lcout => \c0.data_in_field_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1009_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14586\,
            in1 => \N__28348\,
            in2 => \N__17087\,
            in3 => \N__26848\,
            lcout => \c0.n5575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5779_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__16110\,
            in1 => \N__29970\,
            in2 => \N__14571\,
            in3 => \N__27648\,
            lcout => OPEN,
            ltout => \c0.n6147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6147_bdd_4_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__29971\,
            in1 => \N__18963\,
            in2 => \N__14850\,
            in3 => \N__17026\,
            lcout => \c0.n6150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i157_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__14828\,
            in1 => \N__20657\,
            in2 => \N__32916\,
            in3 => \N__32220\,
            lcout => \c0.data_in_frame_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5874_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__17354\,
            in2 => \N__30128\,
            in3 => \N__19281\,
            lcout => OPEN,
            ltout => \c0.n6255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6255_bdd_4_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__29929\,
            in1 => \N__14814\,
            in2 => \N__14793\,
            in3 => \N__16650\,
            lcout => \c0.n5692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5884_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27665\,
            in1 => \N__14781\,
            in2 => \N__30061\,
            in3 => \N__19473\,
            lcout => OPEN,
            ltout => \c0.n6273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6273_bdd_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30029\,
            in1 => \N__19143\,
            in2 => \N__14760\,
            in3 => \N__14757\,
            lcout => OPEN,
            ltout => \c0.n5686_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__14733\,
            in1 => \N__25404\,
            in2 => \N__14727\,
            in3 => \N__25231\,
            lcout => OPEN,
            ltout => \c0.n6261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6261_bdd_4_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__25405\,
            in1 => \N__15327\,
            in2 => \N__14724\,
            in3 => \N__29580\,
            lcout => \c0.n6264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i148_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15746\,
            in1 => \N__35384\,
            in2 => \_gnd_net_\,
            in3 => \N__14694\,
            lcout => data_in_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37535\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5675_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27607\,
            in1 => \N__17372\,
            in2 => \N__29925\,
            in3 => \N__25572\,
            lcout => OPEN,
            ltout => \c0.n6021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6021_bdd_4_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__29786\,
            in1 => \N__14921\,
            in2 => \N__14898\,
            in3 => \N__20809\,
            lcout => \c0.n5797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15122\,
            in1 => \N__14954\,
            in2 => \_gnd_net_\,
            in3 => \N__14883\,
            lcout => \c0.rx.n5855\,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => \c0.rx.n4772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15108\,
            in1 => \N__14996\,
            in2 => \_gnd_net_\,
            in3 => \N__14874\,
            lcout => \c0.rx.n5860\,
            ltout => OPEN,
            carryin => \c0.rx.n4772\,
            carryout => \c0.rx.n4773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15121\,
            in1 => \N__16009\,
            in2 => \_gnd_net_\,
            in3 => \N__14871\,
            lcout => \c0.rx.n5822\,
            ltout => OPEN,
            carryin => \c0.rx.n4773\,
            carryout => \c0.rx.n4774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15107\,
            in1 => \N__15068\,
            in2 => \_gnd_net_\,
            in3 => \N__14862\,
            lcout => \c0.rx.n5856\,
            ltout => OPEN,
            carryin => \c0.rx.n4774\,
            carryout => \c0.rx.n4775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15120\,
            in1 => \_gnd_net_\,
            in2 => \N__15234\,
            in3 => \N__14859\,
            lcout => \c0.rx.n5857\,
            ltout => OPEN,
            carryin => \c0.rx.n4775\,
            carryout => \c0.rx.n4776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15109\,
            in1 => \N__15035\,
            in2 => \_gnd_net_\,
            in3 => \N__14856\,
            lcout => \c0.rx.n5858\,
            ltout => OPEN,
            carryin => \c0.rx.n4776\,
            carryout => \c0.rx.n4777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15123\,
            in1 => \N__15051\,
            in2 => \_gnd_net_\,
            in3 => \N__14853\,
            lcout => \c0.rx.n5854\,
            ltout => OPEN,
            carryin => \c0.rx.n4777\,
            carryout => \c0.rx.n4778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15110\,
            in1 => \N__16172\,
            in2 => \_gnd_net_\,
            in3 => \N__15090\,
            lcout => \c0.rx.n5859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14991\,
            in2 => \_gnd_net_\,
            in3 => \N__14949\,
            lcout => \c0.rx.n5361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15036\,
            in1 => \N__16212\,
            in2 => \_gnd_net_\,
            in3 => \N__15081\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__15050\,
            in1 => \_gnd_net_\,
            in2 => \N__16222\,
            in3 => \N__15075\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_3_lut_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__15067\,
            in1 => \N__15229\,
            in2 => \_gnd_net_\,
            in3 => \N__15049\,
            lcout => OPEN,
            ltout => \c0.rx.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5277_4_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15034\,
            in1 => \N__16011\,
            in2 => \N__15018\,
            in3 => \N__16171\,
            lcout => \c0.rx.n1724\,
            ltout => \c0.rx.n1724_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__14950\,
            in1 => \_gnd_net_\,
            in2 => \N__15000\,
            in3 => \N__14995\,
            lcout => \r_SM_Main_2_N_1824_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16210\,
            in1 => \N__14951\,
            in2 => \_gnd_net_\,
            in3 => \N__14961\,
            lcout => \c0.rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15233\,
            in1 => \N__15240\,
            in2 => \_gnd_net_\,
            in3 => \N__16211\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i8_1_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35640\,
            in1 => \N__28437\,
            in2 => \_gnd_net_\,
            in3 => \N__18236\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i156_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35478\,
            in1 => \N__15173\,
            in2 => \_gnd_net_\,
            in3 => \N__15735\,
            lcout => data_in_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i132_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33246\,
            in1 => \N__32024\,
            in2 => \N__15207\,
            in3 => \N__16371\,
            lcout => \c0.data_in_field_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__19443\,
            in1 => \N__20360\,
            in2 => \N__15177\,
            in3 => \N__17769\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i146_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35477\,
            in1 => \N__15147\,
            in2 => \_gnd_net_\,
            in3 => \N__26726\,
            lcout => data_in_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16335\,
            in1 => \N__18286\,
            in2 => \_gnd_net_\,
            in3 => \N__35450\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i100_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35449\,
            in1 => \N__26333\,
            in2 => \_gnd_net_\,
            in3 => \N__16444\,
            lcout => data_in_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i122_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__28169\,
            in1 => \N__33006\,
            in2 => \N__19529\,
            in3 => \N__31849\,
            lcout => \c0.data_in_field_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5670_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27745\,
            in1 => \N__15265\,
            in2 => \N__30204\,
            in3 => \N__30529\,
            lcout => OPEN,
            ltout => \c0.n6009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6009_bdd_4_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__16598\,
            in1 => \N__15314\,
            in2 => \N__15330\,
            in3 => \N__30170\,
            lcout => \c0.n6012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i7_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31915\,
            in1 => \N__18219\,
            in2 => \N__33155\,
            in3 => \N__16645\,
            lcout => \c0.data_in_field_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_922_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28168\,
            in1 => \N__15313\,
            in2 => \N__30967\,
            in3 => \N__22949\,
            lcout => \c0.n2080\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i69_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__33253\,
            in1 => \N__23457\,
            in2 => \N__32283\,
            in3 => \N__15676\,
            lcout => \c0.data_in_field_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i9_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__15290\,
            in1 => \N__33254\,
            in2 => \N__32282\,
            in3 => \N__18252\,
            lcout => \c0.data_in_field_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_953_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15675\,
            in2 => \_gnd_net_\,
            in3 => \N__15289\,
            lcout => \c0.n2039\,
            ltout => \c0.n2039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_954_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15411\,
            in1 => \N__16587\,
            in2 => \N__15270\,
            in3 => \N__15261\,
            lcout => \c0.n5458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i54_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33252\,
            in1 => \N__32207\,
            in2 => \N__21051\,
            in3 => \N__15412\,
            lcout => \c0.data_in_field_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_945_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21975\,
            in1 => \N__15552\,
            in2 => \N__15516\,
            in3 => \N__20857\,
            lcout => \c0.n1835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_989_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25568\,
            in1 => \N__24942\,
            in2 => \N__30821\,
            in3 => \N__15341\,
            lcout => \c0.n41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5834_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__15414\,
            in1 => \N__27720\,
            in2 => \N__30153\,
            in3 => \N__22363\,
            lcout => \c0.n6213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15458\,
            in1 => \N__15876\,
            in2 => \_gnd_net_\,
            in3 => \N__15360\,
            lcout => \c0.n28_adj_1955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24317\,
            in2 => \_gnd_net_\,
            in3 => \N__22202\,
            lcout => OPEN,
            ltout => \c0.n14_adj_1957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1003_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21391\,
            in1 => \N__16665\,
            in2 => \N__15417\,
            in3 => \N__15413\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1903_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_835_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15894\,
            in1 => \N__30735\,
            in2 => \N__15396\,
            in3 => \N__15393\,
            lcout => OPEN,
            ltout => \c0.n5589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__15636\,
            in1 => \N__15387\,
            in2 => \N__15381\,
            in3 => \N__24621\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_955_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19388\,
            in2 => \_gnd_net_\,
            in3 => \N__15359\,
            lcout => \c0.n1994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_971_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21699\,
            in1 => \N__20741\,
            in2 => \N__26675\,
            in3 => \N__20555\,
            lcout => \c0.n5557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_807_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29408\,
            in1 => \N__16982\,
            in2 => \N__16602\,
            in3 => \N__22896\,
            lcout => OPEN,
            ltout => \c0.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_837_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15653\,
            in1 => \N__15623\,
            in2 => \N__15639\,
            in3 => \N__16950\,
            lcout => \c0.n5574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_845_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18789\,
            in2 => \_gnd_net_\,
            in3 => \N__18877\,
            lcout => \c0.n5572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_860_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20847\,
            lcout => \c0.n2000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i152_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19791\,
            in1 => \N__35348\,
            in2 => \_gnd_net_\,
            in3 => \N__23136\,
            lcout => data_in_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i32_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__32239\,
            in2 => \N__32838\,
            in3 => \N__30522\,
            lcout => \c0.data_in_field_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i72_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32237\,
            in1 => \N__32639\,
            in2 => \N__30775\,
            in3 => \N__15612\,
            lcout => \c0.data_in_field_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i138_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32637\,
            in1 => \N__32238\,
            in2 => \N__15582\,
            in3 => \N__30881\,
            lcout => \c0.data_in_field_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1006_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21178\,
            in1 => \N__28126\,
            in2 => \N__27260\,
            in3 => \N__15758\,
            lcout => OPEN,
            ltout => \c0.n18_adj_1959_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1008_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22712\,
            in1 => \N__15736\,
            in2 => \N__15714\,
            in3 => \N__19101\,
            lcout => OPEN,
            ltout => \c0.n20_adj_1870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19323\,
            in1 => \N__15711\,
            in2 => \N__15702\,
            in3 => \N__17394\,
            lcout => \c0.n5577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i125_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32236\,
            in1 => \N__32638\,
            in2 => \N__30324\,
            in3 => \N__21537\,
            lcout => \c0.data_in_field_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i42_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__16867\,
            in1 => \N__22452\,
            in2 => \N__32987\,
            in3 => \N__32292\,
            lcout => \c0.data_in_field_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i13_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__32290\,
            in1 => \N__23062\,
            in2 => \N__21765\,
            in3 => \N__32773\,
            lcout => \c0.data_in_field_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i103_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32769\,
            in1 => \N__32291\,
            in2 => \N__17793\,
            in3 => \N__17504\,
            lcout => \c0.data_in_field_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21527\,
            in1 => \N__17500\,
            in2 => \N__16868\,
            in3 => \N__21743\,
            lcout => \c0.n2101\,
            ltout => \c0.n2101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_901_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28306\,
            in1 => \N__24868\,
            in2 => \N__15693\,
            in3 => \N__26801\,
            lcout => OPEN,
            ltout => \c0.n6_adj_1917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_848_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17211\,
            in1 => \N__28020\,
            in2 => \N__15690\,
            in3 => \N__15683\,
            lcout => \c0.n5512\,
            ltout => \c0.n5512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_808_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17318\,
            in1 => \N__19074\,
            in2 => \N__15885\,
            in3 => \N__19557\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_929_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17499\,
            lcout => \c0.n2026\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_924_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15943\,
            in2 => \_gnd_net_\,
            in3 => \N__17124\,
            lcout => \c0.n2155\,
            ltout => \c0.n2155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16545\,
            in1 => \N__19589\,
            in2 => \N__15861\,
            in3 => \N__15792\,
            lcout => \c0.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i18_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__18290\,
            in1 => \N__32295\,
            in2 => \N__33068\,
            in3 => \N__15944\,
            lcout => \c0.data_in_field_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_991_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22763\,
            in1 => \N__15833\,
            in2 => \N__15984\,
            in3 => \N__29382\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i130_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32839\,
            in1 => \N__32294\,
            in2 => \N__15822\,
            in3 => \N__17125\,
            lcout => \c0.data_in_field_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i159_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15981\,
            in1 => \N__35347\,
            in2 => \_gnd_net_\,
            in3 => \N__16032\,
            lcout => data_in_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_903_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15791\,
            in1 => \N__17588\,
            in2 => \N__17353\,
            in3 => \N__15773\,
            lcout => \c0.n5491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i151_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15982\,
            in1 => \N__35346\,
            in2 => \_gnd_net_\,
            in3 => \N__16138\,
            lcout => data_in_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i113_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32587\,
            in1 => \N__32286\,
            in2 => \N__19695\,
            in3 => \N__17373\,
            lcout => \c0.data_in_field_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i153_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32285\,
            in1 => \N__32588\,
            in2 => \N__15963\,
            in3 => \N__21910\,
            lcout => \c0.data_in_frame_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i158_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35343\,
            in1 => \N__16047\,
            in2 => \_gnd_net_\,
            in3 => \N__19714\,
            lcout => data_in_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5739_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__27664\,
            in1 => \N__30016\,
            in2 => \N__30845\,
            in3 => \N__15945\,
            lcout => OPEN,
            ltout => \c0.n6093_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6093_bdd_4_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30017\,
            in1 => \N__30975\,
            in2 => \N__15930\,
            in3 => \N__18432\,
            lcout => \c0.n5767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i97_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25756\,
            in1 => \N__35345\,
            in2 => \_gnd_net_\,
            in3 => \N__19670\,
            lcout => data_in_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i131_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35342\,
            in1 => \N__25691\,
            in2 => \_gnd_net_\,
            in3 => \N__15907\,
            lcout => data_in_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20249\,
            in1 => \N__35344\,
            in2 => \_gnd_net_\,
            in3 => \N__27795\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i151_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__16109\,
            in1 => \N__32296\,
            in2 => \N__16146\,
            in3 => \N__32590\,
            lcout => \c0.data_in_frame_18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i152_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32589\,
            in1 => \N__16094\,
            in2 => \N__23156\,
            in3 => \N__32304\,
            lcout => \c0.data_in_frame_18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i50_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36047\,
            in1 => \N__16079\,
            in2 => \_gnd_net_\,
            in3 => \N__22463\,
            lcout => data_in_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_791_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20404\,
            in2 => \_gnd_net_\,
            in3 => \N__19951\,
            lcout => n1764,
            ltout => \n1764_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__20344\,
            in1 => \N__16043\,
            in2 => \N__16050\,
            in3 => \N__15990\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5854_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27613\,
            in1 => \N__18790\,
            in2 => \N__30093\,
            in3 => \N__18828\,
            lcout => \c0.n6237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__20093\,
            in1 => \N__18057\,
            in2 => \N__20361\,
            in3 => \N__16028\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16224\,
            in1 => \N__16010\,
            in2 => \_gnd_net_\,
            in3 => \N__16017\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_26_i4_2_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20004\,
            lcout => n4_adj_1980,
            ltout => \n4_adj_1980_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__16236\,
            in1 => \N__20345\,
            in2 => \N__16239\,
            in3 => \N__20092\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i157_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35349\,
            in1 => \N__16235\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => data_in_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5287_3_lut_4_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__17638\,
            in1 => \N__16307\,
            in2 => \N__18017\,
            in3 => \N__17690\,
            lcout => \c0.rx.n5633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_3_lut_4_lut_4_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001111"
        )
    port map (
            in0 => \N__17637\,
            in1 => \N__16306\,
            in2 => \N__18018\,
            in3 => \N__17689\,
            lcout => OPEN,
            ltout => \n2198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__16308\,
            in1 => \N__35261\,
            in2 => \N__16227\,
            in3 => \N__18003\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16223\,
            in1 => \N__16173\,
            in2 => \_gnd_net_\,
            in3 => \N__16179\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i87_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35255\,
            in1 => \N__19043\,
            in2 => \_gnd_net_\,
            in3 => \N__17461\,
            lcout => data_in_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_4_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__16295\,
            in1 => \N__17684\,
            in2 => \N__18006\,
            in3 => \N__17635\,
            lcout => \c0.rx.n2259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.n6291_bdd_4_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__16155\,
            in1 => \N__17983\,
            in2 => \N__20359\,
            in3 => \N__17598\,
            lcout => OPEN,
            ltout => \c0.rx.n6294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__16296\,
            in1 => \_gnd_net_\,
            in2 => \N__16311\,
            in3 => \_gnd_net_\,
            lcout => \r_SM_Main_0_adj_1991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__16294\,
            in1 => \N__17683\,
            in2 => \N__18005\,
            in3 => \N__17634\,
            lcout => \c0.rx.n1706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i90_2_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__17636\,
            in1 => \_gnd_net_\,
            in2 => \N__17696\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.rx.n75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__16297\,
            in1 => \N__18004\,
            in2 => \N__16251\,
            in3 => \N__16248\,
            lcout => \r_SM_Main_1_adj_1990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33570\,
            in1 => \N__23862\,
            in2 => \_gnd_net_\,
            in3 => \N__21638\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20043\,
            in1 => \N__20417\,
            in2 => \_gnd_net_\,
            in3 => \N__19999\,
            lcout => \c0.rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37581\,
            ce => \N__17927\,
            sr => \N__17898\
        );

    \c0.data_in_0___i67_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35634\,
            in1 => \N__23897\,
            in2 => \_gnd_net_\,
            in3 => \N__16729\,
            lcout => data_in_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i36_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35633\,
            in1 => \N__22108\,
            in2 => \_gnd_net_\,
            in3 => \N__16713\,
            lcout => data_in_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_886_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16488\,
            in1 => \N__18235\,
            in2 => \N__23069\,
            in3 => \N__22055\,
            lcout => \c0.n25_adj_1929\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35632\,
            in1 => \N__21101\,
            in2 => \_gnd_net_\,
            in3 => \N__16489\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16490\,
            in1 => \N__35635\,
            in2 => \_gnd_net_\,
            in3 => \N__18329\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i52_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33268\,
            in1 => \N__31715\,
            in2 => \N__16473\,
            in3 => \N__18726\,
            lcout => \c0.data_in_field_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i92_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35827\,
            in1 => \N__16933\,
            in2 => \_gnd_net_\,
            in3 => \N__16445\,
            lcout => data_in_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16565\,
            in1 => \N__16330\,
            in2 => \_gnd_net_\,
            in3 => \N__35829\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i100_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__31714\,
            in2 => \N__17209\,
            in3 => \N__16446\,
            lcout => \c0.data_in_field_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18509\,
            in1 => \N__23070\,
            in2 => \_gnd_net_\,
            in3 => \N__35828\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35826\,
            in1 => \N__17869\,
            in2 => \_gnd_net_\,
            in3 => \N__25045\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_885_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18508\,
            in1 => \N__16329\,
            in2 => \N__16431\,
            in3 => \N__16561\,
            lcout => \c0.n27_adj_1928\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_985_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20164\,
            in1 => \N__19639\,
            in2 => \N__19790\,
            in3 => \N__16362\,
            lcout => \c0.n22_adj_1886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i10_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31705\,
            in1 => \N__16331\,
            in2 => \N__18423\,
            in3 => \N__33163\,
            lcout => \c0.data_in_field_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i8_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__18105\,
            in1 => \N__31709\,
            in2 => \N__33242\,
            in3 => \N__16594\,
            lcout => \c0.data_in_field_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i2_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31706\,
            in1 => \N__33159\,
            in2 => \N__16566\,
            in3 => \N__30966\,
            lcout => \c0.data_in_field_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i6_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31707\,
            in1 => \N__20211\,
            in2 => \N__22823\,
            in3 => \N__33164\,
            lcout => \c0.data_in_field_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i108_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33158\,
            in1 => \N__31708\,
            in2 => \N__26337\,
            in3 => \N__22959\,
            lcout => \c0.data_in_field_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18186\,
            in1 => \N__35830\,
            in2 => \_gnd_net_\,
            in3 => \N__31443\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i22_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31710\,
            in1 => \N__33086\,
            in2 => \N__17877\,
            in3 => \N__27131\,
            lcout => \c0.data_in_field_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_967_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22813\,
            in1 => \_gnd_net_\,
            in2 => \N__21798\,
            in3 => \N__17154\,
            lcout => \c0.n2104\,
            ltout => \c0.n2104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_871_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16533\,
            in1 => \N__16611\,
            in2 => \N__16527\,
            in3 => \N__20688\,
            lcout => \c0.n5497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i66_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33085\,
            in1 => \N__31712\,
            in2 => \N__16524\,
            in3 => \N__17155\,
            lcout => \c0.data_in_field_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i81_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31711\,
            in1 => \N__33087\,
            in2 => \N__21982\,
            in3 => \N__30452\,
            lcout => \c0.data_in_field_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_966_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22812\,
            in1 => \N__17153\,
            in2 => \N__27137\,
            in3 => \N__16617\,
            lcout => \c0.n5521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_896_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__17311\,
            in1 => \N__18464\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n5476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1002_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18585\,
            in1 => \N__20740\,
            in2 => \N__26645\,
            in3 => \N__22544\,
            lcout => \c0.n20_adj_1958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16767\,
            in1 => \N__26611\,
            in2 => \N__21227\,
            in3 => \N__24437\,
            lcout => OPEN,
            ltout => \c0.n31_adj_1896_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_829_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21693\,
            in1 => \N__22350\,
            in2 => \N__16659\,
            in3 => \N__16656\,
            lcout => \c0.n47_adj_1897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_843_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16646\,
            in1 => \N__20516\,
            in2 => \N__19021\,
            in3 => \N__24707\,
            lcout => \c0.n10_adj_1915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i110_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__26612\,
            in1 => \N__32763\,
            in2 => \N__34491\,
            in3 => \N__31887\,
            lcout => \c0.data_in_field_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i126_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31882\,
            in1 => \N__21309\,
            in2 => \N__32986\,
            in3 => \N__17310\,
            lcout => \c0.data_in_field_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_944_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17309\,
            in1 => \N__18470\,
            in2 => \_gnd_net_\,
            in3 => \N__16766\,
            lcout => \c0.n1913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i65_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__32762\,
            in1 => \N__16788\,
            in2 => \N__32100\,
            in3 => \N__31062\,
            lcout => \c0.data_in_field_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i136_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__22425\,
            in1 => \N__31883\,
            in2 => \N__17283\,
            in3 => \N__32767\,
            lcout => \c0.data_in_field_135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i11_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__22020\,
            in1 => \N__32054\,
            in2 => \N__33276\,
            in3 => \N__16897\,
            lcout => \c0.data_in_field_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i67_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32053\,
            in1 => \N__33263\,
            in2 => \N__16743\,
            in3 => \N__20950\,
            lcout => \c0.data_in_field_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i141_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33261\,
            in1 => \N__32055\,
            in2 => \N__27395\,
            in3 => \N__18881\,
            lcout => \c0.data_in_field_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i44_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32052\,
            in1 => \N__33262\,
            in2 => \N__16712\,
            in3 => \N__19106\,
            lcout => \c0.data_in_field_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5839_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27686\,
            in1 => \N__19338\,
            in2 => \N__30149\,
            in3 => \N__27133\,
            lcout => \c0.n6219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5809_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__22650\,
            in1 => \N__27687\,
            in2 => \N__19164\,
            in3 => \N__30065\,
            lcout => \c0.n6183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_936_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30607\,
            in2 => \_gnd_net_\,
            in3 => \N__27132\,
            lcout => OPEN,
            ltout => \c0.n2062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19260\,
            in1 => \N__18823\,
            in2 => \N__17046\,
            in3 => \N__18624\,
            lcout => \c0.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24746\,
            in1 => \N__17027\,
            in2 => \N__18958\,
            in3 => \N__16836\,
            lcout => \c0.n5503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16911\,
            in1 => \N__16971\,
            in2 => \N__24180\,
            in3 => \N__17237\,
            lcout => \c0.n16_adj_1871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i92_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32089\,
            in1 => \N__16943\,
            in2 => \N__33275\,
            in3 => \N__27951\,
            lcout => \c0.data_in_field_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_863_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20943\,
            in2 => \_gnd_net_\,
            in3 => \N__19159\,
            lcout => \c0.n2021\,
            ltout => \c0.n2021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_864_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16890\,
            in1 => \N__16812\,
            in2 => \N__16872\,
            in3 => \N__26800\,
            lcout => \c0.n2074\,
            ltout => \c0.n2074_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_976_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16860\,
            in1 => \N__22742\,
            in2 => \N__16839\,
            in3 => \N__16835\,
            lcout => \c0.n5527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i27_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32088\,
            in1 => \N__21486\,
            in2 => \N__33274\,
            in3 => \N__16813\,
            lcout => \c0.data_in_field_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i134_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18694\,
            in1 => \N__21347\,
            in2 => \_gnd_net_\,
            in3 => \N__35965\,
            lcout => data_in_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19070\,
            in1 => \N__27210\,
            in2 => \N__17409\,
            in3 => \N__17379\,
            lcout => \c0.n48_adj_1895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_923_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__19207\,
            in2 => \N__19469\,
            in3 => \N__17273\,
            lcout => \c0.n5418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i75_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32293\,
            in1 => \N__32768\,
            in2 => \N__23910\,
            in3 => \N__31000\,
            lcout => \c0.data_in_field_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_898_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27941\,
            in2 => \_gnd_net_\,
            in3 => \N__19461\,
            lcout => \c0.n1908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_919_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17441\,
            in1 => \N__17210\,
            in2 => \N__30768\,
            in3 => \N__24581\,
            lcout => \c0.n1889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i126_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35964\,
            in1 => \N__18695\,
            in2 => \_gnd_net_\,
            in3 => \N__21289\,
            lcout => data_in_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i127_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18813\,
            in1 => \N__17730\,
            in2 => \N__32222\,
            in3 => \N__32602\,
            lcout => \c0.data_in_field_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_910_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25947\,
            in1 => \N__17162\,
            in2 => \_gnd_net_\,
            in3 => \N__17126\,
            lcout => \c0.n5569\,
            ltout => \c0.n5569_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25727\,
            in2 => \N__17094\,
            in3 => \N__17091\,
            lcout => \c0.n20_adj_1882\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_908_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19232\,
            in1 => \N__30993\,
            in2 => \N__23013\,
            in3 => \N__17565\,
            lcout => \c0.n1958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_938_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17566\,
            in1 => \N__23003\,
            in2 => \_gnd_net_\,
            in3 => \N__19233\,
            lcout => \c0.n5388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i79_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__19234\,
            in1 => \N__31193\,
            in2 => \N__32780\,
            in3 => \N__32099\,
            lcout => \c0.data_in_field_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_adj_988_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17400\,
            in1 => \N__19245\,
            in2 => \N__22895\,
            in3 => \N__17390\,
            lcout => \c0.n44_adj_1894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_881_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17371\,
            in1 => \N__18812\,
            in2 => \_gnd_net_\,
            in3 => \N__17564\,
            lcout => \c0.n5524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_926_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17346\,
            in2 => \_gnd_net_\,
            in3 => \N__17435\,
            lcout => \c0.n1917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i160_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19789\,
            in1 => \N__17748\,
            in2 => \_gnd_net_\,
            in3 => \N__36046\,
            lcout => data_in_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i31_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32847\,
            in1 => \N__32288\,
            in2 => \N__17355\,
            in3 => \N__20250\,
            lcout => \c0.data_in_field_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5824_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27663\,
            in1 => \N__22206\,
            in2 => \N__30112\,
            in3 => \N__17322\,
            lcout => \c0.n6201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_986_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22674\,
            in1 => \N__19553\,
            in2 => \N__30264\,
            in3 => \N__17592\,
            lcout => \c0.n18_adj_1887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i77_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__32287\,
            in1 => \N__30390\,
            in2 => \N__17576\,
            in3 => \N__32846\,
            lcout => \c0.data_in_field_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i149_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__17543\,
            in1 => \N__20123\,
            in2 => \N__33069\,
            in3 => \N__32289\,
            lcout => \c0.data_in_frame_18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i141_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20122\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__27379\,
            lcout => data_in_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5859_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27685\,
            in1 => \N__21003\,
            in2 => \N__30184\,
            in3 => \N__17439\,
            lcout => OPEN,
            ltout => \c0.n6243_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6243_bdd_4_lut_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__29513\,
            in1 => \N__19239\,
            in2 => \N__17529\,
            in3 => \N__30125\,
            lcout => OPEN,
            ltout => \c0.n5698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5869_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__25402\,
            in1 => \N__25252\,
            in2 => \N__17526\,
            in3 => \N__17481\,
            lcout => \c0.n6231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6237_bdd_4_lut_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__23691\,
            in2 => \N__17508\,
            in3 => \N__30121\,
            lcout => \c0.n5701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i87_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__17440\,
            in1 => \N__17475\,
            in2 => \N__32303\,
            in3 => \N__32591\,
            lcout => \c0.data_in_field_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i82_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21248\,
            in1 => \_gnd_net_\,
            in2 => \N__35684\,
            in3 => \N__17837\,
            lcout => data_in_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i74_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17836\,
            in1 => \N__35511\,
            in2 => \_gnd_net_\,
            in3 => \N__17804\,
            lcout => data_in_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i95_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__19042\,
            in2 => \_gnd_net_\,
            in3 => \N__17783\,
            lcout => data_in_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i103_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35259\,
            in1 => \N__22915\,
            in2 => \_gnd_net_\,
            in3 => \N__17782\,
            lcout => data_in_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__20349\,
            in2 => \N__17747\,
            in3 => \N__17759\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_27_i4_2_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20045\,
            in2 => \_gnd_net_\,
            in3 => \N__20000\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i119_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35257\,
            in1 => \N__19807\,
            in2 => \_gnd_net_\,
            in3 => \N__17726\,
            lcout => data_in_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i98_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19406\,
            in1 => \N__35258\,
            in2 => \_gnd_net_\,
            in3 => \N__19897\,
            lcout => data_in_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i106_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35256\,
            in1 => \N__19499\,
            in2 => \_gnd_net_\,
            in3 => \N__19405\,
            lcout => data_in_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000111100"
        )
    port map (
            in0 => \N__18035\,
            in1 => \N__17688\,
            in2 => \N__18016\,
            in3 => \N__17646\,
            lcout => \c0.rx.n6291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100110001000"
        )
    port map (
            in0 => \N__20411\,
            in1 => \N__18063\,
            in2 => \N__18039\,
            in3 => \N__17996\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i90_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35448\,
            in1 => \N__21241\,
            in2 => \_gnd_net_\,
            in3 => \N__19898\,
            lcout => data_in_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3393_2_lut_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20033\,
            lcout => n3636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_3_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20032\,
            in1 => \N__20402\,
            in2 => \_gnd_net_\,
            in3 => \N__19989\,
            lcout => \c0.rx.n3850\,
            ltout => \c0.rx.n3850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2116_2_lut_3_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17992\,
            in2 => \N__17931\,
            in3 => \N__17914\,
            lcout => \c0.rx.n2367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20416\,
            in2 => \_gnd_net_\,
            in3 => \N__19998\,
            lcout => \c0.rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37590\,
            ce => \N__17928\,
            sr => \N__17897\
        );

    \c0.i10_4_lut_adj_882_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18328\,
            in1 => \N__21099\,
            in2 => \N__17870\,
            in3 => \N__28432\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21100\,
            in1 => \N__35636\,
            in2 => \_gnd_net_\,
            in3 => \N__22087\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__27896\,
            in2 => \N__35825\,
            in3 => \_gnd_net_\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_877_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18211\,
            in1 => \N__25044\,
            in2 => \N__18104\,
            in3 => \N__18134\,
            lcout => OPEN,
            ltout => \c0.n28_adj_1926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_956_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18312\,
            in1 => \N__18306\,
            in2 => \N__18300\,
            in3 => \N__18297\,
            lcout => \c0.n4795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35928\,
            in1 => \N__18152\,
            in2 => \_gnd_net_\,
            in3 => \N__27819\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_925_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20236\,
            in1 => \N__20184\,
            in2 => \N__18291\,
            in3 => \N__27771\,
            lcout => \c0.n30_adj_1941\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35931\,
            in1 => \N__22264\,
            in2 => \_gnd_net_\,
            in3 => \N__18248\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18151\,
            in1 => \N__35929\,
            in2 => \_gnd_net_\,
            in3 => \N__18212\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_912_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18193\,
            in1 => \N__18150\,
            in2 => \N__24680\,
            in3 => \N__22309\,
            lcout => \c0.n26_adj_1940\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18135\,
            in1 => \N__35930\,
            in2 => \_gnd_net_\,
            in3 => \N__18100\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_958_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__18084\,
            in1 => \N__18078\,
            in2 => \N__18072\,
            in3 => \N__21015\,
            lcout => \c0.n1729\,
            ltout => \c0.n1729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i36_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__22116\,
            in1 => \N__33165\,
            in2 => \N__18474\,
            in3 => \N__18465\,
            lcout => \c0.data_in_field_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i28_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__22092\,
            in1 => \N__31700\,
            in2 => \N__33243\,
            in3 => \N__18605\,
            lcout => \c0.data_in_field_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i55_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18358\,
            in1 => \N__24209\,
            in2 => \N__31944\,
            in3 => \N__33173\,
            lcout => \c0.data_in_field_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_934_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18718\,
            lcout => OPEN,
            ltout => \c0.n5369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_935_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18357\,
            in1 => \N__18914\,
            in2 => \N__18339\,
            in3 => \N__26828\,
            lcout => \c0.n2125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i33_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__26829\,
            in1 => \N__23496\,
            in2 => \N__33244\,
            in3 => \N__31704\,
            lcout => \c0.data_in_field_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i4_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31699\,
            in1 => \N__33166\,
            in2 => \N__18336\,
            in3 => \N__18646\,
            lcout => \c0.data_in_field_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i56_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21070\,
            in1 => \N__35927\,
            in2 => \_gnd_net_\,
            in3 => \N__23267\,
            lcout => data_in_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35926\,
            in1 => \N__24670\,
            in2 => \_gnd_net_\,
            in3 => \N__22019\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i76_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33084\,
            in1 => \N__31713\,
            in2 => \N__18681\,
            in3 => \N__19020\,
            lcout => \c0.data_in_field_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_869_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18640\,
            in2 => \_gnd_net_\,
            in3 => \N__18620\,
            lcout => \c0.n6_adj_1923\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_867_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18601\,
            in2 => \_gnd_net_\,
            in3 => \N__20471\,
            lcout => \c0.n5469\,
            ltout => \c0.n5469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_870_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18573\,
            in1 => \N__18540\,
            in2 => \N__18525\,
            in3 => \N__18522\,
            lcout => \c0.n5548\,
            ltout => \c0.n5548_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22691\,
            in1 => \N__20495\,
            in2 => \N__18516\,
            in3 => \N__24401\,
            lcout => \c0.n45_adj_1892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i5_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__18513\,
            in1 => \N__32059\,
            in2 => \N__33233\,
            in3 => \N__21797\,
            lcout => \c0.data_in_field_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i62_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32056\,
            in1 => \N__33131\,
            in2 => \N__18495\,
            in3 => \N__22346\,
            lcout => \c0.data_in_field_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i116_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33129\,
            in1 => \N__32057\,
            in2 => \N__26373\,
            in3 => \N__20613\,
            lcout => \c0.data_in_field_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i34_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18910\,
            in1 => \N__23181\,
            in2 => \N__32216\,
            in3 => \N__33135\,
            lcout => \c0.data_in_field_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_893_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19190\,
            in1 => \N__18909\,
            in2 => \_gnd_net_\,
            in3 => \N__27952\,
            lcout => \c0.n5403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_892_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18876\,
            in2 => \_gnd_net_\,
            in3 => \N__22345\,
            lcout => \c0.n5391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i41_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33130\,
            in1 => \N__32058\,
            in2 => \N__23523\,
            in3 => \N__26789\,
            lcout => \c0.data_in_field_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_982_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27084\,
            in1 => \N__28058\,
            in2 => \N__18962\,
            in3 => \N__28122\,
            lcout => \c0.n5539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i93_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33118\,
            in1 => \N__31932\,
            in2 => \N__24969\,
            in3 => \N__19191\,
            lcout => \c0.data_in_field_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i104_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__18855\,
            in1 => \N__19136\,
            in2 => \N__32132\,
            in3 => \N__33120\,
            lcout => \c0.data_in_field_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_820_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19116\,
            in1 => \N__18824\,
            in2 => \N__18792\,
            in3 => \N__18736\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22044\,
            in1 => \_gnd_net_\,
            in2 => \N__35963\,
            in3 => \N__21485\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i134_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33117\,
            in1 => \N__31931\,
            in2 => \N__18702\,
            in3 => \N__27157\,
            lcout => \c0.data_in_field_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i53_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31930\,
            in1 => \N__33119\,
            in2 => \N__23400\,
            in3 => \N__19163\,
            lcout => \c0.data_in_field_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_847_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19132\,
            in2 => \_gnd_net_\,
            in3 => \N__27156\,
            lcout => \c0.n2152\,
            ltout => \c0.n2152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_849_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23079\,
            in1 => \N__19105\,
            in2 => \N__19077\,
            in3 => \N__20739\,
            lcout => \c0.n5397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i30_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32090\,
            in1 => \N__19337\,
            in2 => \N__27900\,
            in3 => \N__32807\,
            lcout => \c0.data_in_field_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i95_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32805\,
            in1 => \N__32092\,
            in2 => \N__19053\,
            in3 => \N__21000\,
            lcout => \c0.data_in_field_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_905_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23339\,
            in1 => \N__23306\,
            in2 => \_gnd_net_\,
            in3 => \N__19022\,
            lcout => \c0.n2065\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i143_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32804\,
            in1 => \N__32091\,
            in2 => \N__18990\,
            in3 => \N__18945\,
            lcout => \c0.data_in_field_142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i144_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__27071\,
            in1 => \N__23109\,
            in2 => \N__32221\,
            in3 => \N__32806\,
            lcout => \c0.data_in_field_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_field_143__I_0_1808_2_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18944\,
            in2 => \_gnd_net_\,
            in3 => \N__27070\,
            lcout => OPEN,
            ltout => \c0.tx2_transmit_N_1031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_927_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20163\,
            in1 => \N__25144\,
            in2 => \N__19341\,
            in3 => \N__19336\,
            lcout => \c0.n2030\,
            ltout => \c0.n2030_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20576\,
            in1 => \N__22235\,
            in2 => \N__19314\,
            in3 => \N__22649\,
            lcout => \c0.n5466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i23_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__19274\,
            in2 => \N__27815\,
            in3 => \N__33124\,
            lcout => \c0.data_in_field_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i123_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__33121\,
            in1 => \N__32086\,
            in2 => \N__24603\,
            in3 => \N__19311\,
            lcout => \c0.data_in_field_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i83_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32085\,
            in1 => \N__33123\,
            in2 => \N__30678\,
            in3 => \N__19582\,
            lcout => \c0.data_in_field_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_914_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19273\,
            in1 => \N__19616\,
            in2 => \_gnd_net_\,
            in3 => \N__20977\,
            lcout => \c0.n5436\,
            ltout => \c0.n5436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_900_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19549\,
            in2 => \N__19248\,
            in3 => \N__21440\,
            lcout => \c0.n5509\,
            ltout => \c0.n5509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_874_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19235\,
            in2 => \N__19212\,
            in3 => \N__19208\,
            lcout => \c0.n2053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_918_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__20978\,
            in1 => \_gnd_net_\,
            in2 => \N__21568\,
            in3 => \_gnd_net_\,
            lcout => \c0.n1779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i37_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33122\,
            in1 => \N__32087\,
            in2 => \N__31230\,
            in3 => \N__19617\,
            lcout => \c0.data_in_field_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i117_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31936\,
            in1 => \N__32760\,
            in2 => \N__21572\,
            in3 => \N__26925\,
            lcout => \c0.data_in_field_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_917_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19575\,
            in1 => \N__19860\,
            in2 => \_gnd_net_\,
            in3 => \N__20780\,
            lcout => \c0.n1948\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i114_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35812\,
            in1 => \N__19486\,
            in2 => \_gnd_net_\,
            in3 => \N__19533\,
            lcout => data_in_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i19_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31937\,
            in1 => \N__22054\,
            in2 => \N__23020\,
            in3 => \N__32761\,
            lcout => \c0.data_in_field_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i128_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32759\,
            in1 => \N__31939\,
            in2 => \N__21876\,
            in3 => \N__19468\,
            lcout => \c0.data_in_field_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__19439\,
            in1 => \N__20364\,
            in2 => \N__25496\,
            in3 => \N__20094\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i106_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__31938\,
            in2 => \N__19416\,
            in3 => \N__19376\,
            lcout => \c0.data_in_field_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_824_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19362\,
            in1 => \N__27326\,
            in2 => \N__20124\,
            in3 => \N__25464\,
            lcout => \c0.n20_adj_1888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i98_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31940\,
            in1 => \N__32970\,
            in2 => \N__19905\,
            in3 => \N__19869\,
            lcout => \c0.data_in_field_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i153_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21895\,
            in1 => \N__19923\,
            in2 => \_gnd_net_\,
            in3 => \N__35516\,
            lcout => data_in_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i113_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35515\,
            in1 => \N__19687\,
            in2 => \_gnd_net_\,
            in3 => \N__35069\,
            lcout => data_in_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i97_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32969\,
            in1 => \N__31941\,
            in2 => \N__20802\,
            in3 => \N__25760\,
            lcout => \c0.data_in_field_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i158_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__19832\,
            in1 => \N__19730\,
            in2 => \N__33136\,
            in3 => \N__31943\,
            lcout => \c0.data_in_frame_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i111_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35629\,
            in1 => \N__19814\,
            in2 => \_gnd_net_\,
            in3 => \N__22916\,
            lcout => data_in_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i160_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__19745\,
            in1 => \N__31942\,
            in2 => \N__33137\,
            in3 => \N__19782\,
            lcout => \c0.data_in_frame_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i150_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35518\,
            in1 => \N__21381\,
            in2 => \_gnd_net_\,
            in3 => \N__19729\,
            lcout => data_in_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i105_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35628\,
            in1 => \N__19688\,
            in2 => \_gnd_net_\,
            in3 => \N__19657\,
            lcout => data_in_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__29200\,
            in1 => \N__29115\,
            in2 => \N__29022\,
            in3 => \N__28495\,
            lcout => \c0.tx.n2247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i149_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35517\,
            in1 => \N__20118\,
            in2 => \_gnd_net_\,
            in3 => \N__20653\,
            lcout => data_in_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33868\,
            in2 => \_gnd_net_\,
            in3 => \N__29238\,
            lcout => OPEN,
            ltout => \c0.tx.n40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2105_4_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__29116\,
            in1 => \N__20066\,
            in2 => \N__20097\,
            in3 => \N__29327\,
            lcout => \c0.tx.n2356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_792_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19956\,
            lcout => n1760,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__29334\,
            in1 => \_gnd_net_\,
            in2 => \N__33884\,
            in3 => \N__29239\,
            lcout => \c0.tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => \N__20073\,
            sr => \N__20055\
        );

    \c0.tx.r_Bit_Index_i1_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33869\,
            in2 => \_gnd_net_\,
            in3 => \N__29333\,
            lcout => \c0.tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37582\,
            ce => \N__20073\,
            sr => \N__20055\
        );

    \c0.tx.i1_2_lut_3_lut_4_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__29005\,
            in1 => \N__29203\,
            in2 => \N__28617\,
            in3 => \N__29121\,
            lcout => n1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20049\,
            in1 => \N__19997\,
            in2 => \_gnd_net_\,
            in3 => \N__19952\,
            lcout => n1757,
            ltout => \n1757_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__19916\,
            in1 => \N__20412\,
            in2 => \N__19926\,
            in3 => \N__20363\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20418\,
            in1 => \N__20362\,
            in2 => \N__26390\,
            in3 => \N__20256\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35557\,
            in1 => \N__25058\,
            in2 => \_gnd_net_\,
            in3 => \N__20201\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i47_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35406\,
            in1 => \N__24210\,
            in2 => \_gnd_net_\,
            in3 => \N__23353\,
            lcout => data_in_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30629\,
            in1 => \_gnd_net_\,
            in2 => \N__35558\,
            in3 => \N__20235\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i39_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23354\,
            in1 => \N__35405\,
            in2 => \_gnd_net_\,
            in3 => \N__30628\,
            lcout => data_in_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20200\,
            in2 => \_gnd_net_\,
            in3 => \N__22005\,
            lcout => \c0.n22_adj_1924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i63_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35407\,
            in1 => \N__31170\,
            in2 => \_gnd_net_\,
            in3 => \N__24226\,
            lcout => data_in_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i142_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32122\,
            in1 => \N__33157\,
            in2 => \N__21354\,
            in3 => \N__20150\,
            lcout => \c0.data_in_field_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_928_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22637\,
            lcout => \c0.n5590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_949_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28299\,
            in2 => \_gnd_net_\,
            in3 => \N__24861\,
            lcout => OPEN,
            ltout => \c0.n5394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_825_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29445\,
            in1 => \N__20499\,
            in2 => \N__20478\,
            in3 => \N__20475\,
            lcout => \c0.n19_adj_1889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_821_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__22194\,
            in2 => \N__20430\,
            in3 => \N__22170\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i118_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33156\,
            in1 => \N__32123\,
            in2 => \N__31311\,
            in3 => \N__22195\,
            lcout => \c0.data_in_field_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i56_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33095\,
            in1 => \N__32205\,
            in2 => \N__21080\,
            in3 => \N__26986\,
            lcout => \c0.data_in_field_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i35_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32203\,
            in1 => \N__33097\,
            in2 => \N__21423\,
            in3 => \N__20543\,
            lcout => \c0.data_in_field_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i133_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33094\,
            in1 => \N__32204\,
            in2 => \N__30351\,
            in3 => \N__20714\,
            lcout => \c0.data_in_field_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_961_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30829\,
            in1 => \N__31416\,
            in2 => \N__26990\,
            in3 => \N__30892\,
            lcout => \c0.n5515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_828_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26982\,
            in1 => \N__23622\,
            in2 => \N__21915\,
            in3 => \N__21771\,
            lcout => OPEN,
            ltout => \c0.n40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20760\,
            in1 => \N__21267\,
            in2 => \N__20754\,
            in3 => \N__20751\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i61_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33096\,
            in1 => \N__32206\,
            in2 => \N__23427\,
            in3 => \N__22642\,
            lcout => \c0.data_in_field_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37516\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_861_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20713\,
            in1 => \N__21680\,
            in2 => \_gnd_net_\,
            in3 => \N__20542\,
            lcout => \c0.n1969\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_895_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24380\,
            in1 => \N__20675\,
            in2 => \_gnd_net_\,
            in3 => \N__25105\,
            lcout => \c0.n1855\,
            ltout => \c0.n1855_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_832_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20661\,
            in1 => \N__20615\,
            in2 => \N__20586\,
            in3 => \N__20583\,
            lcout => \c0.n13_adj_1899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i21_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__31104\,
            in1 => \N__32172\,
            in2 => \N__21698\,
            in3 => \N__33271\,
            lcout => \c0.data_in_field_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35853\,
            in1 => \N__23492\,
            in2 => \_gnd_net_\,
            in3 => \N__27843\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i69_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35401\,
            in1 => \N__30386\,
            in2 => \_gnd_net_\,
            in3 => \N__23449\,
            lcout => data_in_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_962_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22574\,
            in1 => \N__22529\,
            in2 => \N__25984\,
            in3 => \N__20541\,
            lcout => \c0.n2092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i140_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__22530\,
            in1 => \N__33270\,
            in2 => \N__21135\,
            in3 => \N__32173\,
            lcout => \c0.data_in_field_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i20_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__33269\,
            in1 => \N__22582\,
            in2 => \N__21111\,
            in3 => \N__32126\,
            lcout => \c0.data_in_field_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i48_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35904\,
            in1 => \N__21081\,
            in2 => \_gnd_net_\,
            in3 => \N__27181\,
            lcout => data_in_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i46_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35901\,
            in1 => \N__21044\,
            in2 => \_gnd_net_\,
            in3 => \N__22501\,
            lcout => data_in_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i45_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23396\,
            in1 => \N__35902\,
            in2 => \_gnd_net_\,
            in3 => \N__27343\,
            lcout => data_in_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_957_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22091\,
            in1 => \N__31102\,
            in2 => \N__22278\,
            in3 => \N__21478\,
            lcout => \c0.n25_adj_1948\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_911_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21002\,
            in1 => \N__20951\,
            in2 => \_gnd_net_\,
            in3 => \N__20923\,
            lcout => \c0.n5545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_979_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21273\,
            in1 => \N__22725\,
            in2 => \N__30734\,
            in3 => \N__23655\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_907_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20858\,
            in2 => \_gnd_net_\,
            in3 => \N__20810\,
            lcout => \c0.n5427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21809\,
            in1 => \N__21539\,
            in2 => \N__25455\,
            in3 => \N__28114\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i94_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__25104\,
            in1 => \N__32006\,
            in2 => \N__27021\,
            in3 => \N__32895\,
            lcout => \c0.data_in_field_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i118_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31297\,
            in1 => \N__35903\,
            in2 => \_gnd_net_\,
            in3 => \N__21308\,
            lcout => data_in_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_rep_100_2_lut_3_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__26642\,
            in2 => \_gnd_net_\,
            in3 => \N__21179\,
            lcout => \c0.n6414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_853_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21808\,
            in2 => \_gnd_net_\,
            in3 => \N__21538\,
            lcout => \c0.n5563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i46_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__21210\,
            in1 => \N__32894\,
            in2 => \N__22506\,
            in3 => \N__32007\,
            lcout => \c0.data_in_field_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i90_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32005\,
            in1 => \N__33227\,
            in2 => \N__21258\,
            in3 => \N__23338\,
            lcout => \c0.data_in_field_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_952_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21211\,
            in2 => \_gnd_net_\,
            in3 => \N__26643\,
            lcout => OPEN,
            ltout => \c0.n2149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21183\,
            in1 => \N__21156\,
            in2 => \N__21150\,
            in3 => \N__22608\,
            lcout => \c0.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36054\,
            in1 => \N__21413\,
            in2 => \_gnd_net_\,
            in3 => \N__21471\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_899_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25094\,
            in2 => \_gnd_net_\,
            in3 => \N__23221\,
            lcout => \c0.n1955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i35_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36055\,
            in1 => \N__21412\,
            in2 => \_gnd_net_\,
            in3 => \N__25628\,
            lcout => data_in_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i142_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36053\,
            in1 => \N__21340\,
            in2 => \_gnd_net_\,
            in3 => \N__21395\,
            lcout => data_in_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i0_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23549\,
            in2 => \N__36792\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \c0.n4754\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21597\,
            in2 => \_gnd_net_\,
            in3 => \N__21324\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n4754\,
            carryout => \c0.n4755\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i2_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23562\,
            in2 => \_gnd_net_\,
            in3 => \N__21321\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n4755\,
            carryout => \c0.n4756\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26099\,
            in2 => \_gnd_net_\,
            in3 => \N__21318\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n4756\,
            carryout => \c0.n4757\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i4_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26021\,
            in2 => \_gnd_net_\,
            in3 => \N__21315\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n4757\,
            carryout => \c0.n4758\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i5_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21585\,
            in2 => \_gnd_net_\,
            in3 => \N__21312\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n4758\,
            carryout => \c0.n4759\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i6_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26081\,
            in2 => \_gnd_net_\,
            in3 => \N__21612\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n4759\,
            carryout => \c0.n4760\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i7_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23535\,
            in2 => \_gnd_net_\,
            in3 => \N__21609\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \c0.n4760\,
            carryout => \c0.n4761\,
            clk => \N__37569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i8_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26039\,
            in2 => \_gnd_net_\,
            in3 => \N__21606\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \c0.n4762\,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i9_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23574\,
            in2 => \_gnd_net_\,
            in3 => \N__21603\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \c0.n4762\,
            carryout => \c0.n4763\,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_528__i10_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21600\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21584\,
            lcout => \c0.n16_adj_1921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5799_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27703\,
            in1 => \N__21573\,
            in2 => \N__30173\,
            in3 => \N__21543\,
            lcout => OPEN,
            ltout => \c0.n6171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6171_bdd_4_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30113\,
            in1 => \N__30260\,
            in2 => \N__21504\,
            in3 => \N__24869\,
            lcout => \c0.n5731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6189_bdd_4_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30100\,
            in1 => \N__21813\,
            in2 => \N__21657\,
            in3 => \N__21770\,
            lcout => \c0.n5722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i3388_2_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29017\,
            in2 => \_gnd_net_\,
            in3 => \N__29092\,
            lcout => OPEN,
            ltout => \c0.tx.n3631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5592_3_lut_4_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__28609\,
            in1 => \N__29173\,
            in2 => \N__21702\,
            in3 => \N__23807\,
            lcout => \c0.tx.n5883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23727\,
            in1 => \N__33605\,
            in2 => \_gnd_net_\,
            in3 => \N__21624\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i17_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__28725\,
            in1 => \N__23847\,
            in2 => \N__36183\,
            in3 => \N__37727\,
            lcout => data_out_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5819_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27612\,
            in1 => \N__28238\,
            in2 => \N__30174\,
            in3 => \N__21697\,
            lcout => \c0.n6189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5604_2_lut_3_lut_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__28477\,
            in1 => \_gnd_net_\,
            in2 => \N__29253\,
            in3 => \N__33888\,
            lcout => OPEN,
            ltout => \c0.tx.n5812_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i28_4_lut_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28613\,
            in1 => \N__29089\,
            in2 => \N__21648\,
            in3 => \N__29326\,
            lcout => OPEN,
            ltout => \c0.tx.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__28478\,
            in1 => \N__29016\,
            in2 => \N__21645\,
            in3 => \N__29175\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__21642\,
            in1 => \N__21623\,
            in2 => \N__33893\,
            in3 => \N__29325\,
            lcout => \c0.tx.n6285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26499\,
            in2 => \_gnd_net_\,
            in3 => \N__21840\,
            lcout => n321,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \c0.tx.n4764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26421\,
            in2 => \_gnd_net_\,
            in3 => \N__21837\,
            lcout => n320,
            ltout => OPEN,
            carryin => \c0.tx.n4764\,
            carryout => \c0.tx.n4765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22134\,
            in1 => \N__23977\,
            in2 => \_gnd_net_\,
            in3 => \N__21834\,
            lcout => \c0.tx.n5885\,
            ltout => OPEN,
            carryin => \c0.tx.n4765\,
            carryout => \c0.tx.n4766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26538\,
            in2 => \_gnd_net_\,
            in3 => \N__21831\,
            lcout => n318,
            ltout => OPEN,
            carryin => \c0.tx.n4766\,
            carryout => \c0.tx.n4767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24068\,
            in2 => \_gnd_net_\,
            in3 => \N__21828\,
            lcout => n317,
            ltout => OPEN,
            carryin => \c0.tx.n4767\,
            carryout => \c0.tx.n4768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23997\,
            in1 => \N__23781\,
            in2 => \_gnd_net_\,
            in3 => \N__21825\,
            lcout => \c0.tx.n5821\,
            ltout => OPEN,
            carryin => \c0.tx.n4768\,
            carryout => \c0.tx.n4769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \_gnd_net_\,
            in3 => \N__21822\,
            lcout => n315,
            ltout => OPEN,
            carryin => \c0.tx.n4769\,
            carryout => \c0.tx.n4770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22133\,
            in1 => \N__24037\,
            in2 => \_gnd_net_\,
            in3 => \N__21819\,
            lcout => \c0.tx.n5884\,
            ltout => OPEN,
            carryin => \c0.tx.n4770\,
            carryout => \c0.tx.n4771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23930\,
            in2 => \_gnd_net_\,
            in3 => \N__21816\,
            lcout => n313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23979\,
            in1 => \N__29010\,
            in2 => \_gnd_net_\,
            in3 => \N__22140\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i33_3_lut_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__29009\,
            in1 => \N__23978\,
            in2 => \_gnd_net_\,
            in3 => \N__23996\,
            lcout => \c0.tx.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24038\,
            in1 => \N__29011\,
            in2 => \_gnd_net_\,
            in3 => \N__22122\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35630\,
            in1 => \N__22115\,
            in2 => \_gnd_net_\,
            in3 => \N__22077\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35978\,
            in1 => \N__22006\,
            in2 => \_gnd_net_\,
            in3 => \N__22056\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_977_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26890\,
            in1 => \N__29503\,
            in2 => \N__23157\,
            in3 => \N__21983\,
            lcout => OPEN,
            ltout => \c0.n42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24555\,
            in1 => \N__25835\,
            in2 => \N__21936\,
            in3 => \N__22589\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i145_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35688\,
            in1 => \N__24168\,
            in2 => \_gnd_net_\,
            in3 => \N__21914\,
            lcout => data_in_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i128_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__35689\,
            in2 => \_gnd_net_\,
            in3 => \N__21853\,
            lcout => data_in_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i136_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35687\,
            in1 => \N__22414\,
            in2 => \_gnd_net_\,
            in3 => \N__23102\,
            lcout => data_in_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_826_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101001"
        )
    port map (
            in0 => \N__22401\,
            in1 => \N__24390\,
            in2 => \N__22395\,
            in3 => \N__24246\,
            lcout => \c0.n22_adj_1890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_855_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24528\,
            in2 => \_gnd_net_\,
            in3 => \N__22365\,
            lcout => \c0.n5384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23180\,
            in1 => \_gnd_net_\,
            in2 => \N__35876\,
            in3 => \N__22300\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__22274\,
            in1 => \N__31997\,
            in2 => \N__33228\,
            in3 => \N__22228\,
            lcout => \c0.data_in_field_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i78_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31996\,
            in1 => \N__33098\,
            in2 => \N__28824\,
            in3 => \N__25983\,
            lcout => \c0.data_in_field_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22188\,
            in1 => \N__23654\,
            in2 => \_gnd_net_\,
            in3 => \N__22166\,
            lcout => OPEN,
            ltout => \c0.n12_adj_1898_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_830_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22604\,
            in1 => \N__22155\,
            in2 => \N__22143\,
            in3 => \N__24135\,
            lcout => OPEN,
            ltout => \c0.n5567_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_834_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111101101111"
        )
    port map (
            in0 => \N__22872\,
            in1 => \N__22860\,
            in2 => \N__22848\,
            in3 => \N__22845\,
            lcout => \c0.n17_adj_1902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6219_bdd_4_lut_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__30200\,
            in1 => \N__25025\,
            in2 => \N__22839\,
            in3 => \N__22824\,
            lcout => \c0.n5707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_948_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22794\,
            in1 => \N__22770\,
            in2 => \N__24999\,
            in3 => \N__22749\,
            lcout => \c0.n5506\,
            ltout => \c0.n5506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_831_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24477\,
            in1 => \N__22719\,
            in2 => \N__22698\,
            in3 => \N__22695\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1010_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22673\,
            in1 => \N__28338\,
            in2 => \N__26859\,
            in3 => \N__22638\,
            lcout => \c0.n5500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_890_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25982\,
            in1 => \N__22575\,
            in2 => \_gnd_net_\,
            in3 => \N__22531\,
            lcout => \c0.n5372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i38_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35981\,
            in1 => \N__25583\,
            in2 => \_gnd_net_\,
            in3 => \N__22502\,
            lcout => data_in_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i42_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22438\,
            in1 => \N__35983\,
            in2 => \_gnd_net_\,
            in3 => \N__22485\,
            lcout => data_in_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i34_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22439\,
            in1 => \N__35982\,
            in2 => \_gnd_net_\,
            in3 => \N__23173\,
            lcout => data_in_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i144_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36052\,
            in1 => \N__23095\,
            in2 => \_gnd_net_\,
            in3 => \N__23149\,
            lcout => data_in_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_964_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23675\,
            in1 => \N__25934\,
            in2 => \N__25454\,
            in3 => \N__25017\,
            lcout => \c0.n6_adj_1918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__31103\,
            in1 => \_gnd_net_\,
            in2 => \N__36073\,
            in3 => \N__23047\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_891_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23676\,
            in1 => \N__25935\,
            in2 => \_gnd_net_\,
            in3 => \N__25018\,
            lcout => OPEN,
            ltout => \c0.n2043_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_992_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23021\,
            in1 => \N__22977\,
            in2 => \N__22971\,
            in3 => \N__22967\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i70_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__26580\,
            in1 => \N__33108\,
            in2 => \N__32171\,
            in3 => \N__25936\,
            lcout => \c0.data_in_field_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i111_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__31994\,
            in1 => \N__23677\,
            in2 => \N__33229\,
            in3 => \N__22923\,
            lcout => \c0.data_in_field_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i102_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__25441\,
            in1 => \N__33107\,
            in2 => \N__34461\,
            in3 => \N__31995\,
            lcout => \c0.data_in_field_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_973_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23298\,
            in1 => \N__26877\,
            in2 => \N__24521\,
            in3 => \N__26951\,
            lcout => \c0.n5443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i49_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__26878\,
            in1 => \N__28800\,
            in2 => \N__32170\,
            in3 => \N__33241\,
            lcout => \c0.data_in_field_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i91_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__23299\,
            in1 => \N__33005\,
            in2 => \N__31260\,
            in3 => \N__32004\,
            lcout => \c0.data_in_field_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_951_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23331\,
            in2 => \_gnd_net_\,
            in3 => \N__23297\,
            lcout => \c0.n1866\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i64_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33238\,
            in1 => \N__32000\,
            in2 => \N__23277\,
            in3 => \N__26952\,
            lcout => \c0.data_in_field_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i63_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31999\,
            in1 => \N__33240\,
            in2 => \N__24529\,
            in3 => \N__24240\,
            lcout => \c0.data_in_field_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i85_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36048\,
            in1 => \N__24959\,
            in2 => \_gnd_net_\,
            in3 => \N__30406\,
            lcout => data_in_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i29_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31998\,
            in1 => \N__33239\,
            in2 => \N__31137\,
            in3 => \N__28224\,
            lcout => \c0.data_in_field_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i38_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33125\,
            in1 => \N__32244\,
            in2 => \N__25599\,
            in3 => \N__23227\,
            lcout => \c0.data_in_field_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i145_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__24176\,
            in2 => \N__33232\,
            in3 => \N__32245\,
            lcout => \c0.data_in_frame_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_943_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27986\,
            in2 => \_gnd_net_\,
            in3 => \N__24781\,
            lcout => \c0.n2077\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6195_bdd_4_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__23610\,
            in1 => \N__23598\,
            in2 => \N__25413\,
            in3 => \N__25158\,
            lcout => \c0.n6198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_852_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23573\,
            in1 => \N__23561\,
            in2 => \N__23550\,
            in3 => \N__23534\,
            lcout => \c0.n18_adj_1919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i41_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35816\,
            in1 => \N__28799\,
            in2 => \_gnd_net_\,
            in3 => \N__23509\,
            lcout => data_in_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i33_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23510\,
            in1 => \N__35819\,
            in2 => \_gnd_net_\,
            in3 => \N__23473\,
            lcout => data_in_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i61_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35818\,
            in1 => \N__23413\,
            in2 => \_gnd_net_\,
            in3 => \N__23456\,
            lcout => data_in_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i51_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33231\,
            in1 => \N__32243\,
            in2 => \N__25662\,
            in3 => \N__24792\,
            lcout => \c0.data_in_field_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i53_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35817\,
            in1 => \N__23414\,
            in2 => \_gnd_net_\,
            in3 => \N__23383\,
            lcout => data_in_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i47_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33230\,
            in1 => \N__32242\,
            in2 => \N__23367\,
            in3 => \N__27994\,
            lcout => \c0.data_in_field_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5299_4_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100000"
        )
    port map (
            in0 => \N__34808\,
            in1 => \N__36230\,
            in2 => \N__36261\,
            in3 => \N__34835\,
            lcout => n5645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5300_4_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011101100"
        )
    port map (
            in0 => \N__34836\,
            in1 => \N__36260\,
            in2 => \N__36234\,
            in3 => \N__34809\,
            lcout => OPEN,
            ltout => \n5646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5301_3_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__36204\,
            in1 => \_gnd_net_\,
            in2 => \N__23721\,
            in3 => \N__23718\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i32_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101101000001"
        )
    port map (
            in0 => \N__37717\,
            in1 => \N__28560\,
            in2 => \N__28713\,
            in3 => \N__26247\,
            lcout => data_out_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i23_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__33669\,
            in1 => \N__34602\,
            in2 => \N__23637\,
            in3 => \N__37715\,
            lcout => data_out_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i25_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__37716\,
            in1 => \N__23831\,
            in2 => \N__33504\,
            in3 => \N__28758\,
            lcout => data_out_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_906_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27987\,
            in1 => \N__24782\,
            in2 => \_gnd_net_\,
            in3 => \N__23684\,
            lcout => \c0.n5533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_931_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35040\,
            in1 => \N__34970\,
            in2 => \_gnd_net_\,
            in3 => \N__34707\,
            lcout => n4_adj_1975,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i17_3_lut_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34326\,
            in1 => \N__28548\,
            in2 => \_gnd_net_\,
            in3 => \N__23633\,
            lcout => OPEN,
            ltout => \c0.n17_adj_1913_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5575_3_lut_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__33781\,
            in1 => \_gnd_net_\,
            in2 => \N__23751\,
            in3 => \N__34072\,
            lcout => \c0.n5830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_894_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33665\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35038\,
            lcout => n4_adj_1982,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i957_4_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000111000100"
        )
    port map (
            in0 => \N__34211\,
            in1 => \N__34070\,
            in2 => \N__28770\,
            in3 => \N__34325\,
            lcout => \c0.n1198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__29282\,
            in1 => \N__23748\,
            in2 => \N__33612\,
            in3 => \N__23808\,
            lcout => \c0.tx.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_904_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34971\,
            lcout => n1991,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5563_3_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__34071\,
            in1 => \N__33780\,
            in2 => \_gnd_net_\,
            in3 => \N__26235\,
            lcout => \c0.n5827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i746_2_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34132\,
            in2 => \_gnd_net_\,
            in3 => \N__34079\,
            lcout => \c0.n1253\,
            ltout => \c0.n1253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__33633\,
            in1 => \N__26169\,
            in2 => \N__23742\,
            in3 => \N__33738\,
            lcout => \tx_data_2_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_841_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100100010"
        )
    port map (
            in0 => \N__34328\,
            in1 => \N__34212\,
            in2 => \N__33396\,
            in3 => \N__34080\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001101"
        )
    port map (
            in0 => \N__33739\,
            in1 => \N__23739\,
            in2 => \N__23730\,
            in3 => \N__34134\,
            lcout => \tx_data_6_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__26295\,
            in1 => \N__23877\,
            in2 => \N__23871\,
            in3 => \N__33740\,
            lcout => \tx_data_7_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5588_4_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__23846\,
            in1 => \N__26200\,
            in2 => \N__23835\,
            in3 => \N__34327\,
            lcout => OPEN,
            ltout => \c0.n5810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__34133\,
            in1 => \N__23817\,
            in2 => \N__23811\,
            in3 => \N__33737\,
            lcout => \c0.tx_data_0_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5281_4_lut_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24096\,
            in1 => \N__23929\,
            in2 => \N__24069\,
            in3 => \N__23778\,
            lcout => \c0.tx.n5627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i6_4_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24066\,
            in1 => \N__24097\,
            in2 => \N__23984\,
            in3 => \N__24033\,
            lcout => OPEN,
            ltout => \c0.tx.n14_adj_1869_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7_4_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24045\,
            in1 => \N__26280\,
            in2 => \N__23796\,
            in3 => \N__23779\,
            lcout => \c0.tx.r_SM_Main_2_N_1767_1\,
            ltout => \c0.tx.r_SM_Main_2_N_1767_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__28976\,
            in1 => \N__29174\,
            in2 => \N__23793\,
            in3 => \N__29090\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__23790\,
            in1 => \N__23780\,
            in2 => \N__23985\,
            in3 => \N__28978\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__26458\,
            in2 => \N__23763\,
            in3 => \N__24098\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__28977\,
            in2 => \N__24081\,
            in3 => \N__24067\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26533\,
            lcout => \c0.tx.n10_adj_1868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5283_3_lut_4_lut_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__26532\,
            in1 => \N__26493\,
            in2 => \N__24039\,
            in3 => \N__26412\,
            lcout => \c0.tx.n5629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29198\,
            in2 => \_gnd_net_\,
            in3 => \N__29070\,
            lcout => n11_adj_1979,
            ltout => \n11_adj_1979_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_adj_805_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28956\,
            in1 => \N__24012\,
            in2 => \N__24006\,
            in3 => \N__24003\,
            lcout => \c0.tx.n3120\,
            ltout => \c0.tx.n3120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__23980\,
            in1 => \_gnd_net_\,
            in2 => \N__23946\,
            in3 => \N__28957\,
            lcout => n782,
            ltout => \n782_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__28958\,
            in1 => \N__23943\,
            in2 => \N__23934\,
            in3 => \N__23931\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i75_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35631\,
            in1 => \N__23890\,
            in2 => \_gnd_net_\,
            in3 => \N__30671\,
            lcout => data_in_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_819_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24453\,
            in1 => \N__24447\,
            in2 => \N__24426\,
            in3 => \N__24411\,
            lcout => \c0.n24_adj_1885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25555\,
            in1 => \N__26739\,
            in2 => \N__25901\,
            in3 => \N__24384\,
            lcout => OPEN,
            ltout => \c0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_822_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24366\,
            in1 => \N__24324\,
            in2 => \N__24273\,
            in3 => \N__24270\,
            lcout => \c0.n5519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28419\,
            in1 => \N__35685\,
            in2 => \_gnd_net_\,
            in3 => \N__27861\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i55_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24202\,
            in1 => \N__35686\,
            in2 => \_gnd_net_\,
            in3 => \N__24239\,
            lcout => data_in_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i45_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__32128\,
            in1 => \N__24890\,
            in2 => \N__27363\,
            in3 => \N__33103\,
            lcout => \c0.data_in_field_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i137_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30694\,
            in1 => \_gnd_net_\,
            in2 => \N__36063\,
            in3 => \N__24169\,
            lcout => data_in_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i101_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__24845\,
            in1 => \N__33102\,
            in2 => \N__24990\,
            in3 => \N__32129\,
            lcout => \c0.data_in_field_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_998_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24144\,
            in1 => \N__24134\,
            in2 => \N__24120\,
            in3 => \N__24914\,
            lcout => \c0.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_856_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24886\,
            in2 => \_gnd_net_\,
            in3 => \N__24832\,
            lcout => \c0.n4_adj_1920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_996_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24802\,
            in1 => \N__24750\,
            in2 => \N__24732\,
            in3 => \N__24714\,
            lcout => OPEN,
            ltout => \c0.n31_adj_1900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_833_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26586\,
            in1 => \N__25068\,
            in2 => \N__24693\,
            in3 => \N__24690\,
            lcout => \c0.n5582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i3_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__33104\,
            in1 => \N__27241\,
            in2 => \N__24684\,
            in3 => \N__32131\,
            lcout => \c0.data_in_field_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37542\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_838_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101101"
        )
    port map (
            in0 => \N__24651\,
            in1 => \N__24645\,
            in2 => \N__24639\,
            in3 => \N__24627\,
            lcout => \c0.n25_adj_1907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_858_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30243\,
            in1 => \N__24612\,
            in2 => \N__27242\,
            in3 => \N__24604\,
            lcout => \c0.n5593\,
            ltout => \c0.n5593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_974_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24527\,
            in1 => \N__26897\,
            in2 => \N__24480\,
            in3 => \N__26960\,
            lcout => \c0.n5430\,
            ltout => \c0.n5430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_999_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27032\,
            in1 => \N__24471\,
            in2 => \N__24465\,
            in3 => \N__24462\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i14_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__33106\,
            in1 => \N__25062\,
            in2 => \N__25026\,
            in3 => \N__32127\,
            lcout => \c0.data_in_field_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25789\,
            in1 => \N__30569\,
            in2 => \N__30935\,
            in3 => \N__30534\,
            lcout => \c0.n6_adj_1939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i101_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24982\,
            in1 => \_gnd_net_\,
            in2 => \N__30291\,
            in3 => \N__35906\,
            lcout => data_in_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i89_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__28339\,
            in1 => \N__32130\,
            in2 => \N__30483\,
            in3 => \N__33105\,
            lcout => \c0.data_in_field_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i65_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25869\,
            in1 => \N__35907\,
            in2 => \_gnd_net_\,
            in3 => \N__31045\,
            lcout => data_in_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i93_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35905\,
            in1 => \N__24958\,
            in2 => \_gnd_net_\,
            in3 => \N__24983\,
            lcout => data_in_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_942_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30926\,
            in2 => \_gnd_net_\,
            in3 => \N__25788\,
            lcout => \c0.n2089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_868_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27443\,
            in2 => \_gnd_net_\,
            in3 => \N__24927\,
            lcout => \c0.n5581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i88_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32992\,
            in1 => \N__32164\,
            in2 => \N__28121\,
            in3 => \N__31367\,
            lcout => \c0.data_in_field_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i73_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32161\,
            in1 => \N__32994\,
            in2 => \N__25868\,
            in3 => \N__25793\,
            lcout => \c0.data_in_field_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i129_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32991\,
            in1 => \N__32163\,
            in2 => \N__35103\,
            in3 => \N__28045\,
            lcout => \c0.data_in_field_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i121_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32990\,
            in1 => \N__32162\,
            in2 => \N__35073\,
            in3 => \N__25543\,
            lcout => \c0.data_in_field_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i43_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32160\,
            in1 => \N__32993\,
            in2 => \N__25629\,
            in3 => \N__25828\,
            lcout => \c0.data_in_field_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_969_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28277\,
            in1 => \N__25542\,
            in2 => \_gnd_net_\,
            in3 => \N__28044\,
            lcout => \c0.n2107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i155_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25894\,
            in1 => \N__25500\,
            in2 => \_gnd_net_\,
            in3 => \N__35918\,
            lcout => data_in_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6201_bdd_4_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__25479\,
            in1 => \N__26646\,
            in2 => \N__30206\,
            in3 => \N__25462\,
            lcout => OPEN,
            ltout => \c0.n5716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_5844_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__25409\,
            in1 => \N__25259\,
            in2 => \N__25161\,
            in3 => \N__25914\,
            lcout => \c0.n6195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5829_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__27743\,
            in1 => \N__25152\,
            in2 => \N__30205\,
            in3 => \N__25113\,
            lcout => OPEN,
            ltout => \c0.n6207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6207_bdd_4_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__25994\,
            in1 => \N__30180\,
            in2 => \N__25950\,
            in3 => \N__25946\,
            lcout => \c0.n5713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i147_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25893\,
            in2 => \N__36022\,
            in3 => \N__25714\,
            lcout => data_in_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i73_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30453\,
            in1 => \N__25861\,
            in2 => \_gnd_net_\,
            in3 => \N__35919\,
            lcout => data_in_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_875_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25821\,
            in2 => \_gnd_net_\,
            in3 => \N__25787\,
            lcout => \c0.n2068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i89_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35821\,
            in1 => \N__25764\,
            in2 => \_gnd_net_\,
            in3 => \N__30469\,
            lcout => data_in_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i139_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25715\,
            in1 => \N__25673\,
            in2 => \_gnd_net_\,
            in3 => \N__35822\,
            lcout => data_in_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i43_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__35823\,
            in2 => \_gnd_net_\,
            in3 => \N__25615\,
            lcout => data_in_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35820\,
            in1 => \N__25595\,
            in2 => \_gnd_net_\,
            in3 => \N__27889\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i88_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35824\,
            in1 => \N__26162\,
            in2 => \_gnd_net_\,
            in3 => \N__31357\,
            lcout => data_in_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33457\,
            in2 => \_gnd_net_\,
            in3 => \N__33336\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26123\,
            in1 => \N__26111\,
            in2 => \_gnd_net_\,
            in3 => \N__34332\,
            lcout => \c0.n17_adj_1908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_968_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36518\,
            in1 => \N__34657\,
            in2 => \_gnd_net_\,
            in3 => \N__35013\,
            lcout => OPEN,
            ltout => \n5448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i29_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__37708\,
            in1 => \N__26124\,
            in2 => \N__26136\,
            in3 => \N__26133\,
            lcout => data_out_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i21_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010001011"
        )
    port map (
            in0 => \N__26112\,
            in1 => \N__37707\,
            in2 => \N__33516\,
            in3 => \N__28692\,
            lcout => data_out_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_859_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26103\,
            in1 => \N__26085\,
            in2 => \N__26067\,
            in3 => \N__26049\,
            lcout => OPEN,
            ltout => \c0.n20_adj_1922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_862_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26043\,
            in1 => \N__26025\,
            in2 => \N__26007\,
            in3 => \N__26004\,
            lcout => n21_adj_1977,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5571_4_lut_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__34324\,
            in1 => \N__26475\,
            in2 => \N__28533\,
            in3 => \N__26201\,
            lcout => \c0.n5833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_865_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36731\,
            in2 => \_gnd_net_\,
            in3 => \N__36825\,
            lcout => n4334,
            ltout => \n4334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i28_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000101"
        )
    port map (
            in0 => \N__28517\,
            in1 => \N__33926\,
            in2 => \N__26256\,
            in3 => \N__26253\,
            lcout => data_out_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26246\,
            in1 => \N__26213\,
            in2 => \_gnd_net_\,
            in3 => \N__34323\,
            lcout => \c0.n17_adj_1950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i27_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__26186\,
            in1 => \N__26229\,
            in2 => \N__28518\,
            in3 => \N__37702\,
            lcout => data_out_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__26202\,
            in1 => \N__33678\,
            in2 => \N__26223\,
            in3 => \N__33722\,
            lcout => \tx_data_4_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i24_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__26214\,
            in1 => \N__36732\,
            in2 => \N__28674\,
            in3 => \N__36826\,
            lcout => data_out_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_997_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__34204\,
            in1 => \N__34130\,
            in2 => \_gnd_net_\,
            in3 => \N__34067\,
            lcout => \c0.n1508\,
            ltout => \c0.n1508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5587_4_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__26187\,
            in1 => \N__26303\,
            in2 => \N__26172\,
            in3 => \N__34331\,
            lcout => \c0.n5840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010011101100"
        )
    port map (
            in0 => \N__34206\,
            in1 => \N__34131\,
            in2 => \N__28650\,
            in3 => \N__34068\,
            lcout => OPEN,
            ltout => \c0.n6309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6309_bdd_4_lut_4_lut_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000111100011"
        )
    port map (
            in0 => \N__34069\,
            in1 => \N__34207\,
            in2 => \N__26307\,
            in3 => \N__34330\,
            lcout => \c0.n6312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i19_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__26304\,
            in1 => \N__37706\,
            in2 => \N__36591\,
            in3 => \N__36440\,
            lcout => data_out_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1006_4_lut_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__34531\,
            in1 => \N__34205\,
            in2 => \N__36519\,
            in3 => \N__34329\,
            lcout => \c0.n1249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__28452\,
            in1 => \N__29091\,
            in2 => \_gnd_net_\,
            in3 => \N__29321\,
            lcout => \c0.tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_857_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34658\,
            lcout => n1768,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33598\,
            in1 => \N__33833\,
            in2 => \_gnd_net_\,
            in3 => \N__26289\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i3401_2_lut_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26494\,
            in2 => \_gnd_net_\,
            in3 => \N__26413\,
            lcout => \c0.tx.n3644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5566_2_lut_3_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29204\,
            in1 => \N__29087\,
            in2 => \_gnd_net_\,
            in3 => \N__28485\,
            lcout => OPEN,
            ltout => \n5818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Done_44_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111000"
        )
    port map (
            in0 => \N__26265\,
            in1 => \N__26274\,
            in2 => \N__26268\,
            in3 => \N__28973\,
            lcout => n4155,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__28968\,
            in1 => \N__26460\,
            in2 => \N__26550\,
            in3 => \N__26537\,
            lcout => \r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__26459\,
            in1 => \N__28969\,
            in2 => \N__26511\,
            in3 => \N__26495\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29205\,
            in1 => \N__29088\,
            in2 => \N__29004\,
            in3 => \N__28486\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i22_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__33624\,
            in1 => \N__26474\,
            in2 => \N__37757\,
            in3 => \N__37726\,
            lcout => data_out_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__26456\,
            in2 => \N__26436\,
            in3 => \N__26417\,
            lcout => \r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i154_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35760\,
            in1 => \N__26391\,
            in2 => \_gnd_net_\,
            in3 => \N__26700\,
            lcout => data_in_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i108_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35693\,
            in1 => \N__26366\,
            in2 => \_gnd_net_\,
            in3 => \N__26321\,
            lcout => data_in_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i129_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__30695\,
            in2 => \_gnd_net_\,
            in3 => \N__35086\,
            lcout => data_in_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i86_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36020\,
            in1 => \N__27014\,
            in2 => \_gnd_net_\,
            in3 => \N__28840\,
            lcout => data_in_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i109_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26918\,
            in1 => \N__36021\,
            in2 => \_gnd_net_\,
            in3 => \N__30280\,
            lcout => data_in_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5661_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__26991\,
            in1 => \N__27754\,
            in2 => \N__30209\,
            in3 => \N__26964\,
            lcout => \c0.n5997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i117_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36019\,
            in1 => \N__26917\,
            in2 => \_gnd_net_\,
            in3 => \N__30308\,
            lcout => data_in_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5685_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__30198\,
            in1 => \N__27755\,
            in2 => \N__26904\,
            in3 => \N__29460\,
            lcout => OPEN,
            ltout => \c0.n6033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n6033_bdd_4_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__26858\,
            in1 => \N__26805\,
            in2 => \N__26754\,
            in3 => \N__30199\,
            lcout => \c0.n5791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_889_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27909\,
            in1 => \N__29361\,
            in2 => \N__28143\,
            in3 => \N__30903\,
            lcout => \c0.n1814\,
            ltout => \c0.n1814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_993_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26710\,
            in1 => \N__26676\,
            in2 => \N__26649\,
            in3 => \N__26644\,
            lcout => \c0.n32_adj_1901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i85_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33070\,
            in1 => \N__32230\,
            in2 => \N__30423\,
            in3 => \N__29542\,
            lcout => \c0.data_in_field_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i70_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35878\,
            in1 => \N__28817\,
            in2 => \_gnd_net_\,
            in3 => \N__26579\,
            lcout => data_in_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i133_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35499\,
            in1 => \N__27399\,
            in2 => \_gnd_net_\,
            in3 => \N__30340\,
            lcout => data_in_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i37_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35877\,
            in1 => \N__31210\,
            in2 => \_gnd_net_\,
            in3 => \N__27356\,
            lcout => data_in_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i25_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__27856\,
            in1 => \N__32229\,
            in2 => \N__33218\,
            in3 => \N__27442\,
            lcout => \c0.data_in_field_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_913_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27435\,
            in1 => \N__30593\,
            in2 => \N__31407\,
            in3 => \N__30561\,
            lcout => \c0.n5560\,
            ltout => \c0.n5560_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27300\,
            in1 => \N__27234\,
            in2 => \N__27213\,
            in3 => \N__30230\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i40_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35923\,
            in1 => \N__31432\,
            in2 => \_gnd_net_\,
            in3 => \N__27188\,
            lcout => data_in_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_947_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27164\,
            in1 => \N__27138\,
            in2 => \N__30606\,
            in3 => \N__27099\,
            lcout => \c0.n5378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i94_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35925\,
            in1 => \N__27007\,
            in2 => \_gnd_net_\,
            in3 => \N__34457\,
            lcout => data_in_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i99_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__33234\,
            in1 => \N__28281\,
            in2 => \N__32241\,
            in3 => \N__31277\,
            lcout => \c0.data_in_field_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i17_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32165\,
            in1 => \N__28433\,
            in2 => \N__33272\,
            in3 => \N__30934\,
            lcout => \c0.data_in_field_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i99_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__35924\,
            in1 => \N__28391\,
            in2 => \N__31281\,
            in3 => \_gnd_net_\,
            lcout => data_in_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_4_lut_adj_1001_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28332\,
            in1 => \N__28270\,
            in2 => \N__28234\,
            in3 => \N__28197\,
            lcout => \c0.n23_adj_1935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_878_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28096\,
            in2 => \_gnd_net_\,
            in3 => \N__28043\,
            lcout => OPEN,
            ltout => \c0.n1965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_887_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28016\,
            in1 => \N__28001\,
            in2 => \N__27960\,
            in3 => \N__27953\,
            lcout => \c0.n24_adj_1930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_876_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27882\,
            in1 => \N__27857\,
            in2 => \N__31130\,
            in3 => \N__27814\,
            lcout => \c0.n28_adj_1925\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_5704_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__27744\,
            in1 => \N__27444\,
            in2 => \N__30194\,
            in3 => \N__30933\,
            lcout => \c0.n6039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i16_3_lut_4_lut_4_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__29202\,
            in1 => \N__29113\,
            in2 => \N__28608\,
            in3 => \N__28497\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010111010"
        )
    port map (
            in0 => \N__28637\,
            in1 => \N__29015\,
            in2 => \N__28506\,
            in3 => \N__29114\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_809_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28503\,
            in2 => \_gnd_net_\,
            in3 => \N__28636\,
            lcout => \c0.n50_adj_1875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_1793_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_adj_804_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__29201\,
            in1 => \N__29112\,
            in2 => \N__29021\,
            in3 => \N__28496\,
            lcout => \c0.tx.n2177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33356\,
            in1 => \N__33332\,
            in2 => \_gnd_net_\,
            in3 => \N__33302\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33456\,
            in2 => \_gnd_net_\,
            in3 => \N__33357\,
            lcout => \c0.byte_transmit_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5640_3_lut_4_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__33488\,
            in1 => \N__28639\,
            in2 => \N__28597\,
            in3 => \N__33524\,
            lcout => n4333,
            ltout => \n4333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i10_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__36828\,
            in1 => \N__36303\,
            in2 => \N__28443\,
            in3 => \N__35008\,
            lcout => data_out_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__28583\,
            in1 => \N__28640\,
            in2 => \_gnd_net_\,
            in3 => \N__36827\,
            lcout => \c0.n81_adj_1872\,
            ltout => \c0.n81_adj_1872_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__33282\,
            in1 => \N__33437\,
            in2 => \N__28440\,
            in3 => \N__33489\,
            lcout => \c0.byte_transmit_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_1794_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33490\,
            in1 => \N__28641\,
            in2 => \N__28598\,
            in3 => \N__33525\,
            lcout => \c0.tx_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_975_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36954\,
            in1 => \N__33972\,
            in2 => \_gnd_net_\,
            in3 => \N__36408\,
            lcout => n135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_873_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36681\,
            lcout => n5482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_994_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34431\,
            in1 => \N__36683\,
            in2 => \_gnd_net_\,
            in3 => \N__36635\,
            lcout => n5433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_813_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__36554\,
            in1 => \_gnd_net_\,
            in2 => \N__35018\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n4_adj_1986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i31_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__37705\,
            in1 => \N__28746\,
            in2 => \N__28551\,
            in3 => \N__28547\,
            lcout => data_out_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i30_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__34917\,
            in1 => \N__37704\,
            in2 => \N__33798\,
            in3 => \N__28532\,
            lcout => data_out_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i18_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__33950\,
            in1 => \N__37703\,
            in2 => \N__34905\,
            in3 => \N__33971\,
            lcout => data_out_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_930_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34659\,
            in1 => \N__34430\,
            in2 => \N__36508\,
            in3 => \N__35012\,
            lcout => n5440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34279\,
            in1 => \_gnd_net_\,
            in2 => \N__36564\,
            in3 => \N__34380\,
            lcout => \c0.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36495\,
            in1 => \N__28745\,
            in2 => \_gnd_net_\,
            in3 => \N__36687\,
            lcout => n8_adj_1987,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_963_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33967\,
            in1 => \N__36413\,
            in2 => \N__36965\,
            in3 => \N__34381\,
            lcout => n5400,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33611\,
            in1 => \N__28734\,
            in2 => \_gnd_net_\,
            in3 => \N__29346\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_987_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36430\,
            in1 => \N__36412\,
            in2 => \N__36966\,
            in3 => \N__34382\,
            lcout => n5364,
            ltout => \n5364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5552_4_lut_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28709\,
            in1 => \N__28688\,
            in2 => \N__28677\,
            in3 => \N__34429\,
            lcout => n5871,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__28665\,
            in1 => \N__33912\,
            in2 => \N__33782\,
            in3 => \N__33736\,
            lcout => \tx_data_3_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__29355\,
            in1 => \_gnd_net_\,
            in2 => \N__28659\,
            in3 => \N__33610\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5572_4_lut_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__36614\,
            in1 => \N__34066\,
            in2 => \N__36414\,
            in3 => \N__34319\,
            lcout => \c0.n5853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0__bdd_4_lut_5889_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__29354\,
            in1 => \N__29345\,
            in2 => \N__33894\,
            in3 => \N__29317\,
            lcout => OPEN,
            ltout => \c0.tx.n6051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n6051_bdd_4_lut_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__29264\,
            in1 => \N__29286\,
            in2 => \N__29268\,
            in3 => \N__33892\,
            lcout => \c0.tx.n6054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33571\,
            in1 => \N__29265\,
            in2 => \_gnd_net_\,
            in3 => \N__33687\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i367827_i1_3_lut_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29252\,
            in1 => \N__29211\,
            in2 => \_gnd_net_\,
            in3 => \N__33804\,
            lcout => OPEN,
            ltout => \c0.tx.o_Tx_Serial_N_1798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i26_3_lut_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29199\,
            in2 => \N__29124\,
            in3 => \N__29117\,
            lcout => OPEN,
            ltout => \c0.tx.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28868\,
            in2 => \N__29025\,
            in3 => \N__28979\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i78_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35880\,
            in1 => \N__28841\,
            in2 => \_gnd_net_\,
            in3 => \N__28816\,
            lcout => data_in_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i49_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35879\,
            in1 => \N__31031\,
            in2 => \_gnd_net_\,
            in3 => \N__28781\,
            lcout => data_in_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i77_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35899\,
            in1 => \N__30367\,
            in2 => \_gnd_net_\,
            in3 => \N__30419\,
            lcout => data_in_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i125_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30307\,
            in1 => \N__35980\,
            in2 => \_gnd_net_\,
            in3 => \N__30341\,
            lcout => data_in_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i109_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33074\,
            in1 => \N__32133\,
            in2 => \N__30290\,
            in3 => \N__30250\,
            lcout => \c0.data_in_field_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i71_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__29484\,
            in1 => \N__33076\,
            in2 => \N__31169\,
            in3 => \N__32232\,
            lcout => \c0.data_in_field_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5997_bdd_4_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__30210\,
            in1 => \N__31411\,
            in2 => \N__29625\,
            in3 => \N__29586\,
            lcout => \c0.n6000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i57_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__29459\,
            in1 => \N__33075\,
            in2 => \N__31032\,
            in3 => \N__32231\,
            lcout => \c0.data_in_field_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_880_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29535\,
            in1 => \N__29483\,
            in2 => \_gnd_net_\,
            in3 => \N__29458\,
            lcout => \c0.n5494\,
            ltout => \c0.n5494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_884_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29429\,
            in1 => \N__29412\,
            in2 => \N__29385\,
            in3 => \N__29378\,
            lcout => \c0.n26_adj_1927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i57_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35979\,
            in1 => \N__31027\,
            in2 => \_gnd_net_\,
            in3 => \N__31058\,
            lcout => data_in_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_888_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31013\,
            in1 => \N__30974\,
            in2 => \N__30936\,
            in3 => \N__30489\,
            lcout => \c0.n25_adj_1931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_965_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31400\,
            in1 => \N__30897\,
            in2 => \N__30846\,
            in3 => \N__30780\,
            lcout => \c0.n5542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i137_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33153\,
            in1 => \N__32134\,
            in2 => \N__30705\,
            in3 => \N__30568\,
            lcout => \c0.data_in_field_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i83_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36074\,
            in1 => \N__31253\,
            in2 => \_gnd_net_\,
            in3 => \N__30658\,
            lcout => data_in_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i39_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__33154\,
            in1 => \N__32135\,
            in2 => \N__30642\,
            in3 => \N__30605\,
            lcout => \c0.data_in_field_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33466\,
            in2 => \_gnd_net_\,
            in3 => \N__33306\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_941_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30560\,
            in2 => \_gnd_net_\,
            in3 => \N__30530\,
            lcout => \c0.n2113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i81_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36015\,
            in1 => \N__30482\,
            in2 => \_gnd_net_\,
            in3 => \N__30439\,
            lcout => data_in_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i40_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__32989\,
            in1 => \N__32169\,
            in2 => \N__31412\,
            in3 => \N__31436\,
            lcout => \c0.data_in_field_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i80_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36014\,
            in1 => \N__31322\,
            in2 => \_gnd_net_\,
            in3 => \N__31368\,
            lcout => data_in_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i110_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35900\,
            in1 => \N__31310\,
            in2 => \_gnd_net_\,
            in3 => \N__34477\,
            lcout => data_in_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i91_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36058\,
            in1 => \N__31246\,
            in2 => \_gnd_net_\,
            in3 => \N__31276\,
            lcout => data_in_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36057\,
            in1 => \N__31223\,
            in2 => \_gnd_net_\,
            in3 => \N__31125\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i71_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36062\,
            in1 => \N__31197\,
            in2 => \_gnd_net_\,
            in3 => \N__31153\,
            lcout => data_in_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36056\,
            in1 => \N__31089\,
            in2 => \_gnd_net_\,
            in3 => \N__31126\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31068\,
            in2 => \N__34278\,
            in3 => \N__37734\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \c0.n4703\,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__37735\,
            in1 => \N__34017\,
            in2 => \_gnd_net_\,
            in3 => \N__33375\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n4703\,
            carryout => \c0.n4704\,
            clk => \N__37595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_4_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34108\,
            in2 => \_gnd_net_\,
            in3 => \N__33372\,
            lcout => \c0.tx_transmit_N_568_2\,
            ltout => OPEN,
            carryin => \c0.n4704\,
            carryout => \c0.n4705\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_5_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34187\,
            in3 => \N__33369\,
            lcout => \c0.tx_transmit_N_568_3\,
            ltout => OPEN,
            carryin => \c0.n4705\,
            carryout => \c0.n4706\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_6_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33713\,
            in2 => \_gnd_net_\,
            in3 => \N__33366\,
            lcout => \c0.tx_transmit_N_568_4\,
            ltout => OPEN,
            carryin => \c0.n4706\,
            carryout => \c0.n4707\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_7_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33363\,
            in2 => \_gnd_net_\,
            in3 => \N__33348\,
            lcout => \c0.tx_transmit_N_568_5\,
            ltout => OPEN,
            carryin => \c0.n4707\,
            carryout => \c0.n4708\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_8_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33345\,
            in2 => \_gnd_net_\,
            in3 => \N__33321\,
            lcout => \c0.tx_transmit_N_568_6\,
            ltout => OPEN,
            carryin => \c0.n4708\,
            carryout => \c0.n4709\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_1824_9_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__33318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33309\,
            lcout => \c0.tx_transmit_N_568_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33436\,
            in2 => \N__33471\,
            in3 => \N__33492\,
            lcout => \c0.byte_transmit_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_842_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33416\,
            in2 => \_gnd_net_\,
            in3 => \N__33290\,
            lcout => \c0.n95\,
            ltout => \c0.n95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i120_2_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33528\,
            in3 => \N__33432\,
            lcout => \c0.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_995_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34533\,
            in1 => \N__33664\,
            in2 => \N__34383\,
            in3 => \N__36120\,
            lcout => n4_adj_1981,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36175\,
            in1 => \N__36641\,
            in2 => \_gnd_net_\,
            in3 => \N__34650\,
            lcout => n7_adj_1988,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__33467\,
            in2 => \N__33438\,
            in3 => \N__33417\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i13_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34962\,
            in1 => \N__36892\,
            in2 => \N__37110\,
            in3 => \N__36752\,
            lcout => data_out_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__33381\,
            in1 => \N__33723\,
            in2 => \N__33408\,
            in3 => \N__34116\,
            lcout => \tx_data_5_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1000_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33656\,
            in1 => \N__36173\,
            in2 => \_gnd_net_\,
            in3 => \N__34375\,
            lcout => n5424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i35_3_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34649\,
            in1 => \N__36119\,
            in2 => \_gnd_net_\,
            in3 => \N__34302\,
            lcout => \c0.n31_adj_1912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i748_4_lut_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100100010"
        )
    port map (
            in0 => \N__34303\,
            in1 => \N__34173\,
            in2 => \N__34395\,
            in3 => \N__34058\,
            lcout => \c0.n989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34945\,
            in1 => \N__33655\,
            in2 => \_gnd_net_\,
            in3 => \N__34301\,
            lcout => OPEN,
            ltout => \c0.n9_adj_1906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i15_4_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001110111"
        )
    port map (
            in0 => \N__34115\,
            in1 => \N__34172\,
            in2 => \N__33681\,
            in3 => \N__34057\,
            lcout => \c0.n15_adj_1909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i951_2_lut_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34171\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34114\,
            lcout => \c0.n1251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i5_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__33657\,
            in1 => \N__36897\,
            in2 => \N__37866\,
            in3 => \N__36748\,
            lcout => data_out_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2044_4_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__36169\,
            in1 => \N__34197\,
            in2 => \N__36964\,
            in3 => \N__34320\,
            lcout => \c0.n2293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i16_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34521\,
            in1 => \N__36898\,
            in2 => \N__37044\,
            in3 => \N__36783\,
            lcout => data_out_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_933_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34695\,
            in1 => \N__34518\,
            in2 => \N__34969\,
            in3 => \N__36111\,
            lcout => n5479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_844_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36499\,
            lcout => n4_adj_1996,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33609\,
            in1 => \N__33906\,
            in2 => \_gnd_net_\,
            in3 => \N__33534\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1005_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34696\,
            in1 => \N__34519\,
            in2 => \N__34968\,
            in3 => \N__36112\,
            lcout => n5421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i8_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__36785\,
            in1 => \N__37791\,
            in2 => \N__36500\,
            in3 => \N__36894\,
            lcout => data_out_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5595_4_lut_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__33951\,
            in1 => \N__34060\,
            in2 => \N__36348\,
            in3 => \N__34322\,
            lcout => \c0.n5845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i4_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__36784\,
            in1 => \N__36639\,
            in2 => \N__37887\,
            in3 => \N__36893\,
            lcout => data_out_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5582_4_lut_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__37641\,
            in1 => \N__34059\,
            in2 => \N__33936\,
            in3 => \N__34321\,
            lcout => \c0.n5837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.n6285_bdd_4_lut_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__33905\,
            in1 => \N__33883\,
            in2 => \N__33834\,
            in3 => \N__33816\,
            lcout => \c0.tx.n6288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i9_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__36786\,
            in1 => \N__36550\,
            in2 => \N__36327\,
            in3 => \N__36895\,
            lcout => data_out_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_897_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36109\,
            lcout => n5415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__33984\,
            in1 => \N__33783\,
            in2 => \N__33753\,
            in3 => \N__33744\,
            lcout => \tx_data_1_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_937_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34705\,
            in1 => \N__36108\,
            in2 => \_gnd_net_\,
            in3 => \N__34532\,
            lcout => n1579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i102_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35999\,
            in1 => \N__34478\,
            in2 => \_gnd_net_\,
            in3 => \N__34444\,
            lcout => data_in_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i6_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34419\,
            in1 => \N__36900\,
            in2 => \N__37842\,
            in3 => \N__36791\,
            lcout => data_out_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34682\,
            in1 => \N__34411\,
            in2 => \_gnd_net_\,
            in3 => \N__34269\,
            lcout => \c0.n9_adj_1911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i1_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__34379\,
            in1 => \N__37023\,
            in2 => \N__36912\,
            in3 => \N__36769\,
            lcout => data_out_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35014\,
            in1 => \N__36666\,
            in2 => \_gnd_net_\,
            in3 => \N__34270\,
            lcout => OPEN,
            ltout => \c0.n9_adj_1891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010010011001"
        )
    port map (
            in0 => \N__34186\,
            in1 => \N__34117\,
            in2 => \N__34083\,
            in3 => \N__34036\,
            lcout => \c0.n15_adj_1893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i7_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34642\,
            in1 => \N__36902\,
            in2 => \N__37818\,
            in3 => \N__36771\,
            lcout => data_out_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i2_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__36770\,
            in1 => \N__37005\,
            in2 => \N__36911\,
            in3 => \N__36667\,
            lcout => data_out_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i14_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__34694\,
            in1 => \N__36901\,
            in2 => \N__37086\,
            in3 => \N__36768\,
            lcout => data_out_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_959_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36174\,
            in1 => \N__34641\,
            in2 => \_gnd_net_\,
            in3 => \N__36566\,
            lcout => n4_adj_1976,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i0_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34593\,
            in2 => \_gnd_net_\,
            in3 => \N__34587\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => n4710,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i1_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34584\,
            in2 => \_gnd_net_\,
            in3 => \N__34578\,
            lcout => n25,
            ltout => OPEN,
            carryin => n4710,
            carryout => n4711,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i2_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34575\,
            in2 => \_gnd_net_\,
            in3 => \N__34569\,
            lcout => n24,
            ltout => OPEN,
            carryin => n4711,
            carryout => n4712,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i3_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34566\,
            in2 => \_gnd_net_\,
            in3 => \N__34560\,
            lcout => n23,
            ltout => OPEN,
            carryin => n4712,
            carryout => n4713,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i4_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34557\,
            in2 => \_gnd_net_\,
            in3 => \N__34551\,
            lcout => n22,
            ltout => OPEN,
            carryin => n4713,
            carryout => n4714,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i5_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34548\,
            in2 => \_gnd_net_\,
            in3 => \N__34542\,
            lcout => n21,
            ltout => OPEN,
            carryin => n4714,
            carryout => n4715,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i6_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34539\,
            in2 => \_gnd_net_\,
            in3 => \N__34782\,
            lcout => n20,
            ltout => OPEN,
            carryin => n4715,
            carryout => n4716,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i7_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34779\,
            in2 => \_gnd_net_\,
            in3 => \N__34773\,
            lcout => n19,
            ltout => OPEN,
            carryin => n4716,
            carryout => n4717,
            clk => \N__37612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i8_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34770\,
            in2 => \_gnd_net_\,
            in3 => \N__34764\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => n4718,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i9_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34761\,
            in2 => \_gnd_net_\,
            in3 => \N__34755\,
            lcout => n17,
            ltout => OPEN,
            carryin => n4718,
            carryout => n4719,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i10_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34752\,
            in2 => \_gnd_net_\,
            in3 => \N__34746\,
            lcout => n16,
            ltout => OPEN,
            carryin => n4719,
            carryout => n4720,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i11_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34743\,
            in2 => \_gnd_net_\,
            in3 => \N__34737\,
            lcout => n15,
            ltout => OPEN,
            carryin => n4720,
            carryout => n4721,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i12_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34734\,
            in2 => \_gnd_net_\,
            in3 => \N__34728\,
            lcout => n14,
            ltout => OPEN,
            carryin => n4721,
            carryout => n4722,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i13_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34725\,
            in2 => \_gnd_net_\,
            in3 => \N__34719\,
            lcout => n13,
            ltout => OPEN,
            carryin => n4722,
            carryout => n4723,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i14_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34716\,
            in2 => \_gnd_net_\,
            in3 => \N__34710\,
            lcout => n12,
            ltout => OPEN,
            carryin => n4723,
            carryout => n4724,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i15_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34890\,
            in2 => \_gnd_net_\,
            in3 => \N__34884\,
            lcout => n11,
            ltout => OPEN,
            carryin => n4724,
            carryout => n4725,
            clk => \N__37617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i16_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34881\,
            in2 => \_gnd_net_\,
            in3 => \N__34875\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => n4726,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i17_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34872\,
            in2 => \_gnd_net_\,
            in3 => \N__34866\,
            lcout => n9,
            ltout => OPEN,
            carryin => n4726,
            carryout => n4727,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i18_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34863\,
            in2 => \_gnd_net_\,
            in3 => \N__34857\,
            lcout => n8,
            ltout => OPEN,
            carryin => n4727,
            carryout => n4728,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i19_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34854\,
            in2 => \_gnd_net_\,
            in3 => \N__34848\,
            lcout => n7,
            ltout => OPEN,
            carryin => n4728,
            carryout => n4729,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i20_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34845\,
            in2 => \_gnd_net_\,
            in3 => \N__34839\,
            lcout => n6,
            ltout => OPEN,
            carryin => n4729,
            carryout => n4730,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i21_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34823\,
            in2 => \_gnd_net_\,
            in3 => \N__34812\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n4730,
            carryout => n4731,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i22_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34796\,
            in2 => \_gnd_net_\,
            in3 => \N__34785\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n4731,
            carryout => n4732,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i23_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \N__36237\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n4732,
            carryout => n4733,
            clk => \N__37619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i24_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36221\,
            in2 => \_gnd_net_\,
            in3 => \N__36210\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => n4734,
            clk => \N__37621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_523__i25_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36194\,
            in2 => \_gnd_net_\,
            in3 => \N__36207\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i3_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__36788\,
            in1 => \N__36150\,
            in2 => \N__36984\,
            in3 => \N__36896\,
            lcout => data_out_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i15_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__36110\,
            in1 => \N__36787\,
            in2 => \N__37065\,
            in3 => \N__36899\,
            lcout => data_out_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i121_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36000\,
            in1 => \N__35051\,
            in2 => \_gnd_net_\,
            in3 => \N__35099\,
            lcout => data_in_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_978_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36935\,
            in1 => \N__36390\,
            in2 => \_gnd_net_\,
            in3 => \N__36565\,
            lcout => \c0.n5409\,
            ltout => \c0.n5409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36507\,
            in1 => \N__35019\,
            in2 => \N__34974\,
            in3 => \N__34961\,
            lcout => n4_adj_1978,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_990_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36682\,
            in1 => \N__36391\,
            in2 => \_gnd_net_\,
            in3 => \N__36640\,
            lcout => n4_adj_1983,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i11_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__36945\,
            in1 => \N__36909\,
            in2 => \N__36282\,
            in3 => \N__36789\,
            lcout => data_out_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i12_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__36392\,
            in1 => \N__36910\,
            in2 => \N__37131\,
            in3 => \N__36790\,
            lcout => data_out_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36680\,
            in1 => \N__36642\,
            in2 => \N__36587\,
            in3 => \N__36567\,
            lcout => n8_adj_1984,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_981_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36506\,
            in1 => \N__36441\,
            in2 => \_gnd_net_\,
            in3 => \N__36399\,
            lcout => OPEN,
            ltout => \n7_adj_1985_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i26_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000011"
        )
    port map (
            in0 => \N__36341\,
            in1 => \N__36357\,
            in2 => \N__36351\,
            in3 => \N__37736\,
            lcout => data_out_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i0_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36317\,
            in2 => \_gnd_net_\,
            in3 => \N__36306\,
            lcout => data_0,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \c0.n4739\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i1_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36296\,
            in2 => \_gnd_net_\,
            in3 => \N__36285\,
            lcout => data_1,
            ltout => OPEN,
            carryin => \c0.n4739\,
            carryout => \c0.n4740\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i2_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36275\,
            in2 => \_gnd_net_\,
            in3 => \N__36264\,
            lcout => data_2,
            ltout => OPEN,
            carryin => \c0.n4740\,
            carryout => \c0.n4741\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i3_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37124\,
            in2 => \_gnd_net_\,
            in3 => \N__37113\,
            lcout => data_3,
            ltout => OPEN,
            carryin => \c0.n4741\,
            carryout => \c0.n4742\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i4_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37100\,
            in2 => \_gnd_net_\,
            in3 => \N__37089\,
            lcout => data_4,
            ltout => OPEN,
            carryin => \c0.n4742\,
            carryout => \c0.n4743\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i5_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37079\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => data_5,
            ltout => OPEN,
            carryin => \c0.n4743\,
            carryout => \c0.n4744\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i6_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37058\,
            in2 => \_gnd_net_\,
            in3 => \N__37047\,
            lcout => data_6,
            ltout => OPEN,
            carryin => \c0.n4744\,
            carryout => \c0.n4745\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i7_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37037\,
            in2 => \_gnd_net_\,
            in3 => \N__37026\,
            lcout => data_7,
            ltout => OPEN,
            carryin => \c0.n4745\,
            carryout => \c0.n4746\,
            clk => \N__37620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i8_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37019\,
            in2 => \_gnd_net_\,
            in3 => \N__37008\,
            lcout => data_8,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => \c0.n4747\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i9_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36998\,
            in2 => \_gnd_net_\,
            in3 => \N__36987\,
            lcout => data_9,
            ltout => OPEN,
            carryin => \c0.n4747\,
            carryout => \c0.n4748\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i10_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36980\,
            in2 => \_gnd_net_\,
            in3 => \N__36969\,
            lcout => data_10,
            ltout => OPEN,
            carryin => \c0.n4748\,
            carryout => \c0.n4749\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i11_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37880\,
            in2 => \_gnd_net_\,
            in3 => \N__37869\,
            lcout => data_11,
            ltout => OPEN,
            carryin => \c0.n4749\,
            carryout => \c0.n4750\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i12_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37856\,
            in2 => \_gnd_net_\,
            in3 => \N__37845\,
            lcout => data_12,
            ltout => OPEN,
            carryin => \c0.n4750\,
            carryout => \c0.n4751\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i13_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37832\,
            in2 => \_gnd_net_\,
            in3 => \N__37821\,
            lcout => data_13,
            ltout => OPEN,
            carryin => \c0.n4751\,
            carryout => \c0.n4752\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i14_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37808\,
            in2 => \_gnd_net_\,
            in3 => \N__37797\,
            lcout => data_14,
            ltout => OPEN,
            carryin => \c0.n4752\,
            carryout => \c0.n4753\,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_527__i15_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37790\,
            in2 => \_gnd_net_\,
            in3 => \N__37794\,
            lcout => data_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0___i20_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100101"
        )
    port map (
            in0 => \N__37776\,
            in1 => \N__37637\,
            in2 => \N__37764\,
            in3 => \N__37737\,
            lcout => data_out_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37623\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
