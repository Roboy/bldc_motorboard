// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Sep 12 19:16:24 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    inout PIN_1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    inout PIN_2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    input PIN_12 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    input PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    input PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    input PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire GND_net, VCC_net, LED_c, tx_o, tx2_o, tx_enable, tx2_enable, 
        rx_i;
    wire [25:0]blink_counter;   // verilog/TinyFPGA_B.v(64[14:27])
    wire [31:0]rand_data;   // verilog/TinyFPGA_B.v(77[14:23])
    wire [31:0]rand_setpoint;   // verilog/TinyFPGA_B.v(78[14:27])
    wire [7:0]byte_transmit_counter;   // coms.v(19[11:32])
    
    wire n3, n15593, n16629, n15562, n1, n3_adj_2406;
    wire [7:0]\data_out[9] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[8] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[6] ;   // coms.v(21[11:19])
    
    wire n10795, n10794;
    wire [7:0]\data_out[3] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    
    wire n17461, tx_active, n10793;
    wire [7:0]\UART_TRANSMITTER.state ;   // coms.v(277[13:18])
    
    wire rx_data_ready;
    wire [7:0]rx_data;   // coms.v(384[13:20])
    wire [7:0]\data_in[3] ;   // coms.v(388[12:19])
    wire [7:0]\data_in[2] ;   // coms.v(388[12:19])
    wire [7:0]\data_in[1] ;   // coms.v(388[12:19])
    wire [7:0]\data_in[0] ;   // coms.v(388[12:19])
    
    wire n16327, n15561, n10, n9460, n9462, n10_adj_2407;
    wire [7:0]\data_in_frame[7] ;   // coms.v(389[12:25])
    wire [7:0]\data_in_frame[6] ;   // coms.v(389[12:25])
    wire [7:0]\data_in_frame[0] ;   // coms.v(389[12:25])
    wire [7:0]\data_out_frame2[18] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[17] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[16] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[15] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[14] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[13] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[12] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[11] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[10] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[9] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[8] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[7] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[6] ;   // coms.v(390[12:27])
    wire [7:0]\data_out_frame2[5] ;   // coms.v(390[12:27])
    
    wire n6;
    wire [31:0]\FRAME_MATCHER.state ;   // coms.v(419[11:16])
    
    wire n10792, n10791, n4, n10790, n10789, n10788, n10787, n10786, 
        n8730, n3_adj_2408, n16795, n16473, n14060, n16863, n10374, 
        n10785, n7866, n13, n10784, n17458, n17457, n15592, n10783, 
        n10782, n4_adj_2409, n10781, n13440, n10780, n10779, n10778, 
        n10777, data_out_9__2__N_367, n15560, n15591, n16671, n17544, 
        n5, n10776, n10775, n10774, n12, n10773, n10772, n17542, 
        n15539, n10373, n10771, n15590, n127, n10770, n10372, 
        n9929, n17537, n10769, n15701, n10768, n15589, n10767, 
        n10766, n10765, n10764, n10763, n10762, n10761, n10760, 
        n7198, n10759, n10371, n119, n118, n117, n116, data_out_10__7__N_110, 
        n10758, n10757, n10756, n10755, n10754, n10753, n10752, 
        n10751, n10750, n10749, n10748, n10747, n10746, n10745, 
        n10744, n10743, n10742, n10741, n10740, n13082, n10739, 
        n10738, n10737, n10736, n10735, n10734, n10733, n10732, 
        n9361, n10731, n10730, n10729, n10728, n10727, n10726, 
        n115, n10725, n114, n13276, n31, n10714, n15538, n15588, 
        n113, n165, n164, n163, n162, n161, n160, n159, n158, 
        n157, n156, n155, n15537, n15536, n15535, n17298, n16856, 
        n16649, n10698, n10697, n12_adj_2410, n10695, n112, n10693, 
        n10692, n10691, n16467, n17144, n1651, n111, n110, n10031, 
        n9403, n1716, n4_adj_2411, n16509, n15559, n15587, n2275;
    wire [31:0]\FRAME_MATCHER.state_31__N_1440 ;
    
    wire n10836, n10835, n10834, n10833, n10832, n10_adj_2412, n16896, 
        n15586, n15558, n12933, n17, n16844, n10_adj_2413, n16463, 
        n16852, n10_adj_2414, n15557, n13510, n16824, n16797, n16623, 
        n14, n10_adj_2415, n15585, n15556, n16607, n17504, n15584, 
        n16459, n15555, n15534, n15583, n15582, n15533, n15532, 
        n15581, n15580, n15531, n15554, n15553, n15530, n15579, 
        n15552, n15551, n15550, n15578, n15577, n15576, n10690, 
        n16828, n10689, n10688, n10687, n10686, n10685, n53, n10684, 
        n10683, n10682, n10681, n9937, n10680, n10679, n10678, 
        n10677, n10676, n10675, n10674, n10673, n10672, n10671, 
        n5029, n10670, n10669, n10668, n9453, n4445, n10667, n10666, 
        n10665, n17494, n10664, n15549, n15575, n10663, n15548, 
        n15574, n15529, n15547, n15528, n10662, n15614, n15546, 
        n10661, n15573, n10660, n10659, n15613, n10658, n10367, 
        n16483, n15612, n10366, n15611, n15610, n15609, n10365, 
        n15572, n15608, n15607, n15571, n15570, n15569, n15606, 
        n15605, n2652, n16625, n10364, n15568, n10362, n15567, 
        n15545, n15544, n15604, n15543, n15603, n16627, n10361, 
        n17_adj_2416, n16854, n4_adj_2417, n3977, n26, n9, n8, 
        n7, n127_adj_2418, n17641, n17640, n10831, n10197, n10803, 
        n10804, n10805, n10806, n10830, n10635, n10829, n10807, 
        n10808, n10810, n10631, n10809, n10811, n10812, n10796, 
        n10797, n15837, n10828, n10813, n16857, n10814, n20, n10798, 
        n17484, n10815, n10625, n10624, n19, n15, n10623, n16893, 
        n10622, n10621, n10620, n10619, n12_adj_2419, n16859, n11, 
        n10817, n10816, n10799, n10800, n10801, n10802, n10141, 
        n10_adj_2420, n10607, n16855, n10599, n10598, n10597, n10596, 
        n16775, n10592, n10591, n10590, n10360, n10359, n10358, 
        n10589, n10357, n10355, n17398, n10588, n10587, n6_adj_2421, 
        n10585, n10584, n10583, n10582, n10581, n17_adj_2422, n10580, 
        n10579, n17636, n25, n24, n23, n22, n491, n10578, n15689, 
        n10577, n17479, n2547, n17634, n10_adj_2423, n21, n445, 
        n18, n16, n14_adj_2424, n16567, n10576, n17631, n10575, 
        n10574, n9472, n17629, n16469, n16479, n16569, n16651, 
        n16673, n16517, n16571, n17395, n16573, n16575, n16577, 
        n16675, n16677, n10055, n17260, n16886, n154, n153, n152, 
        n151, n150, n149, n148, n147, n146, n145, n144, n143, 
        n142, n141, n140, n139, n138, n137, n136, n135, n134, 
        n16683, n10_adj_2425, n17194, n10_adj_2426, n10_adj_2427, 
        n10433, n10432, n17230, n10431, n15566, n17299, n16860, 
        n16547, n9357, n10430, n17222, n17602, n10429, n17601, 
        n10428;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n10827, n10826, n10825, n10427, n10426, n135_adj_2428, 
        n134_adj_2429, n133, n132, n131, n130, n10425, n10423, 
        n16259, r_Rx_Data;
    wire [7:0]r_Clock_Count_adj_2504;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index_adj_2505;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_adj_2506;   // verilog/uart_rx.v(36[17:26])
    
    wire n9452, n10824, n10823, n10822, n15602, n129, n128, n127_adj_2442, 
        n126, n125, n124, n123, n122, n16477;
    wire [2:0]r_SM_Main_adj_2509;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_2510;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_2511;   // verilog/uart_tx.v(33[16:27])
    
    wire n15542, n29;
    wire [2:0]r_SM_Main_2__N_2033_adj_2515;
    
    wire n10821, n10820, n10819, n121, n120, n10399, n10398, n9445, 
        n15601, n15565, n16681, n15600, n4_adj_2458, n15541, n15564, 
        n10396, n8_adj_2459, n17397, n10392, n15599, n17573, n15598, 
        n17394, n18137, n18044, n33, n41, n38, n18038, n35, 
        n17140, n17570, n4_adj_2460, n6_adj_2461, n16776, n18032, 
        n17162, n18026, n17208, n16897, n16810, n134_adj_2462, n135_adj_2463, 
        n136_adj_2464, n137_adj_2465, n138_adj_2466, n139_adj_2467, 
        n140_adj_2468, n141_adj_2469, n142_adj_2470, n143_adj_2471, 
        n144_adj_2472, n145_adj_2473, n146_adj_2474, n147_adj_2475, 
        n148_adj_2476, n149_adj_2477, n150_adj_2478, n151_adj_2479, 
        n152_adj_2480, n153_adj_2481, n154_adj_2482, n155_adj_2483, 
        n156_adj_2484, n157_adj_2485, n158_adj_2486, n159_adj_2487, 
        n160_adj_2488, n161_adj_2489, n162_adj_2490, n163_adj_2491, 
        n164_adj_2492, n165_adj_2493, n9435, n17567, n16255, n15540, 
        n9406, n9477, n16858, n9358, n15597, n15563, n16515, n16867, 
        n16853, n17834, n17154, n15596, n10818, n8828, n16817, 
        n15595, n15594;
    
    VCC i2 (.Y(VCC_net));
    SB_IO tx2_output (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx2_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx2_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx2_output.PIN_TYPE = 6'b101001;
    defparam tx2_output.PULLUP = 1'b1;
    defparam tx2_output.NEG_TRIGGER = 1'b0;
    defparam tx2_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO rx_input (.PACKAGE_PIN(PIN_2), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(rx_i)) /* synthesis lattice_noprune=1, syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam rx_input.PIN_TYPE = 6'b000001;
    defparam rx_input.PULLUP = 1'b1;
    defparam rx_input.NEG_TRIGGER = 1'b0;
    defparam rx_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_1), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i43_4_lut (.I0(n17834), .I1(n4445), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(n17162), .O(n16259));   // coms.v(280[12] 380[6])
    defparam i43_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i31_3_lut (.I0(r_Clock_Count_adj_2510[0]), .I1(n17544), .I2(r_SM_Main_adj_2509[2]), 
            .I3(GND_net), .O(n16623));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n16795), .I1(n9452), .I2(n17), .I3(n2275), 
            .O(n16775));   // coms.v(426[12] 547[6])
    defparam i1_4_lut.LUT_INIT = 16'hf5f7;
    SB_LUT4 i8214_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n16893), 
            .I3(GND_net), .O(n10574));   // coms.v(426[12] 547[6])
    defparam i8214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8451_3_lut (.I0(\data_out_frame2[15] [6]), .I1(rand_data[14]), 
            .I2(n10197), .I3(GND_net), .O(n10811));   // coms.v(426[12] 547[6])
    defparam i8451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8215_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n16893), 
            .I3(GND_net), .O(n10575));   // coms.v(426[12] 547[6])
    defparam i8215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8216_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n16893), 
            .I3(GND_net), .O(n10576));   // coms.v(426[12] 547[6])
    defparam i8216_3_lut.LUT_INIT = 16'hacac;
    SB_DFF rand_setpoint_2351__i0 (.Q(rand_setpoint[0]), .C(CLK_c), .D(n165));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF blink_counter_2352__i0 (.Q(n26), .C(CLK_c), .D(n135_adj_2428));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i8217_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n16897), 
            .I3(GND_net), .O(n10577));   // coms.v(426[12] 547[6])
    defparam i8217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8369_3_lut (.I0(\data_out_frame2[5] [4]), .I1(rand_data[28]), 
            .I2(n10197), .I3(GND_net), .O(n10729));   // coms.v(426[12] 547[6])
    defparam i8369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8218_3_lut (.I0(tx_o), .I1(n3_adj_2406), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n10578));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8219_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n4_adj_2458), .O(n10579));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8219_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i8370_3_lut (.I0(\data_out_frame2[5] [5]), .I1(rand_data[29]), 
            .I2(n10197), .I3(GND_net), .O(n10730));   // coms.v(426[12] 547[6])
    defparam i8370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut (.I0(n17542), .I1(r_Clock_Count[0]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16625));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8371_3_lut (.I0(\data_out_frame2[5] [6]), .I1(rand_data[30]), 
            .I2(n10197), .I3(GND_net), .O(n10731));   // coms.v(426[12] 547[6])
    defparam i8371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8372_3_lut (.I0(\data_out_frame2[5] [7]), .I1(rand_data[31]), 
            .I2(n10197), .I3(GND_net), .O(n10732));   // coms.v(426[12] 547[6])
    defparam i8372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_21_lut (.I0(GND_net), .I1(rand_data[19]), 
            .I2(rand_setpoint[19]), .I3(n15577), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8417_3_lut (.I0(\data_out_frame2[11] [4]), .I1(rand_data[12]), 
            .I2(n10197), .I3(GND_net), .O(n10777));   // coms.v(426[12] 547[6])
    defparam i8417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_765 (.I0(n127_adj_2418), .I1(n1716), .I2(n12933), 
            .I3(n16775), .O(n14));   // coms.v(426[12] 547[6])
    defparam i1_4_lut_adj_765.LUT_INIT = 16'h8808;
    SB_CARRY rand_setpoint_2351_add_4_21 (.CI(n15577), .I0(rand_data[19]), 
            .I1(rand_setpoint[19]), .CO(n15578));
    SB_LUT4 i1_4_lut_adj_766 (.I0(n17208), .I1(n3977), .I2(n14), .I3(n12933), 
            .O(n16797));   // coms.v(426[12] 547[6])
    defparam i1_4_lut_adj_766.LUT_INIT = 16'hf5fd;
    SB_LUT4 i8220_4_lut (.I0(r_SM_Main[2]), .I1(n5), .I2(n14060), .I3(r_SM_Main[0]), 
            .O(n10580));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8220_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 rand_setpoint_2351_add_4_20_lut (.I0(GND_net), .I1(rand_data[18]), 
            .I2(rand_setpoint[18]), .I3(n15576), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_27 (.CI(n15552), .I0(GND_net), .I1(rand_data[25]), 
            .CO(n15553));
    SB_LUT4 i8221_4_lut (.I0(r_SM_Main_adj_2506[2]), .I1(n1), .I2(n13440), 
            .I3(r_SM_Main_adj_2506[1]), .O(n10581));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8221_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i31_3_lut_adj_767 (.I0(r_Clock_Count_adj_2510[1]), .I1(n17504), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16677));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut_adj_767.LUT_INIT = 16'hacac;
    SB_LUT4 rand_data_2350_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[9]), 
            .I3(n15536), .O(n156_adj_2484)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8222_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n16893), 
            .I3(GND_net), .O(n10582));   // coms.v(426[12] 547[6])
    defparam i8222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8223_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n16893), 
            .I3(GND_net), .O(n10583));   // coms.v(426[12] 547[6])
    defparam i8223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8224_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n16893), 
            .I3(GND_net), .O(n10584));   // coms.v(426[12] 547[6])
    defparam i8224_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rand_setpoint_2351_add_4_20 (.CI(n15576), .I0(rand_data[18]), 
            .I1(rand_setpoint[18]), .CO(n15577));
    SB_LUT4 i8225_3_lut (.I0(tx2_o), .I1(n3), .I2(r_SM_Main_adj_2509[2]), 
            .I3(GND_net), .O(n10585));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8225_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14702_3_lut (.I0(n12_adj_2410), .I1(r_SM_Main_adj_2509[1]), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n17140));
    defparam i14702_3_lut.LUT_INIT = 16'hd5d5;
    SB_LUT4 i8373_3_lut (.I0(\data_out_frame2[6] [0]), .I1(rand_data[16]), 
            .I2(n10197), .I3(GND_net), .O(n10733));   // coms.v(426[12] 547[6])
    defparam i8373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14847_4_lut (.I0(n15837), .I1(n9929), .I2(n17140), .I3(n9403), 
            .O(n16817));
    defparam i14847_4_lut.LUT_INIT = 16'h1505;
    SB_LUT4 i8227_4_lut (.I0(r_SM_Main_adj_2509[2]), .I1(n7866), .I2(r_SM_Main_2__N_2033_adj_2515[1]), 
            .I3(r_SM_Main_adj_2509[0]), .O(n10587));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8227_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 rand_data_2350_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[24]), 
            .I3(n15551), .O(n141_adj_2469)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_768 (.I0(n17208), .I1(n8828), .I2(n16776), .I3(\FRAME_MATCHER.state [0]), 
            .O(n16327));   // coms.v(426[12] 547[6])
    defparam i1_4_lut_adj_768.LUT_INIT = 16'hf575;
    SB_LUT4 i8452_3_lut (.I0(\data_out_frame2[15] [7]), .I1(rand_data[15]), 
            .I2(n10197), .I3(GND_net), .O(n10812));   // coms.v(426[12] 547[6])
    defparam i8452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14770_3_lut (.I0(n31), .I1(\FRAME_MATCHER.state [1]), .I2(n9445), 
            .I3(GND_net), .O(n17208));
    defparam i14770_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i8228_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n16893), 
            .I3(GND_net), .O(n10588));   // coms.v(426[12] 547[6])
    defparam i8228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8229_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n16896), 
            .I3(GND_net), .O(n10589));   // coms.v(426[12] 547[6])
    defparam i8229_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8230_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n16896), 
            .I3(GND_net), .O(n10590));   // coms.v(426[12] 547[6])
    defparam i8230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8393_3_lut (.I0(\data_out_frame2[8] [4]), .I1(rand_data[4]), 
            .I2(n10197), .I3(GND_net), .O(n10753));   // coms.v(426[12] 547[6])
    defparam i8393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8231_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n16896), 
            .I3(GND_net), .O(n10591));   // coms.v(426[12] 547[6])
    defparam i8231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8232_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n16896), 
            .I3(GND_net), .O(n10592));   // coms.v(426[12] 547[6])
    defparam i8232_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8236_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n16896), 
            .I3(GND_net), .O(n10596));   // coms.v(426[12] 547[6])
    defparam i8236_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8237_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n16896), 
            .I3(GND_net), .O(n10597));   // coms.v(426[12] 547[6])
    defparam i8237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8418_3_lut (.I0(\data_out_frame2[11] [5]), .I1(rand_data[13]), 
            .I2(n10197), .I3(GND_net), .O(n10778));   // coms.v(426[12] 547[6])
    defparam i8418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8453_3_lut (.I0(\data_out_frame2[16] [0]), .I1(rand_data[0]), 
            .I2(n10197), .I3(GND_net), .O(n10813));   // coms.v(426[12] 547[6])
    defparam i8453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8394_3_lut (.I0(\data_out_frame2[8] [5]), .I1(rand_data[5]), 
            .I2(n10197), .I3(GND_net), .O(n10754));   // coms.v(426[12] 547[6])
    defparam i8394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8238_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n16896), 
            .I3(GND_net), .O(n10598));   // coms.v(426[12] 547[6])
    defparam i8238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8374_3_lut (.I0(\data_out_frame2[6] [1]), .I1(rand_data[17]), 
            .I2(n10197), .I3(GND_net), .O(n10734));   // coms.v(426[12] 547[6])
    defparam i8374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8454_3_lut (.I0(\data_out_frame2[16] [1]), .I1(rand_data[1]), 
            .I2(n10197), .I3(GND_net), .O(n10814));   // coms.v(426[12] 547[6])
    defparam i8454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8375_3_lut (.I0(\data_out_frame2[6] [2]), .I1(rand_data[18]), 
            .I2(n10197), .I3(GND_net), .O(n10735));   // coms.v(426[12] 547[6])
    defparam i8375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8395_3_lut (.I0(\data_out_frame2[8] [6]), .I1(rand_data[6]), 
            .I2(n10197), .I3(GND_net), .O(n10755));   // coms.v(426[12] 547[6])
    defparam i8395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_19_lut (.I0(GND_net), .I1(rand_data[17]), 
            .I2(rand_setpoint[17]), .I3(n15575), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8239_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n16896), 
            .I3(GND_net), .O(n10599));   // coms.v(426[12] 547[6])
    defparam i8239_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rand_data_2350_add_4_26 (.CI(n15551), .I0(GND_net), .I1(rand_data[24]), 
            .CO(n15552));
    SB_LUT4 i8376_3_lut (.I0(\data_out_frame2[6] [3]), .I1(rand_data[19]), 
            .I2(n10197), .I3(GND_net), .O(n10736));   // coms.v(426[12] 547[6])
    defparam i8376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8455_3_lut (.I0(\data_out_frame2[16] [2]), .I1(rand_data[2]), 
            .I2(n10197), .I3(GND_net), .O(n10815));   // coms.v(426[12] 547[6])
    defparam i8455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8377_3_lut (.I0(\data_out_frame2[6] [4]), .I1(rand_data[20]), 
            .I2(n10197), .I3(GND_net), .O(n10737));   // coms.v(426[12] 547[6])
    defparam i8377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8378_3_lut (.I0(\data_out_frame2[6] [5]), .I1(rand_data[21]), 
            .I2(n10197), .I3(GND_net), .O(n10738));   // coms.v(426[12] 547[6])
    defparam i8378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8379_3_lut (.I0(\data_out_frame2[6] [6]), .I1(rand_data[22]), 
            .I2(n10197), .I3(GND_net), .O(n10739));   // coms.v(426[12] 547[6])
    defparam i8379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8380_3_lut (.I0(\data_out_frame2[6] [7]), .I1(rand_data[23]), 
            .I2(n10197), .I3(GND_net), .O(n10740));   // coms.v(426[12] 547[6])
    defparam i8380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8032_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n16893), 
            .I3(GND_net), .O(n10392));   // coms.v(426[12] 547[6])
    defparam i8032_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8434_3_lut (.I0(\data_out_frame2[13] [5]), .I1(rand_data[29]), 
            .I2(n10197), .I3(GND_net), .O(n10794));   // coms.v(426[12] 547[6])
    defparam i8434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8067_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n13082), 
            .I3(n9472), .O(n10427));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8067_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i8068_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n13082), 
            .I3(n9477), .O(n10428));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8068_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i8069_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_2417), 
            .I3(n9472), .O(n10429));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8069_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8070_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_2417), 
            .I3(n9477), .O(n10430));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8070_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8071_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_2460), 
            .I3(n9472), .O(n10431));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8071_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8072_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_2460), 
            .I3(n9477), .O(n10432));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8072_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8073_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_2409), 
            .I3(n9472), .O(n10433));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8073_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8381_3_lut (.I0(\data_out_frame2[7] [0]), .I1(rand_data[8]), 
            .I2(n10197), .I3(GND_net), .O(n10741));   // coms.v(426[12] 547[6])
    defparam i8381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8382_3_lut (.I0(\data_out_frame2[7] [1]), .I1(rand_data[9]), 
            .I2(n10197), .I3(GND_net), .O(n10742));   // coms.v(426[12] 547[6])
    defparam i8382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14960_3_lut (.I0(r_Tx_Data[5]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n17398));
    defparam i14960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14959_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[6]), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n17397));
    defparam i14959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8463_3_lut (.I0(\data_out_frame2[17] [2]), .I1(rand_data[10]), 
            .I2(n10197), .I3(GND_net), .O(n10823));   // coms.v(426[12] 547[6])
    defparam i8463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8396_3_lut (.I0(\data_out_frame2[8] [7]), .I1(rand_data[7]), 
            .I2(n10197), .I3(GND_net), .O(n10756));   // coms.v(426[12] 547[6])
    defparam i8396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8464_3_lut (.I0(\data_out_frame2[17] [3]), .I1(rand_data[11]), 
            .I2(n10197), .I3(GND_net), .O(n10824));   // coms.v(426[12] 547[6])
    defparam i8464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8456_3_lut (.I0(\data_out_frame2[16] [3]), .I1(rand_data[3]), 
            .I2(n10197), .I3(GND_net), .O(n10816));   // coms.v(426[12] 547[6])
    defparam i8456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8397_3_lut (.I0(\data_out_frame2[9] [0]), .I1(rand_data[24]), 
            .I2(n10197), .I3(GND_net), .O(n10757));   // coms.v(426[12] 547[6])
    defparam i8397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8472_3_lut (.I0(\data_out_frame2[18] [3]), .I1(rand_data[3]), 
            .I2(n10197), .I3(GND_net), .O(n10832));   // coms.v(426[12] 547[6])
    defparam i8472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8473_3_lut (.I0(\data_out_frame2[18] [4]), .I1(rand_data[4]), 
            .I2(n10197), .I3(GND_net), .O(n10833));   // coms.v(426[12] 547[6])
    defparam i8473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8419_3_lut (.I0(\data_out_frame2[11] [6]), .I1(rand_data[14]), 
            .I2(n10197), .I3(GND_net), .O(n10779));   // coms.v(426[12] 547[6])
    defparam i8419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8474_3_lut (.I0(\data_out_frame2[18] [5]), .I1(rand_data[5]), 
            .I2(n10197), .I3(GND_net), .O(n10834));   // coms.v(426[12] 547[6])
    defparam i8474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8420_3_lut (.I0(\data_out_frame2[11] [7]), .I1(rand_data[15]), 
            .I2(n10197), .I3(GND_net), .O(n10780));   // coms.v(426[12] 547[6])
    defparam i8420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8475_3_lut (.I0(\data_out_frame2[18] [6]), .I1(rand_data[6]), 
            .I2(n10197), .I3(GND_net), .O(n10835));   // coms.v(426[12] 547[6])
    defparam i8475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8383_3_lut (.I0(\data_out_frame2[7] [2]), .I1(rand_data[10]), 
            .I2(n10197), .I3(GND_net), .O(n10743));   // coms.v(426[12] 547[6])
    defparam i8383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8476_3_lut (.I0(\data_out_frame2[18] [7]), .I1(rand_data[7]), 
            .I2(n10197), .I3(GND_net), .O(n10836));   // coms.v(426[12] 547[6])
    defparam i8476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8384_3_lut (.I0(\data_out_frame2[7] [3]), .I1(rand_data[11]), 
            .I2(n10197), .I3(GND_net), .O(n10744));   // coms.v(426[12] 547[6])
    defparam i8384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8385_3_lut (.I0(\data_out_frame2[7] [4]), .I1(rand_data[12]), 
            .I2(n10197), .I3(GND_net), .O(n10745));   // coms.v(426[12] 547[6])
    defparam i8385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8386_3_lut (.I0(\data_out_frame2[7] [5]), .I1(rand_data[13]), 
            .I2(n10197), .I3(GND_net), .O(n10746));   // coms.v(426[12] 547[6])
    defparam i8386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8436_3_lut (.I0(\data_out_frame2[13] [7]), .I1(rand_data[31]), 
            .I2(n10197), .I3(GND_net), .O(n10796));   // coms.v(426[12] 547[6])
    defparam i8436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8387_3_lut (.I0(\data_out_frame2[7] [6]), .I1(rand_data[14]), 
            .I2(n10197), .I3(GND_net), .O(n10747));   // coms.v(426[12] 547[6])
    defparam i8387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8437_3_lut (.I0(\data_out_frame2[14] [0]), .I1(rand_data[16]), 
            .I2(n10197), .I3(GND_net), .O(n10797));   // coms.v(426[12] 547[6])
    defparam i8437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8388_3_lut (.I0(\data_out_frame2[7] [7]), .I1(rand_data[15]), 
            .I2(n10197), .I3(GND_net), .O(n10748));   // coms.v(426[12] 547[6])
    defparam i8388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8438_3_lut (.I0(\data_out_frame2[14] [1]), .I1(rand_data[17]), 
            .I2(n10197), .I3(GND_net), .O(n10798));   // coms.v(426[12] 547[6])
    defparam i8438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8389_3_lut (.I0(\data_out_frame2[8] [0]), .I1(rand_data[0]), 
            .I2(n10197), .I3(GND_net), .O(n10749));   // coms.v(426[12] 547[6])
    defparam i8389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8439_3_lut (.I0(\data_out_frame2[14] [2]), .I1(rand_data[18]), 
            .I2(n10197), .I3(GND_net), .O(n10799));   // coms.v(426[12] 547[6])
    defparam i8439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8390_3_lut (.I0(\data_out_frame2[8] [1]), .I1(rand_data[1]), 
            .I2(n10197), .I3(GND_net), .O(n10750));   // coms.v(426[12] 547[6])
    defparam i8390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8440_3_lut (.I0(\data_out_frame2[14] [3]), .I1(rand_data[19]), 
            .I2(n10197), .I3(GND_net), .O(n10800));   // coms.v(426[12] 547[6])
    defparam i8440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8391_3_lut (.I0(\data_out_frame2[8] [2]), .I1(rand_data[2]), 
            .I2(n10197), .I3(GND_net), .O(n10751));   // coms.v(426[12] 547[6])
    defparam i8391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8441_3_lut (.I0(\data_out_frame2[14] [4]), .I1(rand_data[20]), 
            .I2(n10197), .I3(GND_net), .O(n10801));   // coms.v(426[12] 547[6])
    defparam i8441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8392_3_lut (.I0(\data_out_frame2[8] [3]), .I1(rand_data[3]), 
            .I2(n10197), .I3(GND_net), .O(n10752));   // coms.v(426[12] 547[6])
    defparam i8392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8442_3_lut (.I0(\data_out_frame2[14] [5]), .I1(rand_data[21]), 
            .I2(n10197), .I3(GND_net), .O(n10802));   // coms.v(426[12] 547[6])
    defparam i8442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8443_3_lut (.I0(\data_out_frame2[14] [6]), .I1(rand_data[22]), 
            .I2(n10197), .I3(GND_net), .O(n10803));   // coms.v(426[12] 547[6])
    defparam i8443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8444_3_lut (.I0(\data_out_frame2[14] [7]), .I1(rand_data[23]), 
            .I2(n10197), .I3(GND_net), .O(n10804));   // coms.v(426[12] 547[6])
    defparam i8444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8445_3_lut (.I0(\data_out_frame2[15] [0]), .I1(rand_data[8]), 
            .I2(n10197), .I3(GND_net), .O(n10805));   // coms.v(426[12] 547[6])
    defparam i8445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8446_3_lut (.I0(\data_out_frame2[15] [1]), .I1(rand_data[9]), 
            .I2(n10197), .I3(GND_net), .O(n10806));   // coms.v(426[12] 547[6])
    defparam i8446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8447_3_lut (.I0(\data_out_frame2[15] [2]), .I1(rand_data[10]), 
            .I2(n10197), .I3(GND_net), .O(n10807));   // coms.v(426[12] 547[6])
    defparam i8447_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_19 (.CI(n15575), .I0(rand_data[17]), 
            .I1(rand_setpoint[17]), .CO(n15576));
    SB_LUT4 i8421_3_lut (.I0(\data_out_frame2[12] [0]), .I1(rand_data[0]), 
            .I2(n10197), .I3(GND_net), .O(n10781));   // coms.v(426[12] 547[6])
    defparam i8421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8422_3_lut (.I0(\data_out_frame2[12] [1]), .I1(rand_data[1]), 
            .I2(n10197), .I3(GND_net), .O(n10782));   // coms.v(426[12] 547[6])
    defparam i8422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8398_3_lut (.I0(\data_out_frame2[9] [1]), .I1(rand_data[25]), 
            .I2(n10197), .I3(GND_net), .O(n10758));   // coms.v(426[12] 547[6])
    defparam i8398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8399_3_lut (.I0(\data_out_frame2[9] [2]), .I1(rand_data[26]), 
            .I2(n10197), .I3(GND_net), .O(n10759));   // coms.v(426[12] 547[6])
    defparam i8399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[23]), 
            .I3(n15550), .O(n142_adj_2470)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8423_3_lut (.I0(\data_out_frame2[12] [2]), .I1(rand_data[2]), 
            .I2(n10197), .I3(GND_net), .O(n10783));   // coms.v(426[12] 547[6])
    defparam i8423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8424_3_lut (.I0(\data_out_frame2[12] [3]), .I1(rand_data[3]), 
            .I2(n10197), .I3(GND_net), .O(n10784));   // coms.v(426[12] 547[6])
    defparam i8424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8400_3_lut (.I0(\data_out_frame2[9] [3]), .I1(rand_data[27]), 
            .I2(n10197), .I3(GND_net), .O(n10760));   // coms.v(426[12] 547[6])
    defparam i8400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14956_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[2]), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n17394));
    defparam i14956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14957_3_lut (.I0(r_Tx_Data[1]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n17395));
    defparam i14957_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2350_add_4_25 (.CI(n15550), .I0(GND_net), .I1(rand_data[23]), 
            .CO(n15551));
    SB_LUT4 i8425_3_lut (.I0(\data_out_frame2[12] [4]), .I1(rand_data[4]), 
            .I2(n10197), .I3(GND_net), .O(n10785));   // coms.v(426[12] 547[6])
    defparam i8425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8401_3_lut (.I0(\data_out_frame2[9] [4]), .I1(rand_data[28]), 
            .I2(n10197), .I3(GND_net), .O(n10761));   // coms.v(426[12] 547[6])
    defparam i8401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_4_lut (.I0(n18026), .I1(n10_adj_2426), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2407));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut (.I0(r_Tx_Data[4]), .I1(n10_adj_2407), .I2(n8730), 
            .I3(byte_transmit_counter[4]), .O(n16681));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8426_3_lut (.I0(\data_out_frame2[12] [5]), .I1(rand_data[5]), 
            .I2(n10197), .I3(GND_net), .O(n10786));   // coms.v(426[12] 547[6])
    defparam i8426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_4_lut_adj_769 (.I0(n18032), .I1(n10_adj_2425), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_4_lut_adj_769.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_770 (.I0(r_Tx_Data[5]), .I1(n10), .I2(n8730), 
            .I3(byte_transmit_counter[4]), .O(n16683));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i23_4_lut_adj_770.LUT_INIT = 16'h0aca;
    SB_LUT4 i24_4_lut_adj_771 (.I0(n18038), .I1(n10_adj_2427), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2413));   // coms.v(19[11:32])
    defparam i24_4_lut_adj_771.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut_adj_772 (.I0(r_Tx_Data[6]), .I1(n10_adj_2413), .I2(n8730), 
            .I3(byte_transmit_counter[4]), .O(n16629));   // coms.v(19[11:32])
    defparam i23_4_lut_adj_772.LUT_INIT = 16'h0aca;
    SB_LUT4 i8402_3_lut (.I0(\data_out_frame2[9] [5]), .I1(rand_data[29]), 
            .I2(n10197), .I3(GND_net), .O(n10762));   // coms.v(426[12] 547[6])
    defparam i8402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_4_lut_adj_773 (.I0(n18044), .I1(n10_adj_2423), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n10_adj_2414));   // coms.v(19[11:32])
    defparam i24_4_lut_adj_773.LUT_INIT = 16'h0aca;
    SB_LUT4 i8427_3_lut (.I0(\data_out_frame2[12] [6]), .I1(rand_data[6]), 
            .I2(n10197), .I3(GND_net), .O(n10787));   // coms.v(426[12] 547[6])
    defparam i8427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_adj_774 (.I0(r_Tx_Data[7]), .I1(n10_adj_2414), .I2(n8730), 
            .I3(byte_transmit_counter[4]), .O(n16627));   // coms.v(19[11:32])
    defparam i23_4_lut_adj_774.LUT_INIT = 16'h0aca;
    SB_LUT4 i8448_3_lut (.I0(\data_out_frame2[15] [3]), .I1(rand_data[11]), 
            .I2(n10197), .I3(GND_net), .O(n10808));   // coms.v(426[12] 547[6])
    defparam i8448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8449_3_lut (.I0(\data_out_frame2[15] [4]), .I1(rand_data[12]), 
            .I2(n10197), .I3(GND_net), .O(n10809));   // coms.v(426[12] 547[6])
    defparam i8449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8428_3_lut (.I0(\data_out_frame2[12] [7]), .I1(rand_data[7]), 
            .I2(n10197), .I3(GND_net), .O(n10788));   // coms.v(426[12] 547[6])
    defparam i8428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8066_4_lut (.I0(n10425), .I1(r_Bit_Index_adj_2505[1]), .I2(r_Bit_Index_adj_2505[0]), 
            .I3(n17260), .O(n10426));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8066_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i8063_4_lut (.I0(n10425), .I1(r_Bit_Index_adj_2505[2]), .I2(n4_adj_2411), 
            .I3(n17260), .O(n10423));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8063_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i8435_3_lut (.I0(\data_out_frame2[13] [6]), .I1(rand_data[30]), 
            .I2(n10197), .I3(GND_net), .O(n10795));   // coms.v(426[12] 547[6])
    defparam i8435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[22]), 
            .I3(n15549), .O(n143_adj_2471)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_11 (.CI(n15536), .I0(GND_net), .I1(rand_data[9]), 
            .CO(n15537));
    SB_LUT4 rand_setpoint_2351_add_4_18_lut (.I0(GND_net), .I1(rand_data[16]), 
            .I2(rand_setpoint[16]), .I3(n15574), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_24 (.CI(n15549), .I0(GND_net), .I1(rand_data[22]), 
            .CO(n15550));
    SB_CARRY rand_setpoint_2351_add_4_18 (.CI(n15574), .I0(rand_data[16]), 
            .I1(rand_setpoint[16]), .CO(n15575));
    SB_LUT4 i8403_3_lut (.I0(\data_out_frame2[9] [6]), .I1(rand_data[30]), 
            .I2(n10197), .I3(GND_net), .O(n10763));   // coms.v(426[12] 547[6])
    defparam i8403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8404_3_lut (.I0(\data_out_frame2[9] [7]), .I1(rand_data[31]), 
            .I2(n10197), .I3(GND_net), .O(n10764));   // coms.v(426[12] 547[6])
    defparam i8404_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 blink_counter_2352_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[25]), .I3(n15614), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2352_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[24]), .I3(n15613), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[8]), 
            .I3(n15535), .O(n157_adj_2485)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_26 (.CI(n15613), .I0(GND_net), .I1(blink_counter[24]), 
            .CO(n15614));
    SB_LUT4 blink_counter_2352_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[23]), .I3(n15612), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_25 (.CI(n15612), .I0(GND_net), .I1(blink_counter[23]), 
            .CO(n15613));
    SB_LUT4 blink_counter_2352_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[22]), .I3(n15611), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY blink_counter_2352_add_4_24 (.CI(n15611), .I0(GND_net), .I1(blink_counter[22]), 
            .CO(n15612));
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /media/external/iCEcube2/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 blink_counter_2352_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[21]), .I3(n15610), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_23 (.CI(n15610), .I0(GND_net), .I1(blink_counter[21]), 
            .CO(n15611));
    SB_LUT4 blink_counter_2352_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_2421), .I3(n15609), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_22 (.CI(n15609), .I0(GND_net), .I1(n6_adj_2421), 
            .CO(n15610));
    SB_LUT4 rand_setpoint_2351_add_4_17_lut (.I0(GND_net), .I1(rand_data[15]), 
            .I2(rand_setpoint[15]), .I3(n15573), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(n491), .I1(\FRAME_MATCHER.state [2]), .I2(n9460), 
            .I3(GND_net), .O(n17));   // coms.v(426[12] 547[6])
    defparam i1_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 blink_counter_2352_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n15608), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[21]), 
            .I3(n15548), .O(n144_adj_2472)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_23 (.CI(n15548), .I0(GND_net), .I1(rand_data[21]), 
            .CO(n15549));
    SB_CARRY rand_data_2350_add_4_10 (.CI(n15535), .I0(GND_net), .I1(rand_data[8]), 
            .CO(n15536));
    SB_CARRY blink_counter_2352_add_4_21 (.CI(n15608), .I0(GND_net), .I1(n7), 
            .CO(n15609));
    SB_LUT4 i15393_3_lut_4_lut (.I0(n29), .I1(\UART_TRANSMITTER.state [2]), 
            .I2(\UART_TRANSMITTER.state [0]), .I3(\UART_TRANSMITTER.state [1]), 
            .O(n17834));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hc888;
    SB_CARRY rand_setpoint_2351_add_4_17 (.CI(n15573), .I0(rand_data[15]), 
            .I1(rand_setpoint[15]), .CO(n15574));
    SB_LUT4 blink_counter_2352_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8), .I3(n15607), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8271_3_lut (.I0(n10425), .I1(r_Bit_Index_adj_2505[0]), .I2(n17260), 
            .I3(GND_net), .O(n10631));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8271_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i8337_3_lut_4_lut (.I0(\data_out[8] [1]), .I1(rand_setpoint[1]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10697));   // coms.v(280[12] 380[6])
    defparam i8337_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8333_3_lut_4_lut (.I0(\data_out[8] [4]), .I1(rand_setpoint[4]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10693));   // coms.v(280[12] 380[6])
    defparam i8333_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8332_3_lut_4_lut (.I0(\data_out[8] [5]), .I1(rand_setpoint[5]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10692));   // coms.v(280[12] 380[6])
    defparam i8332_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8331_3_lut_4_lut (.I0(\data_out[8] [6]), .I1(rand_setpoint[6]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10691));   // coms.v(280[12] 380[6])
    defparam i8331_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_4_lut_adj_775 (.I0(n7198), .I1(n9462), .I2(n17), .I3(n9435), 
            .O(n6));   // coms.v(426[12] 547[6])
    defparam i1_4_lut_adj_775.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_4_lut_adj_776 (.I0(n9453), .I1(n1651), .I2(n3977), .I3(n7198), 
            .O(n4));   // coms.v(426[12] 547[6])
    defparam i1_4_lut_adj_776.LUT_INIT = 16'h5450;
    SB_LUT4 i8330_3_lut_4_lut (.I0(\data_out[8] [7]), .I1(rand_setpoint[7]), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10690));   // coms.v(280[12] 380[6])
    defparam i8330_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8327_3_lut_4_lut (.I0(\data_out[9] [2]), .I1(data_out_9__2__N_367), 
            .I2(\UART_TRANSMITTER.state [2]), .I3(n2547), .O(n10687));   // coms.v(280[12] 380[6])
    defparam i8327_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_4_lut_adj_777 (.I0(n15837), .I1(r_SM_Main_adj_2509[1]), .I2(n10_adj_2412), 
            .I3(n12_adj_2410), .O(n16824));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_777.LUT_INIT = 16'h5150;
    SB_LUT4 i8004_3_lut_4_lut (.I0(\data_out[2] [2]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10364));   // coms.v(280[12] 380[6])
    defparam i8004_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i3_4_lut (.I0(n4), .I1(n17208), .I2(n1651), .I3(n6), .O(n8_adj_2459));   // coms.v(426[12] 547[6])
    defparam i3_4_lut.LUT_INIT = 16'hfbbb;
    SB_LUT4 i2_4_lut_4_lut (.I0(\UART_TRANSMITTER.state [1]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(n41), .I3(n9361), .O(n35));   // coms.v(280[12] 380[6])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_CARRY blink_counter_2352_add_4_20 (.CI(n15607), .I0(GND_net), .I1(n8), 
            .CO(n15608));
    SB_LUT4 i14716_2_lut_3_lut (.I0(\UART_TRANSMITTER.state [0]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n9361), .I3(GND_net), .O(n17154));
    defparam i14716_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i4_4_lut (.I0(\FRAME_MATCHER.state_31__N_1440 [1]), .I1(n8_adj_2459), 
            .I2(n3_adj_2408), .I3(n9452), .O(n18137));   // coms.v(426[12] 547[6])
    defparam i4_4_lut.LUT_INIT = 16'hfcfe;
    SB_LUT4 blink_counter_2352_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n15606), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_19 (.CI(n15606), .I0(GND_net), .I1(n9), 
            .CO(n15607));
    SB_LUT4 blink_counter_2352_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_2420), .I3(n15605), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[20]), 
            .I3(n15547), .O(n145_adj_2473)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(n12), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n9937), .O(n10_adj_2415));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i8007_3_lut_4_lut (.I0(\data_out[1] [6]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n4445), .O(n10367));   // coms.v(280[12] 380[6])
    defparam i8007_3_lut_4_lut.LUT_INIT = 16'haae2;
    SB_DFF blink_counter_2352__i25 (.Q(blink_counter[25]), .C(CLK_c), .D(n110));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i24 (.Q(blink_counter[24]), .C(CLK_c), .D(n111));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i23 (.Q(blink_counter[23]), .C(CLK_c), .D(n112));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i22 (.Q(blink_counter[22]), .C(CLK_c), .D(n113));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i21 (.Q(blink_counter[21]), .C(CLK_c), .D(n114));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i20 (.Q(n6_adj_2421), .C(CLK_c), .D(n115));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i19 (.Q(n7), .C(CLK_c), .D(n116));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i18 (.Q(n8), .C(CLK_c), .D(n117));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i17 (.Q(n9), .C(CLK_c), .D(n118));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i16 (.Q(n10_adj_2420), .C(CLK_c), .D(n119));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i15 (.Q(n11), .C(CLK_c), .D(n120));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i14 (.Q(n12_adj_2419), .C(CLK_c), .D(n121));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i8354_3_lut_4_lut (.I0(r_SM_Main_adj_2509[2]), .I1(r_SM_Main_2__N_2033_adj_2515[1]), 
            .I2(r_SM_Main_adj_2509[0]), .I3(r_SM_Main_adj_2509[1]), .O(n10714));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8354_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 i33_3_lut_adj_778 (.I0(n17631), .I1(r_Clock_Count[5]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16509));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_778.LUT_INIT = 16'hcaca;
    SB_LUT4 i8006_3_lut_4_lut (.I0(\data_out[1] [7]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10366));   // coms.v(280[12] 380[6])
    defparam i8006_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_CARRY blink_counter_2352_add_4_18 (.CI(n15605), .I0(GND_net), .I1(n10_adj_2420), 
            .CO(n15606));
    SB_LUT4 i33_3_lut_adj_779 (.I0(n17573), .I1(r_Clock_Count[4]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16567));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_779.LUT_INIT = 16'hcaca;
    SB_LUT4 i8002_3_lut_4_lut (.I0(\data_out[2] [5]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10362));   // coms.v(280[12] 380[6])
    defparam i8002_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 blink_counter_2352_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n15604), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8001_3_lut_4_lut (.I0(\data_out[2] [7]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10361));   // coms.v(280[12] 380[6])
    defparam i8001_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_DFF blink_counter_2352__i13 (.Q(n13), .C(CLK_c), .D(n122));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i12 (.Q(n14_adj_2424), .C(CLK_c), .D(n123));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i11 (.Q(n15), .C(CLK_c), .D(n124));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i10 (.Q(n16), .C(CLK_c), .D(n125));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i9 (.Q(n17_adj_2422), .C(CLK_c), .D(n126));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i8 (.Q(n18), .C(CLK_c), .D(n127_adj_2442));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i7 (.Q(n19), .C(CLK_c), .D(n128));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i6 (.Q(n20), .C(CLK_c), .D(n129));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i5 (.Q(n21), .C(CLK_c), .D(n130));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i4 (.Q(n22), .C(CLK_c), .D(n131));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i3 (.Q(n23), .C(CLK_c), .D(n132));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i2 (.Q(n24), .C(CLK_c), .D(n133));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_2352__i1 (.Q(n25), .C(CLK_c), .D(n134_adj_2429));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF rand_setpoint_2351__i31 (.Q(rand_setpoint[31]), .C(CLK_c), .D(n134));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i30 (.Q(rand_setpoint[30]), .C(CLK_c), .D(n135));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i29 (.Q(rand_setpoint[29]), .C(CLK_c), .D(n136));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 rand_setpoint_2351_add_4_16_lut (.I0(GND_net), .I1(rand_data[14]), 
            .I2(rand_setpoint[14]), .I3(n15572), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_17 (.CI(n15604), .I0(GND_net), .I1(n11), 
            .CO(n15605));
    SB_LUT4 rand_data_2350_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[7]), 
            .I3(n15534), .O(n158_adj_2486)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8000_3_lut_4_lut (.I0(\data_out[3] [0]), .I1(n2652), .I2(n4445), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n10360));   // coms.v(280[12] 380[6])
    defparam i8000_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 blink_counter_2352_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_2419), .I3(n15603), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7999_3_lut_4_lut (.I0(\data_out[3] [2]), .I1(n2652), .I2(n4445), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n10359));   // coms.v(280[12] 380[6])
    defparam i7999_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_DFF rand_setpoint_2351__i28 (.Q(rand_setpoint[28]), .C(CLK_c), .D(n137));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i27 (.Q(rand_setpoint[27]), .C(CLK_c), .D(n138));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i26 (.Q(rand_setpoint[26]), .C(CLK_c), .D(n139));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_CARRY rand_data_2350_add_4_9 (.CI(n15534), .I0(GND_net), .I1(rand_data[7]), 
            .CO(n15535));
    SB_DFF rand_setpoint_2351__i25 (.Q(rand_setpoint[25]), .C(CLK_c), .D(n140));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i24 (.Q(rand_setpoint[24]), .C(CLK_c), .D(n141));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i23 (.Q(rand_setpoint[23]), .C(CLK_c), .D(n142));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_CARRY blink_counter_2352_add_4_16 (.CI(n15603), .I0(GND_net), .I1(n12_adj_2419), 
            .CO(n15604));
    SB_LUT4 blink_counter_2352_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n15602), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2351__i22 (.Q(rand_setpoint[22]), .C(CLK_c), .D(n143));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i21 (.Q(rand_setpoint[21]), .C(CLK_c), .D(n144));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i20 (.Q(rand_setpoint[20]), .C(CLK_c), .D(n145));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i19 (.Q(rand_setpoint[19]), .C(CLK_c), .D(n146));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i18 (.Q(rand_setpoint[18]), .C(CLK_c), .D(n147));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i17 (.Q(rand_setpoint[17]), .C(CLK_c), .D(n148));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i16 (.Q(rand_setpoint[16]), .C(CLK_c), .D(n149));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i15 (.Q(rand_setpoint[15]), .C(CLK_c), .D(n150));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_CARRY rand_setpoint_2351_add_4_16 (.CI(n15572), .I0(rand_data[14]), 
            .I1(rand_setpoint[14]), .CO(n15573));
    SB_DFF rand_setpoint_2351__i14 (.Q(rand_setpoint[14]), .C(CLK_c), .D(n151));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i13 (.Q(rand_setpoint[13]), .C(CLK_c), .D(n152));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i12 (.Q(rand_setpoint[12]), .C(CLK_c), .D(n153));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i11 (.Q(rand_setpoint[11]), .C(CLK_c), .D(n154));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i10 (.Q(rand_setpoint[10]), .C(CLK_c), .D(n155));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i9 (.Q(rand_setpoint[9]), .C(CLK_c), .D(n156));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i8 (.Q(rand_setpoint[8]), .C(CLK_c), .D(n157));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i7 (.Q(rand_setpoint[7]), .C(CLK_c), .D(n158));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i6 (.Q(rand_setpoint[6]), .C(CLK_c), .D(n159));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 rand_setpoint_2351_add_4_15_lut (.I0(GND_net), .I1(rand_data[13]), 
            .I2(rand_setpoint[13]), .I3(n15571), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_setpoint_2351__i5 (.Q(rand_setpoint[5]), .C(CLK_c), .D(n160));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_LUT4 i7998_3_lut_4_lut (.I0(\data_out[3] [4]), .I1(n2652), .I2(n4445), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n10358));   // coms.v(280[12] 380[6])
    defparam i7998_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i33_3_lut_adj_780 (.I0(n17494), .I1(r_Clock_Count[3]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16649));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_780.LUT_INIT = 16'hcaca;
    SB_LUT4 i7997_3_lut_4_lut (.I0(\data_out[3] [5]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n4445), .O(n10357));   // coms.v(280[12] 380[6])
    defparam i7997_3_lut_4_lut.LUT_INIT = 16'haae2;
    SB_CARRY blink_counter_2352_add_4_15 (.CI(n15602), .I0(GND_net), .I1(n13), 
            .CO(n15603));
    SB_CARRY rand_setpoint_2351_add_4_15 (.CI(n15571), .I0(rand_data[13]), 
            .I1(rand_setpoint[13]), .CO(n15572));
    SB_LUT4 blink_counter_2352_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_2424), .I3(n15601), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_14 (.CI(n15601), .I0(GND_net), .I1(n14_adj_2424), 
            .CO(n15602));
    SB_LUT4 i33_3_lut_adj_781 (.I0(n17484), .I1(r_Clock_Count[2]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16651));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_781.LUT_INIT = 16'hcaca;
    SB_DFF rand_setpoint_2351__i4 (.Q(rand_setpoint[4]), .C(CLK_c), .D(n161));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i3 (.Q(rand_setpoint[3]), .C(CLK_c), .D(n162));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i2 (.Q(rand_setpoint[2]), .C(CLK_c), .D(n163));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_setpoint_2351__i1 (.Q(rand_setpoint[1]), .C(CLK_c), .D(n164));   // verilog/TinyFPGA_B.v(81[21:44])
    SB_DFF rand_data_2350__i31 (.Q(rand_data[31]), .C(CLK_c), .D(n134_adj_2462));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i30 (.Q(rand_data[30]), .C(CLK_c), .D(n135_adj_2463));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i29 (.Q(rand_data[29]), .C(CLK_c), .D(n136_adj_2464));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i28 (.Q(rand_data[28]), .C(CLK_c), .D(n137_adj_2465));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i27 (.Q(rand_data[27]), .C(CLK_c), .D(n138_adj_2466));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i26 (.Q(rand_data[26]), .C(CLK_c), .D(n139_adj_2467));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i25 (.Q(rand_data[25]), .C(CLK_c), .D(n140_adj_2468));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i24 (.Q(rand_data[24]), .C(CLK_c), .D(n141_adj_2469));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 blink_counter_2352_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n15600), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2350__i23 (.Q(rand_data[23]), .C(CLK_c), .D(n142_adj_2470));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i11_4_lut (.I0(rand_setpoint[16]), .I1(\data_out[6] [0]), .I2(n10055), 
            .I3(n2547), .O(n16607));   // coms.v(280[12] 380[6])
    defparam i11_4_lut.LUT_INIT = 16'hac0c;
    SB_CARRY blink_counter_2352_add_4_13 (.CI(n15600), .I0(GND_net), .I1(n15), 
            .CO(n15601));
    SB_LUT4 i8298_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10658));   // coms.v(426[12] 547[6])
    defparam i8298_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2350__i22 (.Q(rand_data[22]), .C(CLK_c), .D(n143_adj_2471));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 i8299_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10659));   // coms.v(426[12] 547[6])
    defparam i8299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8300_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10660));   // coms.v(426[12] 547[6])
    defparam i8300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8259_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n16897), 
            .I3(GND_net), .O(n10619));   // coms.v(426[12] 547[6])
    defparam i8259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8301_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10661));   // coms.v(426[12] 547[6])
    defparam i8301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8302_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10662));   // coms.v(426[12] 547[6])
    defparam i8302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8303_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10663));   // coms.v(426[12] 547[6])
    defparam i8303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8260_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n16897), 
            .I3(GND_net), .O(n10620));   // coms.v(426[12] 547[6])
    defparam i8260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rand_setpoint_2351_add_4_14_lut (.I0(GND_net), .I1(rand_data[12]), 
            .I2(rand_setpoint[12]), .I3(n15570), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2352_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n15599), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_12 (.CI(n15599), .I0(GND_net), .I1(n16), 
            .CO(n15600));
    SB_CARRY rand_setpoint_2351_add_4_14 (.CI(n15570), .I0(rand_data[12]), 
            .I1(rand_setpoint[12]), .CO(n15571));
    SB_CARRY rand_data_2350_add_4_22 (.CI(n15547), .I0(GND_net), .I1(rand_data[20]), 
            .CO(n15548));
    SB_LUT4 blink_counter_2352_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_2422), .I3(n15598), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_13_lut (.I0(GND_net), .I1(rand_data[11]), 
            .I2(rand_setpoint[11]), .I3(n15569), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_11 (.CI(n15598), .I0(GND_net), .I1(n17_adj_2422), 
            .CO(n15599));
    SB_DFF rand_data_2350__i21 (.Q(rand_data[21]), .C(CLK_c), .D(n144_adj_2472));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i20 (.Q(rand_data[20]), .C(CLK_c), .D(n145_adj_2473));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i19 (.Q(rand_data[19]), .C(CLK_c), .D(n146_adj_2474));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i18 (.Q(rand_data[18]), .C(CLK_c), .D(n147_adj_2475));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY rand_setpoint_2351_add_4_13 (.CI(n15569), .I0(rand_data[11]), 
            .I1(rand_setpoint[11]), .CO(n15570));
    SB_DFF rand_data_2350__i17 (.Q(rand_data[17]), .C(CLK_c), .D(n148_adj_2476));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i16 (.Q(rand_data[16]), .C(CLK_c), .D(n149_adj_2477));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i15 (.Q(rand_data[15]), .C(CLK_c), .D(n150_adj_2478));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i14 (.Q(rand_data[14]), .C(CLK_c), .D(n151_adj_2479));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i13 (.Q(rand_data[13]), .C(CLK_c), .D(n152_adj_2480));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i12 (.Q(rand_data[12]), .C(CLK_c), .D(n153_adj_2481));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i11 (.Q(rand_data[11]), .C(CLK_c), .D(n154_adj_2482));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 rand_data_2350_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[6]), 
            .I3(n15533), .O(n159_adj_2487)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2350__i10 (.Q(rand_data[10]), .C(CLK_c), .D(n155_adj_2483));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 rand_data_2350_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[19]), 
            .I3(n15546), .O(n146_adj_2474)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2350__i9 (.Q(rand_data[9]), .C(CLK_c), .D(n156_adj_2484));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY rand_data_2350_add_4_21 (.CI(n15546), .I0(GND_net), .I1(rand_data[19]), 
            .CO(n15547));
    SB_LUT4 blink_counter_2352_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n15597), .O(n127_adj_2442)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF rand_data_2350__i8 (.Q(rand_data[8]), .C(CLK_c), .D(n157_adj_2485));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i7 (.Q(rand_data[7]), .C(CLK_c), .D(n158_adj_2486));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i6 (.Q(rand_data[6]), .C(CLK_c), .D(n159_adj_2487));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i5 (.Q(rand_data[5]), .C(CLK_c), .D(n160_adj_2488));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i4 (.Q(rand_data[4]), .C(CLK_c), .D(n161_adj_2489));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i3 (.Q(rand_data[3]), .C(CLK_c), .D(n162_adj_2490));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i2 (.Q(rand_data[2]), .C(CLK_c), .D(n163_adj_2491));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_DFF rand_data_2350__i1 (.Q(rand_data[1]), .C(CLK_c), .D(n164_adj_2492));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_CARRY rand_data_2350_add_4_8 (.CI(n15533), .I0(GND_net), .I1(rand_data[6]), 
            .CO(n15534));
    SB_LUT4 i8261_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n16897), 
            .I3(GND_net), .O(n10621));   // coms.v(426[12] 547[6])
    defparam i8261_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY blink_counter_2352_add_4_10 (.CI(n15597), .I0(GND_net), .I1(n18), 
            .CO(n15598));
    SB_LUT4 blink_counter_2352_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n15596), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_12_lut (.I0(GND_net), .I1(rand_data[10]), 
            .I2(rand_setpoint[10]), .I3(n15568), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_12 (.CI(n15568), .I0(rand_data[10]), 
            .I1(rand_setpoint[10]), .CO(n15569));
    SB_LUT4 i8262_3_lut (.I0(\data_in_frame[0] [4]), .I1(rx_data[4]), .I2(n16897), 
            .I3(GND_net), .O(n10622));   // coms.v(426[12] 547[6])
    defparam i8262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rand_setpoint_2351_add_4_11_lut (.I0(GND_net), .I1(rand_data[9]), 
            .I2(rand_setpoint[9]), .I3(n15567), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_9 (.CI(n15596), .I0(GND_net), .I1(n19), 
            .CO(n15597));
    SB_LUT4 rand_data_2350_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[18]), 
            .I3(n15545), .O(n147_adj_2475)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15444_4_lut (.I0(r_SM_Main_adj_2506[2]), .I1(n17601), .I2(n17602), 
            .I3(r_SM_Main_adj_2506[1]), .O(n13510));
    defparam i15444_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i25_3_lut (.I0(r_Clock_Count_adj_2510[6]), .I1(n17634), .I2(r_SM_Main_adj_2509[2]), 
            .I3(GND_net), .O(n16483));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rand_setpoint_2351_add_4_11 (.CI(n15567), .I0(rand_data[9]), 
            .I1(rand_setpoint[9]), .CO(n15568));
    SB_LUT4 i8304_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10664));   // coms.v(426[12] 547[6])
    defparam i8304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8263_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n16897), 
            .I3(GND_net), .O(n10623));   // coms.v(426[12] 547[6])
    defparam i8263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8264_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n16897), 
            .I3(GND_net), .O(n10624));   // coms.v(426[12] 547[6])
    defparam i8264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7995_3_lut_4_lut (.I0(\data_out[3] [7]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n4445), .O(n10355));   // coms.v(280[12] 380[6])
    defparam i7995_3_lut_4_lut.LUT_INIT = 16'haae2;
    SB_LUT4 rand_setpoint_2351_add_4_10_lut (.I0(GND_net), .I1(rand_data[8]), 
            .I2(rand_setpoint[8]), .I3(n15566), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8305_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10665));   // coms.v(426[12] 547[6])
    defparam i8305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2352_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n15595), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8306_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10666));   // coms.v(426[12] 547[6])
    defparam i8306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33_3_lut_adj_782 (.I0(n17461), .I1(r_Clock_Count[1]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16671));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i33_3_lut_adj_782.LUT_INIT = 16'hcaca;
    SB_LUT4 i8307_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10667));   // coms.v(426[12] 547[6])
    defparam i8307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8308_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10668));   // coms.v(426[12] 547[6])
    defparam i8308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8265_3_lut (.I0(\data_in_frame[0] [1]), .I1(rx_data[1]), .I2(n16897), 
            .I3(GND_net), .O(n10625));   // coms.v(426[12] 547[6])
    defparam i8265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8429_3_lut (.I0(\data_out_frame2[13] [0]), .I1(rand_data[24]), 
            .I2(n10197), .I3(GND_net), .O(n10789));   // coms.v(426[12] 547[6])
    defparam i8429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8430_3_lut (.I0(\data_out_frame2[13] [1]), .I1(rand_data[25]), 
            .I2(n10197), .I3(GND_net), .O(n10790));   // coms.v(426[12] 547[6])
    defparam i8430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8431_3_lut (.I0(\data_out_frame2[13] [2]), .I1(rand_data[26]), 
            .I2(n10197), .I3(GND_net), .O(n10791));   // coms.v(426[12] 547[6])
    defparam i8431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31_3_lut_adj_783 (.I0(r_Clock_Count_adj_2510[5]), .I1(n17629), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16517));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut_adj_783.LUT_INIT = 16'hacac;
    SB_LUT4 i8432_3_lut (.I0(\data_out_frame2[13] [3]), .I1(rand_data[27]), 
            .I2(n10197), .I3(GND_net), .O(n10792));   // coms.v(426[12] 547[6])
    defparam i8432_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_2352_add_4_8 (.CI(n15595), .I0(GND_net), .I1(n20), 
            .CO(n15596));
    SB_CARRY rand_data_2350_add_4_20 (.CI(n15545), .I0(GND_net), .I1(rand_data[18]), 
            .CO(n15546));
    SB_CARRY rand_setpoint_2351_add_4_10 (.CI(n15566), .I0(rand_data[8]), 
            .I1(rand_setpoint[8]), .CO(n15567));
    SB_LUT4 i31_3_lut_adj_784 (.I0(r_Clock_Count_adj_2510[4]), .I1(n17567), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16577));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut_adj_784.LUT_INIT = 16'hacac;
    SB_LUT4 i8309_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10669));   // coms.v(426[12] 547[6])
    defparam i8309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8405_3_lut (.I0(\data_out_frame2[10] [0]), .I1(rand_data[16]), 
            .I2(n10197), .I3(GND_net), .O(n10765));   // coms.v(426[12] 547[6])
    defparam i8405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8406_3_lut (.I0(\data_out_frame2[10] [1]), .I1(rand_data[17]), 
            .I2(n10197), .I3(GND_net), .O(n10766));   // coms.v(426[12] 547[6])
    defparam i8406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2352_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n15594), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14706_3_lut (.I0(n12), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17144));
    defparam i14706_3_lut.LUT_INIT = 16'hd5d5;
    SB_LUT4 i14845_4_lut (.I0(n15701), .I1(n9937), .I2(n17144), .I3(n9406), 
            .O(n16828));
    defparam i14845_4_lut.LUT_INIT = 16'h1505;
    SB_LUT4 i8310_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10670));   // coms.v(426[12] 547[6])
    defparam i8310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_785 (.I0(n16855), .I1(r_Clock_Count_adj_2504[7]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16469));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_785.LUT_INIT = 16'heaea;
    SB_LUT4 rand_data_2350_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[5]), 
            .I3(n15532), .O(n160_adj_2488)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_7 (.CI(n15594), .I0(GND_net), .I1(n21), 
            .CO(n15595));
    SB_LUT4 blink_counter_2352_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22), .I3(n15593), .O(n131)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_786 (.I0(n16856), .I1(r_Clock_Count_adj_2504[6]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16479));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_786.LUT_INIT = 16'heaea;
    SB_LUT4 i1_3_lut_adj_787 (.I0(n16857), .I1(r_Clock_Count_adj_2504[5]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16515));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_787.LUT_INIT = 16'heaea;
    SB_CARRY blink_counter_2352_add_4_6 (.CI(n15593), .I0(GND_net), .I1(n22), 
            .CO(n15594));
    SB_LUT4 blink_counter_2352_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23), .I3(n15592), .O(n132)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_788 (.I0(n16854), .I1(r_Clock_Count_adj_2504[4]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16569));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_788.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_789 (.I0(n15701), .I1(n13276), .I2(n10_adj_2415), 
            .I3(n12), .O(n16844));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_789.LUT_INIT = 16'h5150;
    SB_LUT4 rand_setpoint_2351_add_4_9_lut (.I0(GND_net), .I1(rand_data[7]), 
            .I2(rand_setpoint[7]), .I3(n15565), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_7 (.CI(n15532), .I0(GND_net), .I1(rand_data[5]), 
            .CO(n15533));
    SB_CARRY blink_counter_2352_add_4_5 (.CI(n15592), .I0(GND_net), .I1(n23), 
            .CO(n15593));
    SB_LUT4 i8275_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_2409), 
            .I3(n9477), .O(n10635));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i8275_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3_1_lut (.I0(n29), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53));   // coms.v(280[12] 380[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rand_setpoint_2351_add_4_9 (.CI(n15565), .I0(rand_data[7]), 
            .I1(rand_setpoint[7]), .CO(n15566));
    SB_LUT4 i14861_4_lut (.I0(blink_counter[22]), .I1(blink_counter[23]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17299));
    defparam i14861_4_lut.LUT_INIT = 16'hfec4;
    SB_LUT4 rand_data_2350_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[17]), 
            .I3(n15544), .O(n148_adj_2476)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14860_4_lut (.I0(blink_counter[23]), .I1(blink_counter[22]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n17298));
    defparam i14860_4_lut.LUT_INIT = 16'hcf08;
    SB_LUT4 i14862_3_lut (.I0(n17298), .I1(n17299), .I2(blink_counter[25]), 
            .I3(GND_net), .O(LED_c));
    defparam i14862_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 blink_counter_2352_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n15591), .O(n133)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_19 (.CI(n15544), .I0(GND_net), .I1(rand_data[17]), 
            .CO(n15545));
    SB_LUT4 i8407_3_lut (.I0(\data_out_frame2[10] [2]), .I1(rand_data[18]), 
            .I2(n10197), .I3(GND_net), .O(n10767));   // coms.v(426[12] 547[6])
    defparam i8407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8311_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10671));   // coms.v(426[12] 547[6])
    defparam i8311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8312_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10672));   // coms.v(426[12] 547[6])
    defparam i8312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8408_3_lut (.I0(\data_out_frame2[10] [3]), .I1(rand_data[19]), 
            .I2(n10197), .I3(GND_net), .O(n10768));   // coms.v(426[12] 547[6])
    defparam i8408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8465_3_lut (.I0(\data_out_frame2[17] [4]), .I1(rand_data[12]), 
            .I2(n10197), .I3(GND_net), .O(n10825));   // coms.v(426[12] 547[6])
    defparam i8465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_790 (.I0(n16858), .I1(r_Clock_Count_adj_2504[3]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16571));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_790.LUT_INIT = 16'heaea;
    SB_LUT4 i8313_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10673));   // coms.v(426[12] 547[6])
    defparam i8313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[16]), 
            .I3(n15543), .O(n149_adj_2477)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_8_lut (.I0(GND_net), .I1(rand_data[6]), 
            .I2(rand_setpoint[6]), .I3(n15564), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[4]), 
            .I3(n15531), .O(n161_adj_2489)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8466_3_lut (.I0(\data_out_frame2[17] [5]), .I1(rand_data[13]), 
            .I2(n10197), .I3(GND_net), .O(n10826));   // coms.v(426[12] 547[6])
    defparam i8466_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2350_add_4_6 (.CI(n15531), .I0(GND_net), .I1(rand_data[4]), 
            .CO(n15532));
    SB_CARRY blink_counter_2352_add_4_4 (.CI(n15591), .I0(GND_net), .I1(n24), 
            .CO(n15592));
    SB_LUT4 i1_3_lut_adj_791 (.I0(n16860), .I1(r_Clock_Count_adj_2504[2]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16573));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_791.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_792 (.I0(n29), .I1(n10031), .I2(n17230), .I3(n9358), 
            .O(n41));   // coms.v(280[12] 380[6])
    defparam i1_4_lut_adj_792.LUT_INIT = 16'hcecc;
    SB_LUT4 i8314_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10674));   // coms.v(426[12] 547[6])
    defparam i8314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8315_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10675));   // coms.v(426[12] 547[6])
    defparam i8315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_793 (.I0(r_SM_Main_adj_2506[2]), .I1(r_SM_Main_adj_2506[1]), 
            .I2(n6_adj_2461), .I3(r_SM_Main_adj_2506[0]), .O(n17_adj_2416));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_793.LUT_INIT = 16'hbaaa;
    SB_LUT4 i8467_3_lut (.I0(\data_out_frame2[17] [6]), .I1(rand_data[14]), 
            .I2(n10197), .I3(GND_net), .O(n10827));   // coms.v(426[12] 547[6])
    defparam i8467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15262_4_lut (.I0(n10031), .I1(n9357), .I2(n29), .I3(n445), 
            .O(n17479));   // coms.v(280[12] 380[6])
    defparam i15262_4_lut.LUT_INIT = 16'h5515;
    SB_LUT4 i8316_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10676));   // coms.v(426[12] 547[6])
    defparam i8316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_794 (.I0(n16853), .I1(r_Clock_Count_adj_2504[1]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16575));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_794.LUT_INIT = 16'heaea;
    SB_LUT4 i57_4_lut (.I0(n16886), .I1(n17479), .I2(\UART_TRANSMITTER.state [1]), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n38));   // coms.v(280[12] 380[6])
    defparam i57_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i8039_4_lut (.I0(n10398), .I1(r_Bit_Index_adj_2511[1]), .I2(r_Bit_Index_adj_2511[0]), 
            .I3(n17194), .O(n10399));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8039_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i8036_4_lut (.I0(n10398), .I1(r_Bit_Index_adj_2511[2]), .I2(n5029), 
            .I3(n17194), .O(n10396));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8036_4_lut.LUT_INIT = 16'h8828;
    SB_LUT4 i15433_4_lut (.I0(\UART_TRANSMITTER.state [2]), .I1(n38), .I2(n35), 
            .I3(n17154), .O(n33));   // coms.v(280[12] 380[6])
    defparam i15433_4_lut.LUT_INIT = 16'haf23;
    SB_LUT4 i8317_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10677));   // coms.v(426[12] 547[6])
    defparam i8317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8318_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10678));   // coms.v(426[12] 547[6])
    defparam i8318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_2352_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(n15590), .O(n134_adj_2429)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25_3_lut_adj_795 (.I0(r_Clock_Count_adj_2510[7]), .I1(n17640), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16473));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_795.LUT_INIT = 16'hacac;
    SB_LUT4 i8319_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10679));   // coms.v(426[12] 547[6])
    defparam i8319_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_8 (.CI(n15564), .I0(rand_data[6]), 
            .I1(rand_setpoint[6]), .CO(n15565));
    SB_CARRY rand_data_2350_add_4_18 (.CI(n15543), .I0(GND_net), .I1(rand_data[16]), 
            .CO(n15544));
    SB_LUT4 i1_4_lut_adj_796 (.I0(r_SM_Main_adj_2506[0]), .I1(n17222), .I2(r_Clock_Count_adj_2504[5]), 
            .I3(n16863), .O(n16810));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_796.LUT_INIT = 16'ha8aa;
    SB_LUT4 i1_3_lut_4_lut_adj_797 (.I0(n12_adj_2410), .I1(r_SM_Main_adj_2509[1]), 
            .I2(r_SM_Main_adj_2509[2]), .I3(n9929), .O(n10_adj_2412));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut_adj_797.LUT_INIT = 16'h080c;
    SB_LUT4 i2_4_lut (.I0(n16867), .I1(n17_adj_2416), .I2(r_SM_Main_adj_2506[1]), 
            .I3(n16810), .O(n16852));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_4_lut.LUT_INIT = 16'h2322;
    SB_LUT4 i1_3_lut_4_lut_adj_798 (.I0(n16795), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n127), .I3(n7198), .O(n3_adj_2408));   // coms.v(426[12] 547[6])
    defparam i1_3_lut_4_lut_adj_798.LUT_INIT = 16'h4500;
    SB_LUT4 i8320_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10680));   // coms.v(426[12] 547[6])
    defparam i8320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8321_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10681));   // coms.v(426[12] 547[6])
    defparam i8321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8322_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10682));   // coms.v(426[12] 547[6])
    defparam i8322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8323_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10683));   // coms.v(426[12] 547[6])
    defparam i8323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8324_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10684));   // coms.v(426[12] 547[6])
    defparam i8324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8409_3_lut (.I0(\data_out_frame2[10] [4]), .I1(rand_data[20]), 
            .I2(n10197), .I3(GND_net), .O(n10769));   // coms.v(426[12] 547[6])
    defparam i8409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31_3_lut_adj_799 (.I0(r_Clock_Count_adj_2510[3]), .I1(n17457), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16673));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut_adj_799.LUT_INIT = 16'hacac;
    SB_LUT4 rand_setpoint_2351_add_4_7_lut (.I0(GND_net), .I1(rand_data[5]), 
            .I2(rand_setpoint[5]), .I3(n15563), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_7 (.CI(n15563), .I0(rand_data[5]), 
            .I1(rand_setpoint[5]), .CO(n15564));
    SB_LUT4 i8325_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10685));   // coms.v(426[12] 547[6])
    defparam i8325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_6_lut (.I0(GND_net), .I1(rand_data[4]), 
            .I2(rand_setpoint[4]), .I3(n15562), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_2352_add_4_3 (.CI(n15590), .I0(GND_net), .I1(n25), 
            .CO(n15591));
    SB_LUT4 i8326_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10686));   // coms.v(426[12] 547[6])
    defparam i8326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[3]), 
            .I3(n15530), .O(n162_adj_2490)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[15]), 
            .I3(n15542), .O(n150_adj_2478)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_6 (.CI(n15562), .I0(rand_data[4]), 
            .I1(rand_setpoint[4]), .CO(n15563));
    SB_CARRY rand_data_2350_add_4_17 (.CI(n15542), .I0(GND_net), .I1(rand_data[15]), 
            .CO(n15543));
    SB_CARRY rand_data_2350_add_4_5 (.CI(n15530), .I0(GND_net), .I1(rand_data[3]), 
            .CO(n15531));
    SB_LUT4 rand_data_2350_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[14]), 
            .I3(n15541), .O(n151_adj_2479)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_5_lut (.I0(GND_net), .I1(rand_data[3]), 
            .I2(rand_setpoint[3]), .I3(n15561), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_2352_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26), .I3(VCC_net), .O(n135_adj_2428)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_2352_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_5 (.CI(n15561), .I0(rand_data[3]), 
            .I1(rand_setpoint[3]), .CO(n15562));
    SB_LUT4 i1_3_lut_adj_800 (.I0(n16859), .I1(r_Clock_Count_adj_2504[0]), 
            .I2(n17_adj_2416), .I3(GND_net), .O(n16547));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_800.LUT_INIT = 16'heaea;
    SB_CARRY blink_counter_2352_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n26), 
            .CO(n15590));
    SB_LUT4 rand_setpoint_2351_add_4_4_lut (.I0(GND_net), .I1(rand_data[2]), 
            .I2(rand_setpoint[2]), .I3(n15560), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_16 (.CI(n15541), .I0(GND_net), .I1(rand_data[14]), 
            .CO(n15542));
    SB_LUT4 rand_data_2350_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[2]), 
            .I3(n15529), .O(n163_adj_2491)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_33_lut (.I0(GND_net), .I1(rand_data[31]), 
            .I2(rand_setpoint[31]), .I3(n15589), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_4 (.CI(n15560), .I0(rand_data[2]), 
            .I1(rand_setpoint[2]), .CO(n15561));
    SB_LUT4 rand_setpoint_2351_add_4_32_lut (.I0(GND_net), .I1(rand_data[30]), 
            .I2(rand_setpoint[30]), .I3(n15588), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_3_lut (.I0(GND_net), .I1(rand_data[1]), 
            .I2(rand_setpoint[1]), .I3(n15559), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8410_3_lut (.I0(\data_out_frame2[10] [5]), .I1(rand_data[21]), 
            .I2(n10197), .I3(GND_net), .O(n10770));   // coms.v(426[12] 547[6])
    defparam i8410_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_3 (.CI(n15559), .I0(rand_data[1]), 
            .I1(rand_setpoint[1]), .CO(n15560));
    SB_LUT4 i8411_3_lut (.I0(\data_out_frame2[10] [6]), .I1(rand_data[22]), 
            .I2(n10197), .I3(GND_net), .O(n10771));   // coms.v(426[12] 547[6])
    defparam i8411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_2_lut (.I0(GND_net), .I1(rand_data[0]), 
            .I2(rand_setpoint[0]), .I3(GND_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8412_3_lut (.I0(\data_out_frame2[10] [7]), .I1(rand_data[23]), 
            .I2(n10197), .I3(GND_net), .O(n10772));   // coms.v(426[12] 547[6])
    defparam i8412_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_2 (.CI(GND_net), .I0(rand_data[0]), 
            .I1(rand_setpoint[0]), .CO(n15559));
    SB_CARRY rand_setpoint_2351_add_4_32 (.CI(n15588), .I0(rand_data[30]), 
            .I1(rand_setpoint[30]), .CO(n15589));
    SB_LUT4 rand_setpoint_2351_add_4_31_lut (.I0(GND_net), .I1(rand_data[29]), 
            .I2(rand_setpoint[29]), .I3(n15587), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_31 (.CI(n15587), .I0(rand_data[29]), 
            .I1(rand_setpoint[29]), .CO(n15588));
    SB_LUT4 rand_data_2350_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[13]), 
            .I3(n15540), .O(n152_adj_2480)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_15 (.CI(n15540), .I0(GND_net), .I1(rand_data[13]), 
            .CO(n15541));
    SB_LUT4 rand_setpoint_2351_add_4_30_lut (.I0(GND_net), .I1(rand_data[28]), 
            .I2(rand_setpoint[28]), .I3(n15586), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8328_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10688));   // coms.v(426[12] 547[6])
    defparam i8328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[12]), 
            .I3(n15539), .O(n153_adj_2481)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8468_3_lut (.I0(\data_out_frame2[17] [7]), .I1(rand_data[15]), 
            .I2(n10197), .I3(GND_net), .O(n10828));   // coms.v(426[12] 547[6])
    defparam i8468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8329_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10689));   // coms.v(426[12] 547[6])
    defparam i8329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8012_3_lut_4_lut (.I0(\data_out[0] [3]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10372));   // coms.v(280[12] 380[6])
    defparam i8012_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_CARRY rand_setpoint_2351_add_4_30 (.CI(n15586), .I0(rand_data[28]), 
            .I1(rand_setpoint[28]), .CO(n15587));
    SB_CARRY rand_data_2350_add_4_14 (.CI(n15539), .I0(GND_net), .I1(rand_data[12]), 
            .CO(n15540));
    SB_CARRY rand_data_2350_add_4_4 (.CI(n15529), .I0(GND_net), .I1(rand_data[2]), 
            .CO(n15530));
    SB_LUT4 i8469_3_lut (.I0(\data_out_frame2[18] [0]), .I1(rand_data[0]), 
            .I2(n10197), .I3(GND_net), .O(n10829));   // coms.v(426[12] 547[6])
    defparam i8469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8011_3_lut_4_lut (.I0(\data_out[0] [5]), .I1(n2652), .I2(n4445), 
            .I3(\UART_TRANSMITTER.state [0]), .O(n10371));   // coms.v(280[12] 380[6])
    defparam i8011_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8470_3_lut (.I0(\data_out_frame2[18] [1]), .I1(rand_data[1]), 
            .I2(n10197), .I3(GND_net), .O(n10830));   // coms.v(426[12] 547[6])
    defparam i8470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8471_3_lut (.I0(\data_out_frame2[18] [2]), .I1(rand_data[2]), 
            .I2(n10197), .I3(GND_net), .O(n10831));   // coms.v(426[12] 547[6])
    defparam i8471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8457_3_lut (.I0(\data_out_frame2[16] [4]), .I1(rand_data[4]), 
            .I2(n10197), .I3(GND_net), .O(n10817));   // coms.v(426[12] 547[6])
    defparam i8457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8458_3_lut (.I0(\data_out_frame2[16] [5]), .I1(rand_data[5]), 
            .I2(n10197), .I3(GND_net), .O(n10818));   // coms.v(426[12] 547[6])
    defparam i8458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8459_3_lut (.I0(\data_out_frame2[16] [6]), .I1(rand_data[6]), 
            .I2(n10197), .I3(GND_net), .O(n10819));   // coms.v(426[12] 547[6])
    defparam i8459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8460_3_lut (.I0(\data_out_frame2[16] [7]), .I1(rand_data[7]), 
            .I2(n10197), .I3(GND_net), .O(n10820));   // coms.v(426[12] 547[6])
    defparam i8460_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rand_data_2350__i0 (.Q(rand_data[0]), .C(CLK_c), .D(n165_adj_2493));   // verilog/TinyFPGA_B.v(80[20:33])
    SB_LUT4 rand_setpoint_2351_add_4_29_lut (.I0(GND_net), .I1(rand_data[27]), 
            .I2(rand_setpoint[27]), .I3(n15585), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8461_3_lut (.I0(\data_out_frame2[17] [0]), .I1(rand_data[8]), 
            .I2(n10197), .I3(GND_net), .O(n10821));   // coms.v(426[12] 547[6])
    defparam i8461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[31]), 
            .I3(n15558), .O(n134_adj_2462)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_29 (.CI(n15585), .I0(rand_data[27]), 
            .I1(rand_setpoint[27]), .CO(n15586));
    SB_LUT4 i8335_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n10695));   // coms.v(426[12] 547[6])
    defparam i8335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8462_3_lut (.I0(\data_out_frame2[17] [1]), .I1(rand_data[9]), 
            .I2(n10197), .I3(GND_net), .O(n10822));   // coms.v(426[12] 547[6])
    defparam i8462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[1]), 
            .I3(n15528), .O(n164_adj_2492)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_setpoint_2351_add_4_28_lut (.I0(GND_net), .I1(rand_data[26]), 
            .I2(rand_setpoint[26]), .I3(n15584), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_3 (.CI(n15528), .I0(GND_net), .I1(rand_data[1]), 
            .CO(n15529));
    SB_LUT4 rand_data_2350_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[0]), 
            .I3(VCC_net), .O(n165_adj_2493)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[30]), 
            .I3(n15557), .O(n135_adj_2463)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(rand_data[0]), 
            .CO(n15528));
    SB_CARRY rand_setpoint_2351_add_4_28 (.CI(n15584), .I0(rand_data[26]), 
            .I1(rand_setpoint[26]), .CO(n15585));
    SB_LUT4 rand_setpoint_2351_add_4_27_lut (.I0(GND_net), .I1(rand_data[25]), 
            .I2(rand_setpoint[25]), .I3(n15583), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_32 (.CI(n15557), .I0(GND_net), .I1(rand_data[30]), 
            .CO(n15558));
    SB_LUT4 i8413_3_lut (.I0(\data_out_frame2[11] [0]), .I1(rand_data[8]), 
            .I2(n10197), .I3(GND_net), .O(n10773));   // coms.v(426[12] 547[6])
    defparam i8413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut (.I0(n10141), .I1(\UART_TRANSMITTER.state [1]), .I2(\UART_TRANSMITTER.state [0]), 
            .I3(GND_net), .O(n16255));   // coms.v(280[12] 380[6])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 rand_data_2350_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[11]), 
            .I3(n15538), .O(n154_adj_2482)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25_3_lut_adj_801 (.I0(r_Clock_Count_adj_2510[8]), .I1(n17458), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16463));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_801.LUT_INIT = 16'hacac;
    GND i1 (.Y(GND_net));
    SB_LUT4 i8433_3_lut (.I0(\data_out_frame2[13] [4]), .I1(rand_data[28]), 
            .I2(n10197), .I3(GND_net), .O(n10793));   // coms.v(426[12] 547[6])
    defparam i8433_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_data_2350_add_4_13 (.CI(n15538), .I0(GND_net), .I1(rand_data[11]), 
            .CO(n15539));
    SB_LUT4 i8013_3_lut_4_lut (.I0(\data_out[0] [1]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10373));   // coms.v(280[12] 380[6])
    defparam i8013_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i8338_3_lut (.I0(\data_out[8] [0]), .I1(rand_setpoint[0]), .I2(data_out_10__7__N_110), 
            .I3(GND_net), .O(n10698));   // coms.v(280[12] 380[6])
    defparam i8338_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_27 (.CI(n15583), .I0(rand_data[25]), 
            .I1(rand_setpoint[25]), .CO(n15584));
    SB_LUT4 i8414_3_lut (.I0(\data_out_frame2[11] [1]), .I1(rand_data[9]), 
            .I2(n10197), .I3(GND_net), .O(n10774));   // coms.v(426[12] 547[6])
    defparam i8414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8365_3_lut (.I0(\data_out_frame2[5] [0]), .I1(rand_data[24]), 
            .I2(n10197), .I3(GND_net), .O(n10725));   // coms.v(426[12] 547[6])
    defparam i8365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_data_2350_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[29]), 
            .I3(n15556), .O(n136_adj_2464)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_31 (.CI(n15556), .I0(GND_net), .I1(rand_data[29]), 
            .CO(n15557));
    SB_LUT4 i2_2_lut_4_lut (.I0(r_SM_Main_adj_2509[1]), .I1(r_SM_Main_adj_2509[2]), 
            .I2(r_SM_Main_2__N_2033_adj_2515[1]), .I3(r_SM_Main_adj_2509[0]), 
            .O(n15689));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i8366_3_lut (.I0(\data_out_frame2[5] [1]), .I1(rand_data[25]), 
            .I2(n10197), .I3(GND_net), .O(n10726));   // coms.v(426[12] 547[6])
    defparam i8366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_26_lut (.I0(GND_net), .I1(rand_data[24]), 
            .I2(rand_setpoint[24]), .I3(n15582), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[10]), 
            .I3(n15537), .O(n155_adj_2483)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[28]), 
            .I3(n15555), .O(n137_adj_2465)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(\UART_TRANSMITTER.state [2]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(GND_net), .O(n4445));   // coms.v(280[12] 380[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_802 (.I0(n9462), .I1(n9453), .I2(n16775), 
            .I3(n3977), .O(n16776));   // coms.v(426[12] 547[6])
    defparam i1_3_lut_4_lut_adj_802.LUT_INIT = 16'hf0f7;
    SB_LUT4 i8247_3_lut (.I0(n10398), .I1(r_Bit_Index_adj_2511[0]), .I2(n17194), 
            .I3(GND_net), .O(n10607));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8247_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i8014_3_lut_4_lut (.I0(\data_out[0] [0]), .I1(\UART_TRANSMITTER.state [0]), 
            .I2(\UART_TRANSMITTER.state [1]), .I3(n4445), .O(n10374));   // coms.v(280[12] 380[6])
    defparam i8014_3_lut_4_lut.LUT_INIT = 16'haae2;
    SB_LUT4 i8005_3_lut_4_lut (.I0(\data_out[2] [0]), .I1(\UART_TRANSMITTER.state [1]), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state [0]), .O(n10365));   // coms.v(280[12] 380[6])
    defparam i8005_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i8367_3_lut (.I0(\data_out_frame2[5] [2]), .I1(rand_data[26]), 
            .I2(n10197), .I3(GND_net), .O(n10727));   // coms.v(426[12] 547[6])
    defparam i8367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8415_3_lut (.I0(\data_out_frame2[11] [2]), .I1(rand_data[10]), 
            .I2(n10197), .I3(GND_net), .O(n10775));   // coms.v(426[12] 547[6])
    defparam i8415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_3_lut_adj_803 (.I0(r_Clock_Count[8]), .I1(n17537), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16459));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_803.LUT_INIT = 16'hacac;
    SB_LUT4 i8368_3_lut (.I0(\data_out_frame2[5] [3]), .I1(rand_data[27]), 
            .I2(n10197), .I3(GND_net), .O(n10728));   // coms.v(426[12] 547[6])
    defparam i8368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_3_lut_adj_804 (.I0(r_Clock_Count[7]), .I1(n17641), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16467));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_804.LUT_INIT = 16'hacac;
    SB_LUT4 i31_3_lut_adj_805 (.I0(r_Clock_Count_adj_2510[2]), .I1(n17570), 
            .I2(r_SM_Main_adj_2509[2]), .I3(GND_net), .O(n16675));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31_3_lut_adj_805.LUT_INIT = 16'hacac;
    SB_LUT4 i25_3_lut_adj_806 (.I0(r_Clock_Count[6]), .I1(n17636), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16477));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i25_3_lut_adj_806.LUT_INIT = 16'hacac;
    SB_CARRY rand_setpoint_2351_add_4_26 (.CI(n15582), .I0(rand_data[24]), 
            .I1(rand_setpoint[24]), .CO(n15583));
    SB_LUT4 i8450_3_lut (.I0(\data_out_frame2[15] [5]), .I1(rand_data[13]), 
            .I2(n10197), .I3(GND_net), .O(n10810));   // coms.v(426[12] 547[6])
    defparam i8450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rand_setpoint_2351_add_4_25_lut (.I0(GND_net), .I1(rand_data[23]), 
            .I2(rand_setpoint[23]), .I3(n15581), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_12 (.CI(n15537), .I0(GND_net), .I1(rand_data[10]), 
            .CO(n15538));
    SB_LUT4 i8416_3_lut (.I0(\data_out_frame2[11] [3]), .I1(rand_data[11]), 
            .I2(n10197), .I3(GND_net), .O(n10776));   // coms.v(426[12] 547[6])
    defparam i8416_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rand_setpoint_2351_add_4_25 (.CI(n15581), .I0(rand_data[23]), 
            .I1(rand_setpoint[23]), .CO(n15582));
    SB_CARRY rand_data_2350_add_4_30 (.CI(n15555), .I0(GND_net), .I1(rand_data[28]), 
            .CO(n15556));
    SB_LUT4 rand_data_2350_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[27]), 
            .I3(n15554), .O(n138_adj_2466)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_29 (.CI(n15554), .I0(GND_net), .I1(rand_data[27]), 
            .CO(n15555));
    SB_LUT4 rand_setpoint_2351_add_4_24_lut (.I0(GND_net), .I1(rand_data[22]), 
            .I2(rand_setpoint[22]), .I3(n15580), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rand_data_2350_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[26]), 
            .I3(n15553), .O(n139_adj_2467)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_28_lut.LUT_INIT = 16'hC33C;
    coms c0 (.n10793(n10793), .\data_out_frame2[13] ({\data_out_frame2[13] }), 
         .CLK_c(CLK_c), .n10792(n10792), .n10791(n10791), .n10790(n10790), 
         .rx_data({rx_data}), .n10789(n10789), .n10788(n10788), .\data_out_frame2[12] ({\data_out_frame2[12] }), 
         .n10787(n10787), .n10786(n10786), .n10785(n10785), .n10784(n10784), 
         .GND_net(GND_net), .\data_out_frame2[17] ({\data_out_frame2[17] }), 
         .\data_out_frame2[16] ({\data_out_frame2[16] }), .n12933(n12933), 
         .n127(n127), .n9435(n9435), .n10783(n10783), .\data_out_frame2[6] ({\data_out_frame2[6] }), 
         .\data_out_frame2[7] ({\data_out_frame2[7] }), .\FRAME_MATCHER.state ({Open_0, 
         Open_1, Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, 
         Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
         Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
         Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, 
         \FRAME_MATCHER.state [2], Open_29, Open_30}), .\data_out[8] ({Open_31, 
         Open_32, Open_33, Open_34, Open_35, Open_36, \data_out[8] [1:0]}), 
         .\byte_transmit_counter[3] (byte_transmit_counter[3]), .\data_out[0][1] (\data_out[0] [1]), 
         .\data_out_frame2[5] ({\data_out_frame2[5] }), .n10782(n10782), 
         .\data_out_frame2[10] ({\data_out_frame2[10] }), .\data_out_frame2[11] ({\data_out_frame2[11] }), 
         .n10781(n10781), .n10780(n10780), .n10779(n10779), .n1716(n1716), 
         .n10373(n10373), .n10778(n10778), .n10777(n10777), .n10776(n10776), 
         .n10775(n10775), .n10774(n10774), .n10773(n10773), .tx_active(tx_active), 
         .n10772(n10772), .n10771(n10771), .n10770(n10770), .n10769(n10769), 
         .n4445(n4445), .n10768(n10768), .n10767(n10767), .n10766(n10766), 
         .n10765(n10765), .n10055(n10055), .\data_out_frame2[9] ({\data_out_frame2[9] }), 
         .\data_out_frame2[8] ({\data_out_frame2[8] }), .\data_out[1][7] (\data_out[1] [7]), 
         .n10764(n10764), .\data_out[2][7] (\data_out[2] [7]), .\data_out[3][7] (\data_out[3] [7]), 
         .n10372(n10372), .\data_out[0][3] (\data_out[0] [3]), .n10763(n10763), 
         .n10371(n10371), .\data_out[0][5] (\data_out[0] [5]), .n10762(n10762), 
         .n10761(n10761), .n10760(n10760), .n2275(n2275), .n10759(n10759), 
         .n10758(n10758), .n10836(n10836), .\data_out_frame2[18] ({\data_out_frame2[18] }), 
         .n10835(n10835), .n10834(n10834), .n10833(n10833), .n10832(n10832), 
         .n10757(n10757), .n10816(n10816), .n10756(n10756), .n10815(n10815), 
         .n10755(n10755), .n10814(n10814), .n10754(n10754), .n10813(n10813), 
         .n10753(n10753), .n10812(n10812), .\data_out_frame2[15] ({\data_out_frame2[15] }), 
         .n10811(n10811), .n10810(n10810), .n10809(n10809), .n10808(n10808), 
         .n10807(n10807), .n10806(n10806), .n10805(n10805), .n10804(n10804), 
         .\data_out_frame2[14] ({\data_out_frame2[14] }), .n10803(n10803), 
         .n10802(n10802), .n10752(n10752), .n10801(n10801), .n10751(n10751), 
         .n10800(n10800), .n10750(n10750), .n10799(n10799), .n10749(n10749), 
         .n10798(n10798), .n10748(n10748), .n10797(n10797), .n10747(n10747), 
         .n10796(n10796), .n10746(n10746), .n10745(n10745), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .r_Tx_Data({r_Tx_Data}), .n8730(n8730), .\byte_transmit_counter[4] (byte_transmit_counter[4]), 
         .n10744(n10744), .n10743(n10743), .n10742(n10742), .n9460(n9460), 
         .\FRAME_MATCHER.state[1] (\FRAME_MATCHER.state [1]), .n10741(n10741), 
         .n16795(n16795), .n10740(n10740), .n10739(n10739), .n10738(n10738), 
         .n10737(n10737), .n10736(n10736), .n10735(n10735), .n10734(n10734), 
         .n10733(n10733), .n10732(n10732), .n10731(n10731), .n10730(n10730), 
         .n10729(n10729), .n10728(n10728), .n10727(n10727), .n10726(n10726), 
         .n10725(n10725), .n16255(n16255), .\UART_TRANSMITTER.state[1] (\UART_TRANSMITTER.state [1]), 
         .\data_in[1] ({\data_in[1] }), .\data_in[3] ({\data_in[3] }), .\UART_TRANSMITTER.state[0] (\UART_TRANSMITTER.state [0]), 
         .n2546({n2547}), .n1651(n1651), .n9453(n9453), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .\data_in_frame[0] ({\data_in_frame[0] }), .n16607(n16607), .VCC_net(VCC_net), 
         .\data_out[6][0] (\data_out[6] [0]), .n18137(n18137), .n16797(n16797), 
         .n10698(n10698), .n10697(n10697), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n10695(n10695), .n10693(n10693), .\data_out[8][4] (\data_out[8] [4]), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in[2] ({\data_in[2] }), 
         .\data_in[0] ({\data_in[0] }), .n3977(n3977), .\data_out[9][2] (\data_out[9] [2]), 
         .n127_adj_4(n127_adj_2418), .n10692(n10692), .\data_out[8][5] (\data_out[8] [5]), 
         .n10691(n10691), .\data_out[8][6] (\data_out[8] [6]), .n9445(n9445), 
         .n10690(n10690), .\data_out[8][7] (\data_out[8] [7]), .n10831(n10831), 
         .n10830(n10830), .n10829(n10829), .n10689(n10689), .n10828(n10828), 
         .n10688(n10688), .n10687(n10687), .n10686(n10686), .n10685(n10685), 
         .n10684(n10684), .n10683(n10683), .n10682(n10682), .n10681(n10681), 
         .n10680(n10680), .n10679(n10679), .n10678(n10678), .n10677(n10677), 
         .n10676(n10676), .n10827(n10827), .n10(n10_adj_2426), .n10675(n10675), 
         .data_out_9__2__N_367(data_out_9__2__N_367), .\UART_TRANSMITTER.state[2] (\UART_TRANSMITTER.state [2]), 
         .n10674(n10674), .n10826(n10826), .n10_adj_5(n10_adj_2425), .n16886(n16886), 
         .n9361(n9361), .n9452(n9452), .n10_adj_6(n10_adj_2427), .n10673(n10673), 
         .n10_adj_7(n10_adj_2423), .n10825(n10825), .n10672(n10672), .n29(n29), 
         .n10671(n10671), .n10670(n10670), .n10367(n10367), .\data_out[1][6] (\data_out[1] [6]), 
         .n10669(n10669), .n10668(n10668), .n10667(n10667), .n10366(n10366), 
         .n10666(n10666), .n10665(n10665), .n10664(n10664), .n2651({n2652}), 
         .n10663(n10663), .n10662(n10662), .n10661(n10661), .n10660(n10660), 
         .n10659(n10659), .n10658(n10658), .n18044(n18044), .n10365(n10365), 
         .\data_out[2][0] (\data_out[2] [0]), .\rand_setpoint[25] (rand_setpoint[25]), 
         .\rand_setpoint[17] (rand_setpoint[17]), .n10364(n10364), .\data_out[2][2] (\data_out[2] [2]), 
         .\rand_setpoint[18] (rand_setpoint[18]), .\rand_setpoint[19] (rand_setpoint[19]), 
         .n33(n33), .\rand_setpoint[20] (rand_setpoint[20]), .n53(n53), 
         .n491(n491), .\rand_setpoint[21] (rand_setpoint[21]), .\rand_setpoint[22] (rand_setpoint[22]), 
         .\rand_setpoint[23] (rand_setpoint[23]), .\rand_setpoint[8] (rand_setpoint[8]), 
         .n9462(n9462), .data_out_10__7__N_110(data_out_10__7__N_110), .\rand_setpoint[2] (rand_setpoint[2]), 
         .\rand_setpoint[3] (rand_setpoint[3]), .n7198(n7198), .n10625(n10625), 
         .n10624(n10624), .n10623(n10623), .n10622(n10622), .n10621(n10621), 
         .n10362(n10362), .\data_out[2][5] (\data_out[2] [5]), .n10361(n10361), 
         .n10360(n10360), .\data_out[3][0] (\data_out[3] [0]), .n10620(n10620), 
         .n10619(n10619), .n10359(n10359), .\data_out[3][2] (\data_out[3] [2]), 
         .n10358(n10358), .\data_out[3][4] (\data_out[3] [4]), .\data_out[3][5] (\data_out[3] [5]), 
         .n10357(n10357), .\rand_setpoint[30] (rand_setpoint[30]), .n17230(n17230), 
         .\rand_setpoint[29] (rand_setpoint[29]), .n10355(n10355), .n18038(n18038), 
         .\rand_setpoint[9] (rand_setpoint[9]), .n9357(n9357), .n445(n445), 
         .\rand_setpoint[10] (rand_setpoint[10]), .n18032(n18032), .n10824(n10824), 
         .n10823(n10823), .n10599(n10599), .n10598(n10598), .n10597(n10597), 
         .n10596(n10596), .n10592(n10592), .n10591(n10591), .n10590(n10590), 
         .n10589(n10589), .n10588(n10588), .n10584(n10584), .n10583(n10583), 
         .n10582(n10582), .n10577(n10577), .n10576(n10576), .n10575(n10575), 
         .n10574(n10574), .n16259(n16259), .n10822(n10822), .\rand_setpoint[11] (rand_setpoint[11]), 
         .n10821(n10821), .n10820(n10820), .n18026(n18026), .n10819(n10819), 
         .n10818(n10818), .\rand_setpoint[28] (rand_setpoint[28]), .\FRAME_MATCHER.state_31__N_1440[1] (\FRAME_MATCHER.state_31__N_1440 [1]), 
         .n10817(n10817), .\rand_setpoint[13] (rand_setpoint[13]), .\rand_setpoint[14] (rand_setpoint[14]), 
         .\rand_setpoint[15] (rand_setpoint[15]), .\rand_setpoint[12] (rand_setpoint[12]), 
         .n16897(n16897), .n31(n31), .n10197(n10197), .n10795(n10795), 
         .n16893(n16893), .n16896(n16896), .\rand_setpoint[27] (rand_setpoint[27]), 
         .\rand_setpoint[26] (rand_setpoint[26]), .\data_out[0][0] (\data_out[0] [0]), 
         .n10031(n10031), .\rand_setpoint[24] (rand_setpoint[24]), .n9358(n9358), 
         .rx_data_ready(rx_data_ready), .n10141(n10141), .\rand_setpoint[31] (rand_setpoint[31]), 
         .n10794(n10794), .n10392(n10392), .n16327(n16327), .n10374(n10374), 
         .n8828(n8828), .r_SM_Main({r_SM_Main}), .n3(n3_adj_2406), .\r_Bit_Index[1] (r_Bit_Index[1]), 
         .n14060(n14060), .n5(n5), .n13276(n13276), .n16671(n16671), 
         .r_Clock_Count({r_Clock_Count}), .n16651(n16651), .n16649(n16649), 
         .n16567(n16567), .n16509(n16509), .n16477(n16477), .n16467(n16467), 
         .n16459(n16459), .n16625(n16625), .n17537(n17537), .n16844(n16844), 
         .n17641(n17641), .n17636(n17636), .n17631(n17631), .n16828(n16828), 
         .n17573(n17573), .n17494(n17494), .n17484(n17484), .n17461(n17461), 
         .n17542(n17542), .n15701(n15701), .n10580(n10580), .n10579(n10579), 
         .n10578(n10578), .tx_o(tx_o), .n9406(n9406), .n4(n4_adj_2458), 
         .n12(n12), .n16627(n16627), .n16629(n16629), .n9937(n9937), 
         .n16683(n16683), .n16681(n16681), .n17395(n17395), .n17394(n17394), 
         .n17397(n17397), .n17398(n17398), .tx_enable(tx_enable), .r_Bit_Index({r_Bit_Index_adj_2511}), 
         .r_SM_Main_adj_41({r_SM_Main_adj_2509}), .n3_adj_12(n3), .\r_SM_Main_2__N_2033[1] (r_SM_Main_2__N_2033_adj_2515[1]), 
         .n7866(n7866), .n16463(n16463), .r_Clock_Count_adj_42({r_Clock_Count_adj_2510}), 
         .n10714(n10714), .n10607(n10607), .n17458(n17458), .n16824(n16824), 
         .n17640(n17640), .n17634(n17634), .n17629(n17629), .n16817(n16817), 
         .n16677(n16677), .n17567(n17567), .n16623(n16623), .n17457(n17457), 
         .n16675(n16675), .n17570(n17570), .n17504(n17504), .n17544(n17544), 
         .n16673(n16673), .n16577(n16577), .n16517(n16517), .n9403(n9403), 
         .n16483(n16483), .n10587(n10587), .n10585(n10585), .tx2_o(tx2_o), 
         .n15837(n15837), .n16473(n16473), .n10396(n10396), .n10399(n10399), 
         .n9929(n9929), .n12_adj_22(n12_adj_2410), .n5029(n5029), .n17194(n17194), 
         .n10398(n10398), .n15689(n15689), .tx2_enable(tx2_enable), .r_Rx_Data(r_Rx_Data), 
         .r_SM_Main_adj_43({r_SM_Main_adj_2506}), .n1(n1), .r_Clock_Count_adj_44({r_Clock_Count_adj_2504}), 
         .n16863(n16863), .n16575(n16575), .n17222(n17222), .n16573(n16573), 
         .n16571(n16571), .r_Bit_Index_adj_45({r_Bit_Index_adj_2505}), .n13082(n13082), 
         .n4_adj_37(n4_adj_2417), .n16569(n16569), .n4_adj_38(n4_adj_2460), 
         .n9472(n9472), .n16515(n16515), .n16479(n16479), .n16469(n16469), 
         .n13510(n13510), .rx_i(rx_i), .n10631(n10631), .n16547(n16547), 
         .n16855(n16855), .n16852(n16852), .n16856(n16856), .n16857(n16857), 
         .n16854(n16854), .n16858(n16858), .n16860(n16860), .n16853(n16853), 
         .n10635(n10635), .n16859(n16859), .n4_adj_39(n4_adj_2411), .n17260(n17260), 
         .n17602(n17602), .n17601(n17601), .n10581(n10581), .n9477(n9477), 
         .n4_adj_40(n4_adj_2409), .n6(n6_adj_2461), .n10423(n10423), .n10426(n10426), 
         .n16867(n16867), .n10433(n10433), .n10432(n10432), .n10431(n10431), 
         .n10430(n10430), .n10429(n10429), .n10428(n10428), .n10427(n10427), 
         .n13440(n13440), .n10425(n10425)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(84[8] 97[4])
    SB_CARRY rand_setpoint_2351_add_4_24 (.CI(n15580), .I0(rand_data[22]), 
            .I1(rand_setpoint[22]), .CO(n15581));
    SB_LUT4 rand_setpoint_2351_add_4_23_lut (.I0(GND_net), .I1(rand_data[21]), 
            .I2(rand_setpoint[21]), .I3(n15579), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14724_2_lut (.I0(\UART_TRANSMITTER.state [1]), .I1(n9361), 
            .I2(GND_net), .I3(GND_net), .O(n17162));
    defparam i14724_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY rand_setpoint_2351_add_4_23 (.CI(n15579), .I0(rand_data[21]), 
            .I1(rand_setpoint[21]), .CO(n15580));
    SB_LUT4 rand_setpoint_2351_add_4_22_lut (.I0(GND_net), .I1(rand_data[20]), 
            .I2(rand_setpoint[20]), .I3(n15578), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_setpoint_2351_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_data_2350_add_4_28 (.CI(n15553), .I0(GND_net), .I1(rand_data[26]), 
            .CO(n15554));
    SB_LUT4 rand_data_2350_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(rand_data[25]), 
            .I3(n15552), .O(n140_adj_2468)) /* synthesis syn_instantiated=1 */ ;
    defparam rand_data_2350_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rand_setpoint_2351_add_4_22 (.CI(n15578), .I0(rand_data[20]), 
            .I1(rand_setpoint[20]), .CO(n15579));
    
endmodule
//
// Verilog Description of module coms
//

module coms (n10793, \data_out_frame2[13] , CLK_c, n10792, n10791, 
            n10790, rx_data, n10789, n10788, \data_out_frame2[12] , 
            n10787, n10786, n10785, n10784, GND_net, \data_out_frame2[17] , 
            \data_out_frame2[16] , n12933, n127, n9435, n10783, \data_out_frame2[6] , 
            \data_out_frame2[7] , \FRAME_MATCHER.state , \data_out[8] , 
            \byte_transmit_counter[3] , \data_out[0][1] , \data_out_frame2[5] , 
            n10782, \data_out_frame2[10] , \data_out_frame2[11] , n10781, 
            n10780, n10779, n1716, n10373, n10778, n10777, n10776, 
            n10775, n10774, n10773, tx_active, n10772, n10771, n10770, 
            n10769, n4445, n10768, n10767, n10766, n10765, n10055, 
            \data_out_frame2[9] , \data_out_frame2[8] , \data_out[1][7] , 
            n10764, \data_out[2][7] , \data_out[3][7] , n10372, \data_out[0][3] , 
            n10763, n10371, \data_out[0][5] , n10762, n10761, n10760, 
            n2275, n10759, n10758, n10836, \data_out_frame2[18] , 
            n10835, n10834, n10833, n10832, n10757, n10816, n10756, 
            n10815, n10755, n10814, n10754, n10813, n10753, n10812, 
            \data_out_frame2[15] , n10811, n10810, n10809, n10808, 
            n10807, n10806, n10805, n10804, \data_out_frame2[14] , 
            n10803, n10802, n10752, n10801, n10751, n10800, n10750, 
            n10799, n10749, n10798, n10748, n10797, n10747, n10796, 
            n10746, n10745, \byte_transmit_counter[2] , r_Tx_Data, n8730, 
            \byte_transmit_counter[4] , n10744, n10743, n10742, n9460, 
            \FRAME_MATCHER.state[1] , n10741, n16795, n10740, n10739, 
            n10738, n10737, n10736, n10735, n10734, n10733, n10732, 
            n10731, n10730, n10729, n10728, n10727, n10726, n10725, 
            n16255, \UART_TRANSMITTER.state[1] , \data_in[1] , \data_in[3] , 
            \UART_TRANSMITTER.state[0] , n2546, n1651, n9453, \FRAME_MATCHER.state[0] , 
            \data_in_frame[0] , n16607, VCC_net, \data_out[6][0] , n18137, 
            n16797, n10698, n10697, \data_in_frame[7] , n10695, n10693, 
            \data_out[8][4] , \data_in_frame[6] , \data_in[2] , \data_in[0] , 
            n3977, \data_out[9][2] , n127_adj_4, n10692, \data_out[8][5] , 
            n10691, \data_out[8][6] , n9445, n10690, \data_out[8][7] , 
            n10831, n10830, n10829, n10689, n10828, n10688, n10687, 
            n10686, n10685, n10684, n10683, n10682, n10681, n10680, 
            n10679, n10678, n10677, n10676, n10827, n10, n10675, 
            data_out_9__2__N_367, \UART_TRANSMITTER.state[2] , n10674, 
            n10826, n10_adj_5, n16886, n9361, n9452, n10_adj_6, 
            n10673, n10_adj_7, n10825, n10672, n29, n10671, n10670, 
            n10367, \data_out[1][6] , n10669, n10668, n10667, n10366, 
            n10666, n10665, n10664, n2651, n10663, n10662, n10661, 
            n10660, n10659, n10658, n18044, n10365, \data_out[2][0] , 
            \rand_setpoint[25] , \rand_setpoint[17] , n10364, \data_out[2][2] , 
            \rand_setpoint[18] , \rand_setpoint[19] , n33, \rand_setpoint[20] , 
            n53, n491, \rand_setpoint[21] , \rand_setpoint[22] , \rand_setpoint[23] , 
            \rand_setpoint[8] , n9462, data_out_10__7__N_110, \rand_setpoint[2] , 
            \rand_setpoint[3] , n7198, n10625, n10624, n10623, n10622, 
            n10621, n10362, \data_out[2][5] , n10361, n10360, \data_out[3][0] , 
            n10620, n10619, n10359, \data_out[3][2] , n10358, \data_out[3][4] , 
            \data_out[3][5] , n10357, \rand_setpoint[30] , n17230, \rand_setpoint[29] , 
            n10355, n18038, \rand_setpoint[9] , n9357, n445, \rand_setpoint[10] , 
            n18032, n10824, n10823, n10599, n10598, n10597, n10596, 
            n10592, n10591, n10590, n10589, n10588, n10584, n10583, 
            n10582, n10577, n10576, n10575, n10574, n16259, n10822, 
            \rand_setpoint[11] , n10821, n10820, n18026, n10819, n10818, 
            \rand_setpoint[28] , \FRAME_MATCHER.state_31__N_1440[1] , n10817, 
            \rand_setpoint[13] , \rand_setpoint[14] , \rand_setpoint[15] , 
            \rand_setpoint[12] , n16897, n31, n10197, n10795, n16893, 
            n16896, \rand_setpoint[27] , \rand_setpoint[26] , \data_out[0][0] , 
            n10031, \rand_setpoint[24] , n9358, rx_data_ready, n10141, 
            \rand_setpoint[31] , n10794, n10392, n16327, n10374, n8828, 
            r_SM_Main, n3, \r_Bit_Index[1] , n14060, n5, n13276, 
            n16671, r_Clock_Count, n16651, n16649, n16567, n16509, 
            n16477, n16467, n16459, n16625, n17537, n16844, n17641, 
            n17636, n17631, n16828, n17573, n17494, n17484, n17461, 
            n17542, n15701, n10580, n10579, n10578, tx_o, n9406, 
            n4, n12, n16627, n16629, n9937, n16683, n16681, n17395, 
            n17394, n17397, n17398, tx_enable, r_Bit_Index, r_SM_Main_adj_41, 
            n3_adj_12, \r_SM_Main_2__N_2033[1] , n7866, n16463, r_Clock_Count_adj_42, 
            n10714, n10607, n17458, n16824, n17640, n17634, n17629, 
            n16817, n16677, n17567, n16623, n17457, n16675, n17570, 
            n17504, n17544, n16673, n16577, n16517, n9403, n16483, 
            n10587, n10585, tx2_o, n15837, n16473, n10396, n10399, 
            n9929, n12_adj_22, n5029, n17194, n10398, n15689, tx2_enable, 
            r_Rx_Data, r_SM_Main_adj_43, n1, r_Clock_Count_adj_44, n16863, 
            n16575, n17222, n16573, n16571, r_Bit_Index_adj_45, n13082, 
            n4_adj_37, n16569, n4_adj_38, n9472, n16515, n16479, 
            n16469, n13510, rx_i, n10631, n16547, n16855, n16852, 
            n16856, n16857, n16854, n16858, n16860, n16853, n10635, 
            n16859, n4_adj_39, n17260, n17602, n17601, n10581, n9477, 
            n4_adj_40, n6, n10423, n10426, n16867, n10433, n10432, 
            n10431, n10430, n10429, n10428, n10427, n13440, n10425) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n10793;
    output [7:0]\data_out_frame2[13] ;
    input CLK_c;
    input n10792;
    input n10791;
    input n10790;
    output [7:0]rx_data;
    input n10789;
    input n10788;
    output [7:0]\data_out_frame2[12] ;
    input n10787;
    input n10786;
    input n10785;
    input n10784;
    input GND_net;
    output [7:0]\data_out_frame2[17] ;
    output [7:0]\data_out_frame2[16] ;
    output n12933;
    output n127;
    output n9435;
    input n10783;
    output [7:0]\data_out_frame2[6] ;
    output [7:0]\data_out_frame2[7] ;
    output [31:0]\FRAME_MATCHER.state ;
    output [7:0]\data_out[8] ;
    output \byte_transmit_counter[3] ;
    output \data_out[0][1] ;
    output [7:0]\data_out_frame2[5] ;
    input n10782;
    output [7:0]\data_out_frame2[10] ;
    output [7:0]\data_out_frame2[11] ;
    input n10781;
    input n10780;
    input n10779;
    output n1716;
    input n10373;
    input n10778;
    input n10777;
    input n10776;
    input n10775;
    input n10774;
    input n10773;
    output tx_active;
    input n10772;
    input n10771;
    input n10770;
    input n10769;
    input n4445;
    input n10768;
    input n10767;
    input n10766;
    input n10765;
    output n10055;
    output [7:0]\data_out_frame2[9] ;
    output [7:0]\data_out_frame2[8] ;
    output \data_out[1][7] ;
    input n10764;
    output \data_out[2][7] ;
    output \data_out[3][7] ;
    input n10372;
    output \data_out[0][3] ;
    input n10763;
    input n10371;
    output \data_out[0][5] ;
    input n10762;
    input n10761;
    input n10760;
    output n2275;
    input n10759;
    input n10758;
    input n10836;
    output [7:0]\data_out_frame2[18] ;
    input n10835;
    input n10834;
    input n10833;
    input n10832;
    input n10757;
    input n10816;
    input n10756;
    input n10815;
    input n10755;
    input n10814;
    input n10754;
    input n10813;
    input n10753;
    input n10812;
    output [7:0]\data_out_frame2[15] ;
    input n10811;
    input n10810;
    input n10809;
    input n10808;
    input n10807;
    input n10806;
    input n10805;
    input n10804;
    output [7:0]\data_out_frame2[14] ;
    input n10803;
    input n10802;
    input n10752;
    input n10801;
    input n10751;
    input n10800;
    input n10750;
    input n10799;
    input n10749;
    input n10798;
    input n10748;
    input n10797;
    input n10747;
    input n10796;
    input n10746;
    input n10745;
    output \byte_transmit_counter[2] ;
    output [7:0]r_Tx_Data;
    output n8730;
    output \byte_transmit_counter[4] ;
    input n10744;
    input n10743;
    input n10742;
    output n9460;
    output \FRAME_MATCHER.state[1] ;
    input n10741;
    output n16795;
    input n10740;
    input n10739;
    input n10738;
    input n10737;
    input n10736;
    input n10735;
    input n10734;
    input n10733;
    input n10732;
    input n10731;
    input n10730;
    input n10729;
    input n10728;
    input n10727;
    input n10726;
    input n10725;
    input n16255;
    output \UART_TRANSMITTER.state[1] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[3] ;
    output \UART_TRANSMITTER.state[0] ;
    output [0:0]n2546;
    output n1651;
    output n9453;
    output \FRAME_MATCHER.state[0] ;
    output [7:0]\data_in_frame[0] ;
    input n16607;
    input VCC_net;
    output \data_out[6][0] ;
    input n18137;
    input n16797;
    input n10698;
    input n10697;
    output [7:0]\data_in_frame[7] ;
    input n10695;
    input n10693;
    output \data_out[8][4] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[0] ;
    output n3977;
    output \data_out[9][2] ;
    output n127_adj_4;
    input n10692;
    output \data_out[8][5] ;
    input n10691;
    output \data_out[8][6] ;
    output n9445;
    input n10690;
    output \data_out[8][7] ;
    input n10831;
    input n10830;
    input n10829;
    input n10689;
    input n10828;
    input n10688;
    input n10687;
    input n10686;
    input n10685;
    input n10684;
    input n10683;
    input n10682;
    input n10681;
    input n10680;
    input n10679;
    input n10678;
    input n10677;
    input n10676;
    input n10827;
    output n10;
    input n10675;
    output data_out_9__2__N_367;
    output \UART_TRANSMITTER.state[2] ;
    input n10674;
    input n10826;
    output n10_adj_5;
    output n16886;
    output n9361;
    output n9452;
    output n10_adj_6;
    input n10673;
    output n10_adj_7;
    input n10825;
    input n10672;
    output n29;
    input n10671;
    input n10670;
    input n10367;
    output \data_out[1][6] ;
    input n10669;
    input n10668;
    input n10667;
    input n10366;
    input n10666;
    input n10665;
    input n10664;
    output [0:0]n2651;
    input n10663;
    input n10662;
    input n10661;
    input n10660;
    input n10659;
    input n10658;
    output n18044;
    input n10365;
    output \data_out[2][0] ;
    input \rand_setpoint[25] ;
    input \rand_setpoint[17] ;
    input n10364;
    output \data_out[2][2] ;
    input \rand_setpoint[18] ;
    input \rand_setpoint[19] ;
    input n33;
    input \rand_setpoint[20] ;
    input n53;
    output n491;
    input \rand_setpoint[21] ;
    input \rand_setpoint[22] ;
    input \rand_setpoint[23] ;
    input \rand_setpoint[8] ;
    output n9462;
    output data_out_10__7__N_110;
    input \rand_setpoint[2] ;
    input \rand_setpoint[3] ;
    output n7198;
    input n10625;
    input n10624;
    input n10623;
    input n10622;
    input n10621;
    input n10362;
    output \data_out[2][5] ;
    input n10361;
    input n10360;
    output \data_out[3][0] ;
    input n10620;
    input n10619;
    input n10359;
    output \data_out[3][2] ;
    input n10358;
    output \data_out[3][4] ;
    output \data_out[3][5] ;
    input n10357;
    input \rand_setpoint[30] ;
    output n17230;
    input \rand_setpoint[29] ;
    input n10355;
    output n18038;
    input \rand_setpoint[9] ;
    output n9357;
    output n445;
    input \rand_setpoint[10] ;
    output n18032;
    input n10824;
    input n10823;
    input n10599;
    input n10598;
    input n10597;
    input n10596;
    input n10592;
    input n10591;
    input n10590;
    input n10589;
    input n10588;
    input n10584;
    input n10583;
    input n10582;
    input n10577;
    input n10576;
    input n10575;
    input n10574;
    input n16259;
    input n10822;
    input \rand_setpoint[11] ;
    input n10821;
    input n10820;
    output n18026;
    input n10819;
    input n10818;
    input \rand_setpoint[28] ;
    output \FRAME_MATCHER.state_31__N_1440[1] ;
    input n10817;
    input \rand_setpoint[13] ;
    input \rand_setpoint[14] ;
    input \rand_setpoint[15] ;
    input \rand_setpoint[12] ;
    output n16897;
    output n31;
    output n10197;
    input n10795;
    output n16893;
    output n16896;
    input \rand_setpoint[27] ;
    input \rand_setpoint[26] ;
    output \data_out[0][0] ;
    output n10031;
    input \rand_setpoint[24] ;
    output n9358;
    output rx_data_ready;
    output n10141;
    input \rand_setpoint[31] ;
    input n10794;
    input n10392;
    input n16327;
    input n10374;
    output n8828;
    output [2:0]r_SM_Main;
    output n3;
    output \r_Bit_Index[1] ;
    output n14060;
    output n5;
    output n13276;
    input n16671;
    output [8:0]r_Clock_Count;
    input n16651;
    input n16649;
    input n16567;
    input n16509;
    input n16477;
    input n16467;
    input n16459;
    input n16625;
    output n17537;
    input n16844;
    output n17641;
    output n17636;
    output n17631;
    input n16828;
    output n17573;
    output n17494;
    output n17484;
    output n17461;
    output n17542;
    output n15701;
    input n10580;
    input n10579;
    input n10578;
    output tx_o;
    output n9406;
    output n4;
    output n12;
    input n16627;
    input n16629;
    output n9937;
    input n16683;
    input n16681;
    input n17395;
    input n17394;
    input n17397;
    input n17398;
    output tx_enable;
    output [2:0]r_Bit_Index;
    output [2:0]r_SM_Main_adj_41;
    output n3_adj_12;
    output \r_SM_Main_2__N_2033[1] ;
    output n7866;
    input n16463;
    output [8:0]r_Clock_Count_adj_42;
    input n10714;
    input n10607;
    output n17458;
    input n16824;
    output n17640;
    output n17634;
    output n17629;
    input n16817;
    input n16677;
    output n17567;
    input n16623;
    output n17457;
    input n16675;
    output n17570;
    output n17504;
    output n17544;
    input n16673;
    input n16577;
    input n16517;
    output n9403;
    input n16483;
    input n10587;
    input n10585;
    output tx2_o;
    output n15837;
    input n16473;
    input n10396;
    input n10399;
    output n9929;
    output n12_adj_22;
    output n5029;
    output n17194;
    output n10398;
    input n15689;
    output tx2_enable;
    output r_Rx_Data;
    output [2:0]r_SM_Main_adj_43;
    output n1;
    output [7:0]r_Clock_Count_adj_44;
    output n16863;
    input n16575;
    output n17222;
    input n16573;
    input n16571;
    output [2:0]r_Bit_Index_adj_45;
    output n13082;
    output n4_adj_37;
    input n16569;
    output n4_adj_38;
    output n9472;
    input n16515;
    input n16479;
    input n16469;
    input n13510;
    input rx_i;
    input n10631;
    input n16547;
    output n16855;
    input n16852;
    output n16856;
    output n16857;
    output n16854;
    output n16858;
    output n16860;
    output n16853;
    input n10635;
    output n16859;
    output n4_adj_39;
    output n17260;
    output n17602;
    output n17601;
    input n10581;
    output n9477;
    output n4_adj_40;
    output n6;
    input n10423;
    input n10426;
    output n16867;
    input n10433;
    input n10432;
    input n10431;
    input n10430;
    input n10429;
    input n10428;
    input n10427;
    output n13440;
    output n10425;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n8, n16882;
    wire [7:0]\data_in_frame[10] ;   // coms.v(389[12:25])
    
    wire n10377, n10470;
    wire [14:0]delay_counter;   // coms.v(272[12:25])
    wire [7:0]\data_out_frame2[0] ;   // coms.v(390[12:27])
    wire [7:0]byte_transmit_counter2;   // coms.v(409[12:34])
    
    wire n17579, n17999, n18002, n2, n4_c, n5_c, n17454, n17452, 
        n9451, n7;
    wire [31:0]\FRAME_MATCHER.state_c ;   // coms.v(419[11:16])
    
    wire n16377, n16383;
    wire [7:0]byte_transmit_counter;   // coms.v(19[11:32])
    wire [7:0]\data_out[9] ;   // coms.v(21[11:19])
    
    wire n18077;
    wire [7:0]\data_out[1] ;   // coms.v(21[11:19])
    
    wire n18080, n6_c, n18071;
    wire [7:0]n37;
    
    wire n15618, n127_adj_2136, n15619, n10473, n17969, n17972, 
        tx_active_prev, n15617, n16838;
    wire [2:0]r_SM_Main_2__N_2036;
    wire [0:0]n1846;
    
    wire n10054;
    wire [7:0]\data_out[7] ;   // coms.v(21[11:19])
    wire [0:0]n1881;
    wire [0:0]n1916;
    wire [0:0]n1951;
    wire [0:0]n1986;
    wire [7:0]\data_out[6] ;   // coms.v(21[11:19])
    wire [0:0]n2021;
    wire [0:0]n2056;
    wire [0:0]n2091;
    wire [0:0]n2126;
    wire [0:0]n2161;
    wire [0:0]n2196;
    wire [0:0]n2476;
    wire [7:0]\data_out[5] ;   // coms.v(21[11:19])
    
    wire n18074, n17585;
    wire [0:0]n3071;
    
    wire n2_adj_2137, n10370;
    wire [7:0]\data_out[0] ;   // coms.v(21[11:19])
    wire [31:0]\FRAME_MATCHER.i ;   // coms.v(422[11:12])
    
    wire n9346, n10867, n10479, n10865, n10485, n10488, n10491, 
        n10494, n8_adj_2138;
    wire [7:0]\data_out[10] ;   // coms.v(21[11:19])
    
    wire n10_c, n18098, n10_adj_2139, n16595, n10860, n47, n56, 
        n60, n33_c, n17258, n28, n9, n18065, n6_adj_2140, n10378, 
        n18068, n16905, n16879;
    wire [7:0]\data_out_frame2[19] ;   // coms.v(390[12:27])
    
    wire n18059, n17240, n9490, n9482, n15616, n10052, n10297, 
        n17592;
    wire [7:0]\data_out[2] ;   // coms.v(21[11:19])
    
    wire n17593, n5_adj_2141, n17495, n50, n48, n49, n5_adj_2142, 
        n9_adj_2143, n2338, n10379, n47_adj_2144, n30, n46, n45, 
        n17575, n1419, n2351, n2352, n18062, n26, n10696;
    wire [7:0]\data_out[8]_c ;   // coms.v(21[11:19])
    
    wire n17322, n17323, n18053, n2336, n9541, n20, n23, n10694, 
        n17347, n17346, n18056, n23_adj_2145, n56_adj_2146, n29_c, 
        n16533, n22, n9585, n27, n2334, n18, n51, n17266, n17268, 
        n2342, n26_adj_2147, n30_adj_2148, n9485, n10_adj_2149, n12_c, 
        n21, n15, n18014, n12_adj_2150, n16639, n17, n16148, n2340, 
        n17264;
    wire [7:0]\data_in_frame[1] ;   // coms.v(389[12:25])
    
    wire n17001, n16943, n9493, n16876, n17013, n6_adj_2152, n18047, 
        n9488, n17004, n18050, n17274, n9743, n8_adj_2153, n17638, 
        n10_adj_2154, n18020, n10_adj_2155, n16954, n15615, n16679, 
        n10369;
    wire [7:0]\data_in_frame[9] ;   // coms.v(389[12:25])
    
    wire n15938, n17014, n23_adj_2156, n17172, n8_adj_2157, n12_adj_2158, 
        n17262, n2_adj_2159, n3_c, n19, n16949, n17043, data_out_9__3__N_356, 
        n15939, n10368, n8_adj_2160, n10_adj_2162, n15518, n15519;
    wire [7:0]\data_out[3] ;   // coms.v(21[11:19])
    
    wire n10356, n44_adj_2163, n22_adj_2164, n42_adj_2165, n8_adj_2166, 
        n17574;
    wire [31:0]\FRAME_MATCHER.i_31__N_1280 ;
    
    wire n2_adj_2168, n8_adj_2169, n21_adj_2171, n2_adj_2172, n2_adj_2173, 
        n18_adj_2174, n2_adj_2175, n8_adj_2176, n17993, n17015, n16869, 
        n10859, n15525, n2_adj_2179, n2_adj_2180, n2_adj_2181, n2_adj_2182, 
        n28_adj_2183, n15929, n26_adj_2184, n10858, n17960, n17954, 
        n18125, n2_adj_2185, n2_adj_2186, n6_adj_2187, n17576, n18128, 
        n17569, n5_adj_2188, n18041, n12_adj_2189, n61, n59, n16133, 
        n17942, n17936, n18119, n2_adj_2190, n10_adj_2191, n2_adj_2192, 
        n17085, n17073, n17127, n14, n9688, n17128, n9692, n9810, 
        n16, n16923, n9819, n17031, n17_adj_2193, n17124, n17125, 
        n16926, n17022, n22_adj_2194, n2_adj_2195, n15930, n27_adj_2196, 
        n9913, n16_adj_2197, n24, n18_adj_2198, n25, n17256, n19_adj_2199, 
        n12_adj_2200, n6_adj_2201, n17578, n18122, n16772, n17079, 
        n20_adj_2202, n17115, n17126, n15526, n15846, tx2_transmit_N_1997, 
        n2_adj_2204, n12993, n13298, n9892, n20_adj_2205, n12991, 
        n2_adj_2206, n16247, n9859, n9555, n22_adj_2207, n17543, 
        n5_adj_2208, n18011, n2_adj_2209, n3_adj_2210, n2_adj_2211, 
        n2_adj_2212, n6_adj_2213, n5545, n17352, n2_adj_2214, n3_adj_2215, 
        n2_adj_2216, n3_adj_2217, n2_adj_2218, n3_adj_2219, n2_adj_2220, 
        n3_adj_2221, n2_adj_2222, n3_adj_2223, n2_adj_2224, n3_adj_2225, 
        n2_adj_2226, n3_adj_2227, n2_adj_2228, n3_adj_2229, n2_adj_2230, 
        n3_adj_2231, n2_adj_2232, n3_adj_2233, n2_adj_2234, n3_adj_2235, 
        n2_adj_2236, n3_adj_2237, n2_adj_2238, n3_adj_2239, n3_adj_2240, 
        n3_adj_2241, n3_adj_2242, n3_adj_2243, n3_adj_2244, n3_adj_2245, 
        n3_adj_2246, n3_adj_2247, n3_adj_2248, n3_adj_2249, n3_adj_2250, 
        n5543, n17354, n16946, n18_adj_2251, n17040, n17123, n17121, 
        n17924, n17918, n18107, n16871, n9678, n16940, n20_adj_2252, 
        n3_adj_2253;
    wire [14:0]n6517;
    
    wire n15524, n9901, n9754, n19_adj_2254, n16994, n17082, n17052, 
        n21_adj_2255, n18110, n17122, n16908, n3_adj_2256, n3_adj_2257, 
        n18101, n3_adj_2258, n3_adj_2259, n18104, n3_adj_2260;
    wire [0:0]n4130;
    wire [2:0]r_SM_Main_2__N_2036_adj_2400;
    
    wire n13496, n16898, n5_adj_2262, n16966, n9728, data_out_9__0__N_389, 
        n17393, n17894, n17963, n52, n9763, n17506;
    wire [0:0]n2502;
    
    wire data_out_6__1__N_537, n10259, n9853, n16960, n12_adj_2263, 
        n9886, n17053, n15517, n17103, n9919, n14_adj_2264, n17632, 
        n5_adj_2265, n18095, n2_adj_2266, n17581;
    wire [0:0]n2432;
    
    wire n20_adj_2267;
    wire [0:0]n2397;
    
    wire n9496, n9716, n10_adj_2268, data_out_9__1__N_378, n17507, 
        n16957, n15_adj_2269, n17046, n17097, n17105, n9758, n19_adj_2270, 
        n17514, n21_adj_2271, n24_adj_2272, n17049, n17091, n26_adj_2273, 
        n6_adj_2274, n16761, n17058, n16969, data_out_9__4__N_345, 
        n16987, n9814, n17010, n25_adj_2275, n17055, data_out_9__5__N_334, 
        n9530, n10_adj_2276, n18089, n17133, n27_adj_2277, n16981, 
        data_out_9__6__N_324, n6_adj_2278, n17561, n18092, n6_adj_2280, 
        n17571, n17966, n16972, n10_adj_2281, n17518, n17957, n17951, 
        n17637, n16912, n16978, n16975, n16998, n20_adj_2282, n7212, 
        n17522, n17061, n17104, n17945, n17948, n9522, n19_adj_2283, 
        n17939, n10363, n17528, n17933, n17007, n17028, n17094, 
        n21_adj_2284, n17927, data_out_9__7__N_272, n17930, data_out_7__2__N_447, 
        data_out_7__3__N_441, n17921, n9783, n17070, n9737, n17076, 
        n12_adj_2285, n17915, n17532, n17909, n17109, data_out_10__0__N_219, 
        n17912, n17534, n18008, n18083, n9707, n6_adj_2286, n10839, 
        n28_adj_2287, n9695, n10_adj_2288, n16918;
    wire [0:0]n2362;
    
    wire n16990, n17064, n12_adj_2289, n9916, data_out_10__1__N_168, 
        n6_adj_2290, n17563, n18086, n2_adj_2291, n17594, n9505, 
        n9839, n9589, n10_adj_2292, data_out_10__3__N_146, n17016, 
        n9671, n6_adj_2293, n9509, data_out_10__4__N_135, n9749, n28_adj_2294, 
        n32, n17025, data_out_10__5__N_124, n17034, n30_adj_2295, 
        n17067, n17100, n17118, n31_c, data_out_10__6__N_113;
    wire [7:0]tx_transmit_N_1949;
    
    wire n8938, n456, n29_adj_2296, n10618, n17135, n10464, n32_adj_2297, 
        data_out_10__7__N_101, n17589, n2_adj_2298, n10617;
    wire [0:0]n2292;
    
    wire n5_adj_2299, n8603, n17555, n5_adj_2300, n18035, n17548;
    wire [7:0]\data_in_frame[2] ;   // coms.v(389[12:25])
    
    wire n22_adj_2301, n10616, n10615, n10614, n10613, n10612, n10851, 
        n16915, n16933, n20_adj_2302, n10611, n19_adj_2303, n17106, 
        n21_adj_2304, n1_c, n17107, n17588;
    wire [0:0]n2327;
    
    wire n9826, n12_adj_2305, n11, n17236, n9865, n6_adj_2306, n17276, 
        n9843, n17987, n17990, n17278, n9910, n9579, n10_adj_2307, 
        n17112, n14_adj_2308, n23_adj_2309, n16839, n10380, n10381, 
        n17113, n17897, n10610, n8_adj_2310, n10384, n18029, n17445, 
        n4_adj_2311, n446, n10385, n17450, n13272, n16891, n10181, 
        n10382, n16_adj_2312, n15659, n15658, n15657, n10386, n15656, 
        n1439, n17037, n17088, n17_adj_2313, n17114, n15655, n15654;
    wire [31:0]\FRAME_MATCHER.i_31__N_1312 ;
    
    wire n17019, n26_adj_2314, n24_adj_2315, n25_adj_2316, n10387, 
        n8621, n5_adj_2317, n23_adj_2318, n17132, n15653, n10388, 
        n65, n17889, n15652, n16963, n15651, n9776, n15523, n15650, 
        n15649, data_out_10__2__N_157, n10609, n5_adj_2319, n15_adj_2320, 
        n10608, n5_adj_2321, n5_adj_2322, n14_adj_2323, n17131, n10604, 
        n10603, n10602, n10601, n10600, n15648, n16385, n16379, 
        n16387, n16381, n16389, n16353, n16391, n16355, n9895, 
        n16393, n16357, n16395, n16359, n16397, n16361, n16399, 
        n16363, n16401, n16365, n16403, n16367, n16405, n16369, 
        n16407, n16371, n16409, n16343, n16411, n16345, n16413, 
        n16347, n16415, n16349, n16417, n16351, n16419, n16447, 
        n16421, n16449, n16423, n16451, n16425, n16453, n16427, 
        n16455, n16429, n16445, n16431, n16443, n16433, n16441, 
        n16435, n16335, n16437, n16339, n16439, n16331;
    wire [0:0]n2257;
    
    wire n17254, n17460, n25_adj_2324, n6_adj_2325, n17456, n17547, 
        n5_adj_2326, n18023, n16_adj_2327, n17635, n17_adj_2328, n15647, 
        n17011, n10_adj_2329, n16895, n10389, n62, n13464, n10849, 
        n17591, n17590, n2_adj_2330, n10390, n15646, n16936, n15645, 
        n15644, n15643, n10846, n10391, n18005, n10467, n17351, 
        n10843, n18_adj_2331, n16_adj_2332, n20_adj_2333, n17108, 
        n17328, n17330, n17331, n15642, n5_adj_2334, n17333, n6_adj_2335, 
        n10383, n17560, n15522, n10_adj_2336, n17301, n17334, n17336;
    wire [7:0]\data_out_frame2[20] ;   // coms.v(390[12:27])
    
    wire n22_adj_2337, n17303, n16269, n16283, n16261, n16267, n16285, 
        n16281, n16257, n17345, n5_adj_2339, n16814, n20_adj_2340, 
        n23_adj_2341, n27_adj_2342, n18_adj_2343, n26_adj_2344, n30_adj_2345, 
        n17_adj_2346;
    wire [7:0]tx2_data;   // coms.v(412[13:21])
    
    wire n17337, n17769, n17339, n15516, n17639, n15641, n15521, 
        n17340, n17342, n9_adj_2347, n8_adj_2348, n17900, n5_adj_2349, 
        n5_adj_2350, n17546, n18017, n15640, n17343, n15515, n17290, 
        n17475, n17349, n5_adj_2351, n15639, n22_adj_2352, n22_adj_2353, 
        n17984, n22_adj_2354, n15638, n22_adj_2355, n15637, n15_adj_2356, 
        n15636, n22_adj_2357, n17981, n15520, n15635, n22_adj_2358, 
        n15634, n22_adj_2359, n15633, n15868, n8631, n9393, n17891, 
        n15632, n15514, n15631, n15630, n4_adj_2360, n15629, n15628, 
        n15627, n15527, n15626, n15625, n15624, n15623, n10376, 
        n15622, n15621, n15620;
    
    SB_DFF data_out_frame2_0___i109 (.Q(\data_out_frame2[13] [4]), .C(CLK_c), 
           .D(n10793));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i108 (.Q(\data_out_frame2[13] [3]), .C(CLK_c), 
           .D(n10792));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i107 (.Q(\data_out_frame2[13] [2]), .C(CLK_c), 
           .D(n10791));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i106 (.Q(\data_out_frame2[13] [1]), .C(CLK_c), 
           .D(n10790));   // coms.v(426[12] 547[6])
    SB_LUT4 i8017_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n10377));
    defparam i8017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame2_0___i105 (.Q(\data_out_frame2[13] [0]), .C(CLK_c), 
           .D(n10789));   // coms.v(426[12] 547[6])
    SB_DFF delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .D(n10470));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i104 (.Q(\data_out_frame2[12] [7]), .C(CLK_c), 
           .D(n10788));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i103 (.Q(\data_out_frame2[12] [6]), .C(CLK_c), 
           .D(n10787));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i102 (.Q(\data_out_frame2[12] [5]), .C(CLK_c), 
           .D(n10786));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i101 (.Q(\data_out_frame2[12] [4]), .C(CLK_c), 
           .D(n10785));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i100 (.Q(\data_out_frame2[12] [3]), .C(CLK_c), 
           .D(n10784));   // coms.v(426[12] 547[6])
    SB_LUT4 i15309_3_lut (.I0(\data_out_frame2[0] [1]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17579));
    defparam i15309_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 n17999_bdd_4_lut (.I0(n17999), .I1(\data_out_frame2[17] [6]), 
            .I2(\data_out_frame2[16] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18002));
    defparam n17999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut (.I0(n2), .I1(n12933), .I2(n127), .I3(n9435), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'hbaaa;
    SB_DFF data_out_frame2_0___i99 (.Q(\data_out_frame2[12] [2]), .C(CLK_c), 
           .D(n10783));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame2[6] [1]), 
            .I1(\data_out_frame2[7] [1]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_c));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut (.I0(n17454), .I1(n17452), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n9451), .O(n7));
    defparam i18_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state_c [31]), .I1(n4_c), .I2(GND_net), 
            .I3(GND_net), .O(n16377));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_403 (.I0(\FRAME_MATCHER.state_c [31]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16383));
    defparam i1_2_lut_adj_403.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out[8] [1]), .I2(\data_out[9] [1]), .I3(\byte_transmit_counter[3] ), 
            .O(n18077));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18077_bdd_4_lut (.I0(n18077), .I1(\data_out[1] [1]), .I2(\data_out[0][1] ), 
            .I3(\byte_transmit_counter[3] ), .O(n18080));
    defparam n18077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut (.I0(\data_out_frame2[5] [1]), 
            .I1(n5_c), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_c));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_out_frame2_0___i98 (.Q(\data_out_frame2[12] [1]), .C(CLK_c), 
           .D(n10782));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15621 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [7]), .I2(\data_out_frame2[11] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18071));
    defparam byte_transmit_counter2_0__bdd_4_lut_15621.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame2_0___i97 (.Q(\data_out_frame2[12] [0]), .C(CLK_c), 
           .D(n10781));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i96 (.Q(\data_out_frame2[11] [7]), .C(CLK_c), 
           .D(n10780));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_2353_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[4]), .I3(n15618), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame2_0___i95 (.Q(\data_out_frame2[11] [6]), .C(CLK_c), 
           .D(n10779));   // coms.v(426[12] 547[6])
    SB_LUT4 i10724_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n127_adj_2136), 
            .I2(n127), .I3(GND_net), .O(n1716));   // coms.v(440[13] 443[7])
    defparam i10724_3_lut.LUT_INIT = 16'hb3b3;
    SB_CARRY byte_transmit_counter2_2353_add_4_6 (.CI(n15618), .I0(GND_net), 
            .I1(byte_transmit_counter2[4]), .CO(n15619));
    SB_DFF \data_out_0[[1__2243  (.Q(\data_out[0][1] ), .C(CLK_c), .D(n10373));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i94 (.Q(\data_out_frame2[11] [5]), .C(CLK_c), 
           .D(n10778));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i93 (.Q(\data_out_frame2[11] [4]), .C(CLK_c), 
           .D(n10777));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i92 (.Q(\data_out_frame2[11] [3]), .C(CLK_c), 
           .D(n10776));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i91 (.Q(\data_out_frame2[11] [2]), .C(CLK_c), 
           .D(n10775));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i90 (.Q(\data_out_frame2[11] [1]), .C(CLK_c), 
           .D(n10774));   // coms.v(426[12] 547[6])
    SB_DFF delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .D(n10473));   // coms.v(280[12] 380[6])
    SB_LUT4 n17969_bdd_4_lut (.I0(n17969), .I1(\data_out_frame2[17] [4]), 
            .I2(\data_out_frame2[16] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n17972));
    defparam n17969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i89 (.Q(\data_out_frame2[11] [0]), .C(CLK_c), 
           .D(n10773));   // coms.v(426[12] 547[6])
    SB_DFF tx_active_prev_2155 (.Q(tx_active_prev), .C(CLK_c), .D(tx_active));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i88 (.Q(\data_out_frame2[10] [7]), .C(CLK_c), 
           .D(n10772));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i87 (.Q(\data_out_frame2[10] [6]), .C(CLK_c), 
           .D(n10771));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i86 (.Q(\data_out_frame2[10] [5]), .C(CLK_c), 
           .D(n10770));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_2353_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[3]), .I3(n15617), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame2_0___i85 (.Q(\data_out_frame2[10] [4]), .C(CLK_c), 
           .D(n10769));   // coms.v(426[12] 547[6])
    SB_DFFSR tx_transmit_2156 (.Q(r_SM_Main_2__N_2036[0]), .C(CLK_c), .D(n16838), 
            .R(n4445));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i84 (.Q(\data_out_frame2[10] [3]), .C(CLK_c), 
           .D(n10768));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i83 (.Q(\data_out_frame2[10] [2]), .C(CLK_c), 
           .D(n10767));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i82 (.Q(\data_out_frame2[10] [1]), .C(CLK_c), 
           .D(n10766));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i81 (.Q(\data_out_frame2[10] [0]), .C(CLK_c), 
           .D(n10765));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_7[[3__2185  (.Q(\data_out[7] [3]), .C(CLK_c), .E(n10054), 
            .D(n1846[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_7[[2__2186  (.Q(\data_out[7] [2]), .C(CLK_c), .E(n10054), 
            .D(n1881[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_7[[1__2187  (.Q(\data_out[7] [1]), .C(CLK_c), .E(n10054), 
            .D(n1916[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_7[[0__2188  (.Q(\data_out[7] [0]), .C(CLK_c), .E(n10054), 
            .D(n1951[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[7__2189  (.Q(\data_out[6] [7]), .C(CLK_c), .E(n10055), 
            .D(n1986[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[6__2190  (.Q(\data_out[6] [6]), .C(CLK_c), .E(n10055), 
            .D(n2021[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[5__2191  (.Q(\data_out[6] [5]), .C(CLK_c), .E(n10055), 
            .D(n2056[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[4__2192  (.Q(\data_out[6] [4]), .C(CLK_c), .E(n10055), 
            .D(n2091[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[3__2193  (.Q(\data_out[6] [3]), .C(CLK_c), .E(n10055), 
            .D(n2126[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[2__2194  (.Q(\data_out[6] [2]), .C(CLK_c), .E(n10055), 
            .D(n2161[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_6[[1__2195  (.Q(\data_out[6] [1]), .C(CLK_c), .E(n10055), 
            .D(n2196[0]));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_5[[1__2203  (.Q(\data_out[5] [1]), .C(CLK_c), .E(n10055), 
            .D(n2476[0]));   // coms.v(280[12] 380[6])
    SB_LUT4 n18071_bdd_4_lut (.I0(n18071), .I1(\data_out_frame2[9] [7]), 
            .I2(\data_out_frame2[8] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18074));
    defparam n18071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15355_2_lut (.I0(\data_out[1][7] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17585));
    defparam i15355_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFE \data_out_1[[1__2235  (.Q(\data_out[1] [1]), .C(CLK_c), .E(n10055), 
            .D(n3071[0]));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i80 (.Q(\data_out_frame2[9] [7]), .C(CLK_c), 
           .D(n10764));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i2_3_lut (.I0(\data_out[2][7] ), 
            .I1(\data_out[3][7] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2137));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \data_out_0[[3__2241  (.Q(\data_out[0][3] ), .C(CLK_c), .D(n10372));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i79 (.Q(\data_out_frame2[9] [6]), .C(CLK_c), 
           .D(n10763));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_0[[5__2239  (.Q(\data_out[0][5] ), .C(CLK_c), .D(n10371));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i78 (.Q(\data_out_frame2[9] [5]), .C(CLK_c), 
           .D(n10762));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_0[[6__2238  (.Q(\data_out[0] [6]), .C(CLK_c), .D(n10370));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i77 (.Q(\data_out_frame2[9] [4]), .C(CLK_c), 
           .D(n10761));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i76 (.Q(\data_out_frame2[9] [3]), .C(CLK_c), 
           .D(n10760));   // coms.v(426[12] 547[6])
    SB_LUT4 i10695_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n9346), .I3(\FRAME_MATCHER.i [1]), .O(n2275));   // coms.v(453[9:60])
    defparam i10695_4_lut.LUT_INIT = 16'h3230;
    SB_DFF data_out_frame2_0___i75 (.Q(\data_out_frame2[9] [2]), .C(CLK_c), 
           .D(n10759));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i74 (.Q(\data_out_frame2[9] [1]), .C(CLK_c), 
           .D(n10758));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i152 (.Q(\data_out_frame2[18] [7]), .C(CLK_c), 
           .D(n10836));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i151 (.Q(\data_out_frame2[18] [6]), .C(CLK_c), 
           .D(n10835));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i150 (.Q(\data_out_frame2[18] [5]), .C(CLK_c), 
           .D(n10834));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i149 (.Q(\data_out_frame2[18] [4]), .C(CLK_c), 
           .D(n10833));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i148 (.Q(\data_out_frame2[18] [3]), .C(CLK_c), 
           .D(n10832));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i73 (.Q(\data_out_frame2[9] [0]), .C(CLK_c), 
           .D(n10757));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i132 (.Q(\data_out_frame2[16] [3]), .C(CLK_c), 
           .D(n10816));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i72 (.Q(\data_out_frame2[8] [7]), .C(CLK_c), 
           .D(n10756));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i131 (.Q(\data_out_frame2[16] [2]), .C(CLK_c), 
           .D(n10815));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i71 (.Q(\data_out_frame2[8] [6]), .C(CLK_c), 
           .D(n10755));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i130 (.Q(\data_out_frame2[16] [1]), .C(CLK_c), 
           .D(n10814));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i70 (.Q(\data_out_frame2[8] [5]), .C(CLK_c), 
           .D(n10754));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i129 (.Q(\data_out_frame2[16] [0]), .C(CLK_c), 
           .D(n10813));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i69 (.Q(\data_out_frame2[8] [4]), .C(CLK_c), 
           .D(n10753));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i128 (.Q(\data_out_frame2[15] [7]), .C(CLK_c), 
           .D(n10812));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i127 (.Q(\data_out_frame2[15] [6]), .C(CLK_c), 
           .D(n10811));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i126 (.Q(\data_out_frame2[15] [5]), .C(CLK_c), 
           .D(n10810));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i125 (.Q(\data_out_frame2[15] [4]), .C(CLK_c), 
           .D(n10809));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i124 (.Q(\data_out_frame2[15] [3]), .C(CLK_c), 
           .D(n10808));   // coms.v(426[12] 547[6])
    SB_DFF delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .D(n10867));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .D(n10479));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .D(n10865));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .D(n10485));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .D(n10488));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .D(n10491));   // coms.v(280[12] 380[6])
    SB_DFF delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .D(n10494));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i123 (.Q(\data_out_frame2[15] [2]), .C(CLK_c), 
           .D(n10807));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i122 (.Q(\data_out_frame2[15] [1]), .C(CLK_c), 
           .D(n10806));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i121 (.Q(\data_out_frame2[15] [0]), .C(CLK_c), 
           .D(n10805));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i120 (.Q(\data_out_frame2[14] [7]), .C(CLK_c), 
           .D(n10804));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i119 (.Q(\data_out_frame2[14] [6]), .C(CLK_c), 
           .D(n10803));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i118 (.Q(\data_out_frame2[14] [5]), .C(CLK_c), 
           .D(n10802));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i68 (.Q(\data_out_frame2[8] [3]), .C(CLK_c), 
           .D(n10752));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i117 (.Q(\data_out_frame2[14] [4]), .C(CLK_c), 
           .D(n10801));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i67 (.Q(\data_out_frame2[8] [2]), .C(CLK_c), 
           .D(n10751));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i116 (.Q(\data_out_frame2[14] [3]), .C(CLK_c), 
           .D(n10800));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i66 (.Q(\data_out_frame2[8] [1]), .C(CLK_c), 
           .D(n10750));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i115 (.Q(\data_out_frame2[14] [2]), .C(CLK_c), 
           .D(n10799));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i65 (.Q(\data_out_frame2[8] [0]), .C(CLK_c), 
           .D(n10749));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i114 (.Q(\data_out_frame2[14] [1]), .C(CLK_c), 
           .D(n10798));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i64 (.Q(\data_out_frame2[7] [7]), .C(CLK_c), 
           .D(n10748));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i113 (.Q(\data_out_frame2[14] [0]), .C(CLK_c), 
           .D(n10797));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i63 (.Q(\data_out_frame2[7] [6]), .C(CLK_c), 
           .D(n10747));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i112 (.Q(\data_out_frame2[13] [7]), .C(CLK_c), 
           .D(n10796));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i62 (.Q(\data_out_frame2[7] [5]), .C(CLK_c), 
           .D(n10746));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i61 (.Q(\data_out_frame2[7] [4]), .C(CLK_c), 
           .D(n10745));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i8_3_lut (.I0(\data_out[8] [0]), 
            .I1(\data_out[9] [0]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2138));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i10_4_lut (.I0(n8_adj_2138), 
            .I1(\data_out[10] [0]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_c));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i24_4_lut (.I0(n18098), .I1(n10_c), .I2(\byte_transmit_counter[3] ), 
            .I3(\byte_transmit_counter[2] ), .O(n10_adj_2139));   // coms.v(19[11:32])
    defparam i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i23_4_lut (.I0(r_Tx_Data[0]), .I1(n10_adj_2139), .I2(n8730), 
            .I3(\byte_transmit_counter[4] ), .O(n16595));   // coms.v(19[11:32])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_out_frame2_0___i60 (.Q(\data_out_frame2[7] [3]), .C(CLK_c), 
           .D(n10744));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i59 (.Q(\data_out_frame2[7] [2]), .C(CLK_c), 
           .D(n10743));   // coms.v(426[12] 547[6])
    SB_DFF delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .D(n10860));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i58 (.Q(\data_out_frame2[7] [1]), .C(CLK_c), 
           .D(n10742));   // coms.v(426[12] 547[6])
    SB_LUT4 i14820_4_lut (.I0(n47), .I1(n56), .I2(n60), .I3(n33_c), 
            .O(n17258));
    defparam i14820_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33_3_lut (.I0(n9451), .I1(n9460), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n28));
    defparam i33_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(\FRAME_MATCHER.state_c [24]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n9));
    defparam i3_3_lut.LUT_INIT = 16'h5454;
    SB_DFF data_out_frame2_0___i57 (.Q(\data_out_frame2[7] [0]), .C(CLK_c), 
           .D(n10741));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_4_lut_adj_404 (.I0(n12933), .I1(n9), .I2(n28), .I3(n17258), 
            .O(n16795));
    defparam i1_4_lut_adj_404.LUT_INIT = 16'h5fdf;
    SB_DFF data_out_frame2_0___i56 (.Q(\data_out_frame2[6] [7]), .C(CLK_c), 
           .D(n10740));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15597 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [7]), .I2(\data_out_frame2[15] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18065));
    defparam byte_transmit_counter2_0__bdd_4_lut_15597.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame2_0___i55 (.Q(\data_out_frame2[6] [6]), .C(CLK_c), 
           .D(n10739));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i54 (.Q(\data_out_frame2[6] [5]), .C(CLK_c), 
           .D(n10738));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i53 (.Q(\data_out_frame2[6] [4]), .C(CLK_c), 
           .D(n10737));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i52 (.Q(\data_out_frame2[6] [3]), .C(CLK_c), 
           .D(n10736));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i51 (.Q(\data_out_frame2[6] [2]), .C(CLK_c), 
           .D(n10735));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i50 (.Q(\data_out_frame2[6] [1]), .C(CLK_c), 
           .D(n10734));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i49 (.Q(\data_out_frame2[6] [0]), .C(CLK_c), 
           .D(n10733));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i48 (.Q(\data_out_frame2[5] [7]), .C(CLK_c), 
           .D(n10732));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i47 (.Q(\data_out_frame2[5] [6]), .C(CLK_c), 
           .D(n10731));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i46 (.Q(\data_out_frame2[5] [5]), .C(CLK_c), 
           .D(n10730));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i45 (.Q(\data_out_frame2[5] [4]), .C(CLK_c), 
           .D(n10729));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i44 (.Q(\data_out_frame2[5] [3]), .C(CLK_c), 
           .D(n10728));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i43 (.Q(\data_out_frame2[5] [2]), .C(CLK_c), 
           .D(n10727));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i42 (.Q(\data_out_frame2[5] [1]), .C(CLK_c), 
           .D(n10726));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i41 (.Q(\data_out_frame2[5] [0]), .C(CLK_c), 
           .D(n10725));   // coms.v(426[12] 547[6])
    SB_DFF \UART_TRANSMITTER.state_i0_i1  (.Q(\UART_TRANSMITTER.state[1] ), 
           .C(CLK_c), .D(n16255));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_405 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2140));   // coms.v(448[5:27])
    defparam i1_2_lut_adj_405.LUT_INIT = 16'heeee;
    SB_LUT4 i8018_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n10378));
    defparam i8018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY byte_transmit_counter2_2353_add_4_5 (.CI(n15617), .I0(GND_net), 
            .I1(byte_transmit_counter2[3]), .CO(n15618));
    SB_LUT4 n18065_bdd_4_lut (.I0(n18065), .I1(\data_out_frame2[13] [7]), 
            .I2(\data_out_frame2[12] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18068));
    defparam n18065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut (.I0(\FRAME_MATCHER.state_c [4]), .I1(n16905), .I2(n16879), 
            .I3(n6_adj_2140), .O(n9451));   // coms.v(448[5:27])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15592 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [7]), .I2(\data_out_frame2[19] [7]), 
            .I3(byte_transmit_counter2[1]), .O(n18059));
    defparam byte_transmit_counter2_0__bdd_4_lut_15592.LUT_INIT = 16'he4aa;
    SB_LUT4 i14802_2_lut (.I0(\data_in[1] [2]), .I1(\data_in[3] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n17240));
    defparam i14802_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4030_2_lut (.I0(\UART_TRANSMITTER.state[0] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n2546[0]));   // coms.v(283[4] 379[11])
    defparam i4030_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(\data_in[1] [1]), .I1(n9490), .I2(n9482), .I3(n17240), 
            .O(n127));
    defparam i3_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i10728_2_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n127), .I2(GND_net), 
            .I3(GND_net), .O(n1651));   // coms.v(440[13] 443[7])
    defparam i10728_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_406 (.I0(\FRAME_MATCHER.state [2]), .I1(n9451), 
            .I2(GND_net), .I3(GND_net), .O(n9453));   // coms.v(502[5:21])
    defparam i1_2_lut_adj_406.LUT_INIT = 16'hdddd;
    SB_LUT4 i15423_4_lut (.I0(n4445), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n10055));
    defparam i15423_4_lut.LUT_INIT = 16'h4444;
    SB_LUT4 byte_transmit_counter2_2353_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[2]), .I3(n15616), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR byte_transmit_counter2_2353__i1 (.Q(byte_transmit_counter2[1]), 
            .C(CLK_c), .E(n10052), .D(n37[1]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [16]), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(GND_net), .O(n16905));   // coms.v(448[5:27])
    defparam i1_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFFESR byte_transmit_counter2_2353__i2 (.Q(byte_transmit_counter2[2]), 
            .C(CLK_c), .E(n10052), .D(n37[2]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_DFFESR byte_transmit_counter2_2353__i3 (.Q(byte_transmit_counter2[3]), 
            .C(CLK_c), .E(n10052), .D(n37[3]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_DFFESR byte_transmit_counter2_2353__i4 (.Q(byte_transmit_counter2[4]), 
            .C(CLK_c), .E(n10052), .D(n37[4]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_DFFESR byte_transmit_counter2_2353__i5 (.Q(byte_transmit_counter2[5]), 
            .C(CLK_c), .E(n10052), .D(n37[5]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_DFFESR byte_transmit_counter2_2353__i6 (.Q(byte_transmit_counter2[6]), 
            .C(CLK_c), .E(n10052), .D(n37[6]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_DFFESR byte_transmit_counter2_2353__i7 (.Q(byte_transmit_counter2[7]), 
            .C(CLK_c), .E(n10052), .D(n37[7]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_LUT4 i15344_2_lut (.I0(\data_out[0][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17592));
    defparam i15344_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15290_2_lut (.I0(\data_out[2] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17593));
    defparam i15290_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame2[6] [4]), 
            .I1(\data_out_frame2[7] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2141));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15368_2_lut (.I0(\data_out_frame2[5] [4]), .I1(byte_transmit_counter2[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17495));
    defparam i15368_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [6]), .I3(\FRAME_MATCHER.i [9]), .O(n50));   // coms.v(450[7:23])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [15]), .O(n48));   // coms.v(450[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [23]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n49));   // coms.v(450[7:23])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out[6] [1]), 
            .I1(\data_out[7] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2142));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10915_2_lut (.I0(\data_out[10] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_2143));   // coms.v(257[28:49])
    defparam i10915_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1032_2_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n2338));   // coms.v(67[15:26])
    defparam i1032_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8019_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n10379));
    defparam i8019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_407 (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i [30]), 
            .I2(\FRAME_MATCHER.i [27]), .I3(\FRAME_MATCHER.i [8]), .O(n47_adj_2144));   // coms.v(450[7:23])
    defparam i18_4_lut_adj_407.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_408 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(GND_net), .I3(GND_net), .O(n30));   // coms.v(450[7:23])
    defparam i1_2_lut_adj_408.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [24]), .O(n46));   // coms.v(450[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [12]), .O(n45));   // coms.v(450[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9279_3_lut (.I0(delay_counter[12]), .I1(n17575), .I2(n1419), 
            .I3(GND_net), .O(n10860));
    defparam i9279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1046_2_lut (.I0(n2351), .I1(\data_in_frame[0] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n2352));   // coms.v(76[16:69])
    defparam i1046_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n18059_bdd_4_lut (.I0(n18059), .I1(\data_out_frame2[17] [7]), 
            .I2(\data_out_frame2[16] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n18062));
    defparam n18059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \data_out_6[[0__2196  (.Q(\data_out[6][0] ), .C(CLK_c), .E(VCC_net), 
            .D(n16607));   // coms.v(280[12] 380[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state[1] ), .C(CLK_c), 
           .D(n18137));   // coms.v(426[12] 547[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n16797));   // coms.v(426[12] 547[6])
    SB_LUT4 i53_4_lut (.I0(\data_out[5] [1]), .I1(n5_adj_2142), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n26));   // coms.v(19[11:32])
    defparam i53_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF \data_out_8[[0__2180  (.Q(\data_out[8] [0]), .C(CLK_c), .D(n10698));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_8[[1__2179  (.Q(\data_out[8] [1]), .C(CLK_c), .D(n10697));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_8[[2__2178  (.Q(\data_out[8]_c [2]), .C(CLK_c), .D(n10696));   // coms.v(280[12] 380[6])
    SB_LUT4 byte_transmit_counter2_1__bdd_4_lut (.I0(byte_transmit_counter2[1]), 
            .I1(n17322), .I2(n17323), .I3(byte_transmit_counter2[2]), 
            .O(n18053));
    defparam byte_transmit_counter2_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_409 (.I0(\data_in_frame[7] [3]), .I1(n2336), .I2(n9541), 
            .I3(\data_in_frame[7] [5]), .O(n20));
    defparam i4_4_lut_adj_409.LUT_INIT = 16'h7bde;
    SB_LUT4 i50_4_lut (.I0(n18080), .I1(n9_adj_2143), .I2(byte_transmit_counter[1]), 
            .I3(\byte_transmit_counter[3] ), .O(n23));   // coms.v(19[11:32])
    defparam i50_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF \data_in_3[[7__2250  (.Q(\data_in[3] [7]), .C(CLK_c), .D(n10695));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_8[[3__2177  (.Q(\data_out[8]_c [3]), .C(CLK_c), .D(n10694));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_8[[4__2176  (.Q(\data_out[8][4] ), .C(CLK_c), .D(n10693));   // coms.v(280[12] 380[6])
    SB_LUT4 n18053_bdd_4_lut (.I0(n18053), .I1(n17347), .I2(n17346), .I3(byte_transmit_counter2[2]), 
            .O(n18056));
    defparam n18053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[0] [7]), .I1(n2352), .I2(\data_in_frame[6] [1]), 
            .I3(\data_in_frame[6] [7]), .O(n23_adj_2145));
    defparam i7_4_lut.LUT_INIT = 16'hde7b;
    SB_LUT4 i27_4_lut (.I0(n47_adj_2144), .I1(n49), .I2(n48), .I3(n50), 
            .O(n56_adj_2146));   // coms.v(450[7:23])
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52_4_lut (.I0(n23), .I1(\byte_transmit_counter[3] ), .I2(\byte_transmit_counter[2] ), 
            .I3(n26), .O(n29_c));   // coms.v(19[11:32])
    defparam i52_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i51_4_lut (.I0(r_Tx_Data[1]), .I1(n29_c), .I2(n8730), .I3(\byte_transmit_counter[4] ), 
            .O(n16533));   // coms.v(19[11:32])
    defparam i51_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[6] [2]), .I1(n22), .I2(\data_in_frame[7] [2]), 
            .I3(n9585), .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hdffd;
    SB_LUT4 i2_4_lut (.I0(n2351), .I1(n2334), .I2(\data_in_frame[7] [1]), 
            .I3(\data_in_frame[7] [4]), .O(n18));
    defparam i2_4_lut.LUT_INIT = 16'hb7ed;
    SB_LUT4 i22_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n30), .O(n51));   // coms.v(450[7:23])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28_4_lut (.I0(n51), .I1(n56_adj_2146), .I2(n45), .I3(n46), 
            .O(n9346));   // coms.v(450[7:23])
    defparam i28_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14828_4_lut (.I0(\data_in[2] [7]), .I1(\data_in[2] [2]), .I2(\data_in[0] [1]), 
            .I3(\data_in[2] [5]), .O(n17266));
    defparam i14828_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i14830_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[0] [3]), .I2(\data_in[2] [0]), 
            .I3(GND_net), .O(n17268));
    defparam i14830_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10_4_lut (.I0(n2342), .I1(n20), .I2(\data_in_frame[6] [5]), 
            .I3(\data_in_frame[6] [0]), .O(n26_adj_2147));
    defparam i10_4_lut.LUT_INIT = 16'hefdf;
    SB_LUT4 i14_4_lut (.I0(n27), .I1(n23_adj_2145), .I2(\data_in_frame[6] [3]), 
            .I3(\data_in_frame[6] [4]), .O(n30_adj_2148));
    defparam i14_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i4_4_lut_adj_410 (.I0(\data_in[0] [0]), .I1(\data_in[1] [6]), 
            .I2(n9485), .I3(\data_in[3] [5]), .O(n10_adj_2149));
    defparam i4_4_lut_adj_410.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(\data_in[3] [7]), .I1(n10_adj_2149), .I2(n17268), 
            .I3(n17266), .O(n9482));
    defparam i5_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i10680_2_lut (.I0(n9346), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n3977));   // coms.v(507[9:40])
    defparam i10680_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_411 (.I0(\data_in[3] [0]), .I1(\data_in[3] [4]), 
            .I2(\data_in[0] [5]), .I3(n9482), .O(n12_c));
    defparam i5_4_lut_adj_411.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_3_lut (.I0(\data_out[8]_c [2]), .I1(\data_out[9][2] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n21));   // coms.v(19[11:32])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30_4_lut (.I0(n21), .I1(\data_out[10] [2]), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n15));
    defparam i30_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31_4_lut (.I0(n18014), .I1(n15), .I2(\byte_transmit_counter[3] ), 
            .I3(\byte_transmit_counter[2] ), .O(n12_adj_2150));
    defparam i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29_4_lut (.I0(r_Tx_Data[2]), .I1(n12_adj_2150), .I2(n8730), 
            .I3(\byte_transmit_counter[4] ), .O(n16639));
    defparam i29_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_412 (.I0(n2352), .I1(n2338), .I2(\data_in_frame[7] [0]), 
            .I3(\data_in_frame[7] [6]), .O(n17));
    defparam i1_4_lut_adj_412.LUT_INIT = 16'h7bde;
    SB_LUT4 i15_4_lut (.I0(n17), .I1(n30_adj_2148), .I2(n26_adj_2147), 
            .I3(n18), .O(n16148));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1034_2_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n2340));   // coms.v(68[15:26])
    defparam i1034_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14826_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[0] [6]), .I2(\data_in[1] [4]), 
            .I3(GND_net), .O(n17264));
    defparam i14826_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_413 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17001));   // coms.v(513[9:61])
    defparam i1_2_lut_adj_413.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_414 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(n9541), .O(n16943));   // coms.v(76[16:62])
    defparam i3_4_lut_adj_414.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n17264), .I1(n12_c), .I2(n9493), .I3(\data_in[3] [2]), 
            .O(n127_adj_4));
    defparam i6_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1030_2_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n2336));   // coms.v(66[15:26])
    defparam i1030_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_415 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n16876), 
            .I2(GND_net), .I3(GND_net), .O(n60));   // coms.v(457[5:29])
    defparam i1_2_lut_adj_415.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_416 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n9541));   // coms.v(76[16:62])
    defparam i1_2_lut_adj_416.LUT_INIT = 16'h6666;
    SB_LUT4 i1028_2_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n2334));   // coms.v(65[15:26])
    defparam i1028_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1036_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2342));   // coms.v(69[15:26])
    defparam i1036_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(n56), .I1(\FRAME_MATCHER.state_c [24]), .I2(n60), 
            .I3(GND_net), .O(n16879));   // coms.v(457[5:29])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut (.I0(\FRAME_MATCHER.state_c [8]), .I1(\FRAME_MATCHER.state_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_c));   // coms.v(457[5:29])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF \data_out_8[[5__2175  (.Q(\data_out[8][5] ), .C(CLK_c), .D(n10692));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_417 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9585));   // coms.v(117[16:35])
    defparam i1_2_lut_adj_417.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_418 (.I0(\FRAME_MATCHER.state_c [16]), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n47));   // coms.v(457[5:29])
    defparam i2_3_lut_adj_418.LUT_INIT = 16'hfefe;
    SB_DFF \data_out_8[[6__2174  (.Q(\data_out[8][6] ), .C(CLK_c), .D(n10691));   // coms.v(280[12] 380[6])
    SB_LUT4 i3_4_lut_adj_419 (.I0(n47), .I1(\FRAME_MATCHER.state [2]), .I2(n33_c), 
            .I3(n16879), .O(n9445));   // coms.v(457[5:29])
    defparam i3_4_lut_adj_419.LUT_INIT = 16'hfffe;
    SB_DFF \data_out_8[[7__2173  (.Q(\data_out[8][7] ), .C(CLK_c), .D(n10690));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i147 (.Q(\data_out_frame2[18] [2]), .C(CLK_c), 
           .D(n10831));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_420 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17013));   // coms.v(130[17:124])
    defparam i1_2_lut_adj_420.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_421 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n6_adj_2152));   // coms.v(513[9:61])
    defparam i1_3_lut_adj_421.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame2_0___i146 (.Q(\data_out_frame2[18] [1]), .C(CLK_c), 
           .D(n10830));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15587 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [6]), .I2(\data_out_frame2[11] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18047));
    defparam byte_transmit_counter2_0__bdd_4_lut_15587.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_422 (.I0(\FRAME_MATCHER.state[1] ), .I1(n9445), 
            .I2(GND_net), .I3(GND_net), .O(n9488));   // coms.v(434[90:101])
    defparam i1_2_lut_adj_422.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_423 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17004));   // coms.v(513[9:61])
    defparam i1_2_lut_adj_423.LUT_INIT = 16'h6666;
    SB_LUT4 n18047_bdd_4_lut (.I0(n18047), .I1(\data_out_frame2[9] [6]), 
            .I2(\data_out_frame2[8] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18050));
    defparam n18047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame2_0___i145 (.Q(\data_out_frame2[18] [0]), .C(CLK_c), 
           .D(n10829));   // coms.v(426[12] 547[6])
    SB_LUT4 i14836_4_lut (.I0(\data_in[0] [5]), .I1(\data_in[3] [0]), .I2(\data_in[3] [4]), 
            .I3(\data_in[3] [2]), .O(n17274));
    defparam i14836_4_lut.LUT_INIT = 16'h8000;
    SB_DFF \data_in_3[[5__2252  (.Q(\data_in[3] [5]), .C(CLK_c), .D(n10689));   // coms.v(426[12] 547[6])
    SB_LUT4 i3_4_lut_adj_424 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(\data_in[2] [3]), .I3(n17274), .O(n9490));
    defparam i3_4_lut_adj_424.LUT_INIT = 16'hfeff;
    SB_DFF data_out_frame2_0___i144 (.Q(\data_out_frame2[17] [7]), .C(CLK_c), 
           .D(n10828));   // coms.v(426[12] 547[6])
    SB_LUT4 i4_4_lut_adj_425 (.I0(n16943), .I1(n17004), .I2(n17001), .I3(n6_adj_2152), 
            .O(n9743));   // coms.v(513[9:61])
    defparam i4_4_lut_adj_425.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i8_3_lut (.I0(\data_out[8]_c [3]), 
            .I1(\data_out[9] [3]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2153));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12741_3_lut (.I0(delay_counter[7]), .I1(n17638), .I2(n1419), 
            .I3(GND_net), .O(n10865));
    defparam i12741_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY byte_transmit_counter2_2353_add_4_4 (.CI(n15616), .I0(GND_net), 
            .I1(byte_transmit_counter2[2]), .CO(n15617));
    SB_DFF \data_in_3[[6__2251  (.Q(\data_in[3] [6]), .C(CLK_c), .D(n10688));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i10_4_lut (.I0(n8_adj_2153), 
            .I1(\data_out[10] [3]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_2154));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i24_4_lut_adj_426 (.I0(n18020), .I1(n10_adj_2154), .I2(\byte_transmit_counter[3] ), 
            .I3(\byte_transmit_counter[2] ), .O(n10_adj_2155));
    defparam i24_4_lut_adj_426.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_4_lut_adj_427 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [6]), 
            .I2(n9743), .I3(\data_in_frame[10] [1]), .O(n16954));   // coms.v(130[17:124])
    defparam i2_4_lut_adj_427.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_2353_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[1]), .I3(n15615), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF \data_out_9[[2__2170  (.Q(\data_out[9][2] ), .C(CLK_c), .D(n10687));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_3[[4__2253  (.Q(\data_in[3] [4]), .C(CLK_c), .D(n10686));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_3[[3__2254  (.Q(\data_in[3] [3]), .C(CLK_c), .D(n10685));   // coms.v(426[12] 547[6])
    SB_LUT4 i23_4_lut_adj_428 (.I0(r_Tx_Data[3]), .I1(n10_adj_2155), .I2(n8730), 
            .I3(\byte_transmit_counter[4] ), .O(n16679));
    defparam i23_4_lut_adj_428.LUT_INIT = 16'h0aca;
    SB_DFF \data_out_1[[2__2234  (.Q(\data_out[1] [2]), .C(CLK_c), .D(n10369));   // coms.v(280[12] 380[6])
    SB_LUT4 i2_3_lut_adj_429 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n15938));   // coms.v(513[9:61])
    defparam i2_3_lut_adj_429.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_430 (.I0(\data_in_frame[1] [6]), .I1(n9743), .I2(\data_in_frame[9] [7]), 
            .I3(n17013), .O(n17014));   // coms.v(130[17:124])
    defparam i3_4_lut_adj_430.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_431 (.I0(\data_in_frame[9] [3]), .I1(n15938), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[1] [2]), .O(n23_adj_2156));   // coms.v(513[9:61])
    defparam i7_4_lut_adj_431.LUT_INIT = 16'hedde;
    SB_LUT4 i14734_2_lut (.I0(\data_in[1] [3]), .I1(\data_in[1] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n17172));
    defparam i14734_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_432 (.I0(\data_in[2] [6]), .I1(\data_in[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_2157));   // coms.v(437[16:89])
    defparam i1_2_lut_adj_432.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_433 (.I0(\data_in[2] [4]), .I1(\data_in[0] [2]), 
            .I2(\data_in[3] [1]), .I3(\data_in[2] [1]), .O(n12_adj_2158));   // coms.v(437[16:89])
    defparam i5_4_lut_adj_433.LUT_INIT = 16'hfffe;
    SB_LUT4 i14824_4_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [5]), .I2(\data_in[0] [4]), 
            .I3(n17172), .O(n17262));
    defparam i14824_4_lut.LUT_INIT = 16'h8000;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2_adj_2159), .S(n3_c));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_3[[2__2255  (.Q(\data_in[3] [2]), .C(CLK_c), .D(n10684));   // coms.v(426[12] 547[6])
    SB_LUT4 i3_4_lut_adj_434 (.I0(n2342), .I1(\data_in_frame[9] [5]), .I2(\data_in_frame[9] [0]), 
            .I3(n17004), .O(n19));   // coms.v(513[9:61])
    defparam i3_4_lut_adj_434.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out[5] [1]), .I1(\data_out[8][7] ), 
            .I2(n16949), .I3(n17043), .O(data_out_9__3__N_356));   // coms.v(181[17:93])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF \data_in_3[[1__2256  (.Q(\data_in[3] [1]), .C(CLK_c), .D(n10683));   // coms.v(426[12] 547[6])
    SB_LUT4 i2_3_lut_adj_435 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n15939));   // coms.v(513[9:61])
    defparam i2_3_lut_adj_435.LUT_INIT = 16'h9696;
    SB_DFF \data_in_3[[0__2257  (.Q(\data_in[3] [0]), .C(CLK_c), .D(n10682));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_2[[7__2258  (.Q(\data_in[2] [7]), .C(CLK_c), .D(n10681));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_2[[6__2259  (.Q(\data_in[2] [6]), .C(CLK_c), .D(n10680));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_2[[5__2260  (.Q(\data_in[2] [5]), .C(CLK_c), .D(n10679));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_2[[4__2261  (.Q(\data_in[2] [4]), .C(CLK_c), .D(n10678));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_2[[3__2262  (.Q(\data_in[2] [3]), .C(CLK_c), .D(n10677));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_1[[4__2232  (.Q(\data_out[1] [4]), .C(CLK_c), .D(n10368));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_2[[2__2263  (.Q(\data_in[2] [2]), .C(CLK_c), .D(n10676));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i143 (.Q(\data_out_frame2[17] [6]), .C(CLK_c), 
           .D(n10827));   // coms.v(426[12] 547[6])
    SB_CARRY byte_transmit_counter2_2353_add_4_3 (.CI(n15615), .I0(GND_net), 
            .I1(byte_transmit_counter2[1]), .CO(n15616));
    SB_LUT4 i1_4_lut_adj_436 (.I0(n17262), .I1(n9488), .I2(n12_adj_2158), 
            .I3(n8_adj_2157), .O(n9485));   // coms.v(437[16:89])
    defparam i1_4_lut_adj_436.LUT_INIT = 16'hfffd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i8_3_lut (.I0(\data_out[8][4] ), 
            .I1(\data_out[9] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2160));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i10_4_lut (.I0(n8_adj_2160), 
            .I1(\data_out[10] [4]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF \data_in_2[[1__2264  (.Q(\data_in[2] [1]), .C(CLK_c), .D(n10675));   // coms.v(426[12] 547[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out[5] [1]), .I1(\data_out[8][7] ), 
            .I2(\data_out[10] [6]), .I3(n10_adj_2162), .O(data_out_9__2__N_367));   // coms.v(181[17:93])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2495_7 (.CI(n15518), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n15519));
    SB_LUT4 i7996_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10055), .I3(\data_out[3] [6]), .O(n10356));   // coms.v(283[4] 379[11])
    defparam i7996_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_4_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n44_adj_2163), .I3(n22_adj_2164), .O(n42_adj_2165));   // coms.v(283[4] 379[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'he2c0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i8_3_lut (.I0(\data_out[8][5] ), 
            .I1(\data_out[9] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2166));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9277_3_lut (.I0(delay_counter[5]), .I1(n17574), .I2(n1419), 
            .I3(GND_net), .O(n10867));
    defparam i9277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_437 (.I0(\data_in[1] [2]), .I1(\data_in[1] [1]), 
            .I2(\data_in[3] [6]), .I3(GND_net), .O(n9493));   // coms.v(434[7:86])
    defparam i2_3_lut_adj_437.LUT_INIT = 16'hfbfb;
    SB_DFF \data_in_2[[0__2265  (.Q(\data_in[2] [0]), .C(CLK_c), .D(n10674));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i142 (.Q(\data_out_frame2[17] [5]), .C(CLK_c), 
           .D(n10826));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i10_4_lut (.I0(n8_adj_2166), 
            .I1(\data_out[10] [5]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_5));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8009_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10055), .I3(\data_out[1] [2]), .O(n10369));   // coms.v(283[4] 379[11])
    defparam i8009_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(n16886), .O(n9361));   // coms.v(283[4] 379[11])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 select_238_Select_1_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [1]), .I3(GND_net), .O(n2_adj_2168));
    defparam select_238_Select_1_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i8_3_lut (.I0(\data_out[8][6] ), 
            .I1(\data_out[9] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2169));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i10_4_lut (.I0(n8_adj_2169), 
            .I1(\data_out[10] [6]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_6));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_4_lut_adj_438 (.I0(\data_in_frame[9] [2]), .I1(n15939), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[1] [1]), .O(n21_adj_2171));   // coms.v(513[9:61])
    defparam i5_4_lut_adj_438.LUT_INIT = 16'hedde;
    SB_LUT4 select_238_Select_2_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [2]), .I3(GND_net), .O(n2_adj_2172));
    defparam select_238_Select_2_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_in_1[[7__2266  (.Q(\data_in[1] [7]), .C(CLK_c), .D(n10673));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_3_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [3]), .I3(GND_net), .O(n2_adj_2173));
    defparam select_238_Select_3_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i2_3_lut_adj_439 (.I0(n16954), .I1(n2334), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n18_adj_2174));   // coms.v(513[9:61])
    defparam i2_3_lut_adj_439.LUT_INIT = 16'hbebe;
    SB_LUT4 select_238_Select_4_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [4]), .I3(GND_net), .O(n2_adj_2175));
    defparam select_238_Select_4_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i8_3_lut (.I0(\data_out[8][7] ), 
            .I1(\data_out[9] [7]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n8_adj_2176));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i10_4_lut (.I0(n8_adj_2176), 
            .I1(\data_out[10] [7]), .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n10_adj_7));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15538 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [5]), .I2(\data_out_frame2[11] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n17993));
    defparam byte_transmit_counter2_0__bdd_4_lut_15538.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut_adj_440 (.I0(n17013), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[1] [5]), .I3(n9743), .O(n17015));   // coms.v(130[17:124])
    defparam i2_4_lut_adj_440.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame2_0___i141 (.Q(\data_out_frame2[17] [4]), .C(CLK_c), 
           .D(n10825));   // coms.v(426[12] 547[6])
    SB_LUT4 i2_3_lut_4_lut_adj_441 (.I0(\FRAME_MATCHER.state_c [18]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(\FRAME_MATCHER.state_c [17]), .I3(n16869), .O(n56));   // coms.v(492[5:16])
    defparam i2_3_lut_4_lut_adj_441.LUT_INIT = 16'hfffe;
    SB_DFF delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .D(n10859));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_1[[6__2267  (.Q(\data_in[1] [6]), .C(CLK_c), .D(n10672));   // coms.v(426[12] 547[6])
    SB_LUT4 add_2495_14_lut (.I0(n29), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n15525), .O(n17575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_14_lut.LUT_INIT = 16'h8228;
    SB_DFF \data_in_1[[5__2268  (.Q(\data_in[1] [5]), .C(CLK_c), .D(n10671));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_1[[4__2269  (.Q(\data_in[1] [4]), .C(CLK_c), .D(n10670));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_1[[6__2230  (.Q(\data_out[1][6] ), .C(CLK_c), .D(n10367));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_1[[3__2270  (.Q(\data_in[1] [3]), .C(CLK_c), .D(n10669));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_5_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [5]), .I3(GND_net), .O(n2_adj_2179));
    defparam select_238_Select_5_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_in_1[[2__2271  (.Q(\data_in[1] [2]), .C(CLK_c), .D(n10668));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_1[[1__2272  (.Q(\data_in[1] [1]), .C(CLK_c), .D(n10667));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_6_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [6]), .I3(GND_net), .O(n2_adj_2180));
    defparam select_238_Select_6_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_7_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [7]), .I3(GND_net), .O(n2_adj_2181));
    defparam select_238_Select_7_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_out_1[[7__2229  (.Q(\data_out[1][7] ), .C(CLK_c), .D(n10366));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_1[[0__2273  (.Q(\data_in[1] [0]), .C(CLK_c), .D(n10666));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_8_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [8]), .I3(GND_net), .O(n2_adj_2182));
    defparam select_238_Select_8_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i12_4_lut (.I0(n23_adj_2156), .I1(\data_in_frame[9] [1]), .I2(n17014), 
            .I3(n17001), .O(n28_adj_2183));   // coms.v(513[9:61])
    defparam i12_4_lut.LUT_INIT = 16'hbfef;
    SB_LUT4 i10_4_lut_adj_442 (.I0(n19), .I1(n15929), .I2(n2336), .I3(\data_in_frame[10] [5]), 
            .O(n26_adj_2184));   // coms.v(513[9:61])
    defparam i10_4_lut_adj_442.LUT_INIT = 16'hbffb;
    SB_DFF delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .D(n10858));   // coms.v(280[12] 380[6])
    SB_DFF \data_in_0[[7__2274  (.Q(\data_in[0] [7]), .C(CLK_c), .D(n10665));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut (.I0(byte_transmit_counter2[2]), 
            .I1(n17960), .I2(n17954), .I3(byte_transmit_counter2[3]), 
            .O(n18125));
    defparam byte_transmit_counter2_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 select_238_Select_9_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [9]), .I3(GND_net), .O(n2_adj_2185));
    defparam select_238_Select_9_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_10_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [10]), .I3(GND_net), .O(n2_adj_2186));
    defparam select_238_Select_10_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_in_0[[6__2275  (.Q(\data_in[0] [6]), .C(CLK_c), .D(n10664));   // coms.v(426[12] 547[6])
    SB_LUT4 n18125_bdd_4_lut (.I0(n18125), .I1(n6_adj_2187), .I2(n17576), 
            .I3(byte_transmit_counter2[3]), .O(n18128));
    defparam n18125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1210_i1_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n2651[0]));   // coms.v(283[4] 379[11])
    defparam mux_1210_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15616 (.I0(byte_transmit_counter[1]), 
            .I1(n17569), .I2(n5_adj_2188), .I3(\byte_transmit_counter[2] ), 
            .O(n18041));
    defparam byte_transmit_counter_1__bdd_4_lut_15616.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [18]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(n12_adj_2189), .I3(n16905), .O(n9460));   // coms.v(492[5:16])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \data_in_0[[5__2276  (.Q(\data_in[0] [5]), .C(CLK_c), .D(n10663));   // coms.v(426[12] 547[6])
    SB_LUT4 i2_3_lut_4_lut_adj_443 (.I0(\FRAME_MATCHER.state_c [18]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(n61), .I3(n59), .O(n16133));   // coms.v(492[5:16])
    defparam i2_3_lut_4_lut_adj_443.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15641 (.I0(byte_transmit_counter2[2]), 
            .I1(n17942), .I2(n17936), .I3(byte_transmit_counter2[3]), 
            .O(n18119));
    defparam byte_transmit_counter2_2__bdd_4_lut_15641.LUT_INIT = 16'he4aa;
    SB_LUT4 select_238_Select_11_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [11]), .I3(GND_net), .O(n2_adj_2190));
    defparam select_238_Select_11_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i2_2_lut_adj_444 (.I0(\data_out_frame2[0] [6]), .I1(\data_out_frame2[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_2191));   // coms.v(234[16:291])
    defparam i2_2_lut_adj_444.LUT_INIT = 16'h6666;
    SB_LUT4 select_238_Select_12_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [12]), .I3(GND_net), .O(n2_adj_2192));
    defparam select_238_Select_12_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i6_4_lut_adj_445 (.I0(\data_out_frame2[9] [3]), .I1(n17085), 
            .I2(n17073), .I3(n17127), .O(n14));   // coms.v(234[16:291])
    defparam i6_4_lut_adj_445.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_446 (.I0(n9688), .I1(n14), .I2(n10_adj_2191), 
            .I3(\data_out_frame2[12] [7]), .O(n17128));   // coms.v(234[16:291])
    defparam i7_4_lut_adj_446.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_447 (.I0(\data_out_frame2[14] [5]), .I1(n9692), 
            .I2(\data_out_frame2[7] [5]), .I3(GND_net), .O(n17085));   // coms.v(233[16:291])
    defparam i2_3_lut_adj_447.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_448 (.I0(n9810), .I1(\data_out_frame2[9] [6]), 
            .I2(\data_out_frame2[7] [4]), .I3(\data_out_frame2[8] [0]), 
            .O(n16));   // coms.v(233[16:291])
    defparam i6_4_lut_adj_448.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_449 (.I0(\data_out_frame2[10] [0]), .I1(n16923), 
            .I2(n9819), .I3(n17031), .O(n17_adj_2193));   // coms.v(233[16:291])
    defparam i7_4_lut_adj_449.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17_adj_2193), .I1(n17085), .I2(n16), .I3(n17124), 
            .O(n17125));   // coms.v(233[16:291])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_450 (.I0(\data_out_frame2[0] [4]), .I1(\data_out_frame2[14] [4]), 
            .I2(\data_out_frame2[15] [4]), .I3(GND_net), .O(n17124));   // coms.v(233[16:291])
    defparam i2_3_lut_adj_450.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_451 (.I0(\data_out_frame2[7] [7]), .I1(n16926), 
            .I2(\data_out_frame2[14] [3]), .I3(n17022), .O(n22_adj_2194));   // coms.v(232[16:229])
    defparam i9_4_lut_adj_451.LUT_INIT = 16'h6996;
    SB_LUT4 select_238_Select_13_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [13]), .I3(GND_net), .O(n2_adj_2195));
    defparam select_238_Select_13_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_in_0[[4__2277  (.Q(\data_in[0] [4]), .C(CLK_c), .D(n10662));   // coms.v(426[12] 547[6])
    SB_LUT4 i11_4_lut_adj_452 (.I0(n21_adj_2171), .I1(n15930), .I2(n2340), 
            .I3(\data_in_frame[10] [7]), .O(n27_adj_2196));   // coms.v(513[9:61])
    defparam i11_4_lut_adj_452.LUT_INIT = 16'hbffb;
    SB_LUT4 i11_4_lut_adj_453 (.I0(n9913), .I1(n22_adj_2194), .I2(n16_adj_2197), 
            .I3(\data_out_frame2[9] [3]), .O(n24));   // coms.v(232[16:229])
    defparam i11_4_lut_adj_453.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_454 (.I0(n9485), .I1(\data_in[2] [0]), .I2(\data_in[0] [1]), 
            .I3(n9490), .O(n18_adj_2198));
    defparam i7_4_lut_adj_454.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_455 (.I0(n17015), .I1(n18_adj_2174), .I2(n2338), 
            .I3(\data_in_frame[10] [6]), .O(n25));   // coms.v(513[9:61])
    defparam i9_4_lut_adj_455.LUT_INIT = 16'hdffd;
    SB_LUT4 i14818_4_lut (.I0(\data_in[0] [0]), .I1(\data_in[3] [5]), .I2(\data_in[1] [6]), 
            .I3(\data_in[3] [7]), .O(n17256));
    defparam i14818_4_lut.LUT_INIT = 16'h8000;
    SB_DFF \data_in_0[[3__2278  (.Q(\data_in[0] [3]), .C(CLK_c), .D(n10661));   // coms.v(426[12] 547[6])
    SB_LUT4 i8_4_lut (.I0(\data_in[0] [3]), .I1(\data_in[2] [2]), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [7]), .O(n19_adj_2199));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_456 (.I0(n19_adj_2199), .I1(n17256), .I2(n18_adj_2198), 
            .I3(n12_adj_2200), .O(n127_adj_2136));
    defparam i10_4_lut_adj_456.LUT_INIT = 16'hfffb;
    SB_LUT4 n18119_bdd_4_lut (.I0(n18119), .I1(n6_adj_2201), .I2(n17578), 
            .I3(byte_transmit_counter2[3]), .O(n18122));
    defparam n18119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_457 (.I0(\FRAME_MATCHER.state_c [7]), .I1(\FRAME_MATCHER.state_c [15]), 
            .I2(\FRAME_MATCHER.state_c [13]), .I3(\FRAME_MATCHER.state_c [11]), 
            .O(n16772));   // coms.v(457[5:29])
    defparam i3_4_lut_adj_457.LUT_INIT = 16'hfffe;
    SB_DFF \data_in_0[[2__2279  (.Q(\data_in[0] [2]), .C(CLK_c), .D(n10660));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_458 (.I0(\FRAME_MATCHER.state_c [29]), .I1(\FRAME_MATCHER.state_c [27]), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // coms.v(426[12] 547[6])
    defparam i1_2_lut_adj_458.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_459 (.I0(n17079), .I1(n24), .I2(n20_adj_2202), 
            .I3(n17115), .O(n17126));   // coms.v(232[16:229])
    defparam i12_4_lut_adj_459.LUT_INIT = 16'h9669;
    SB_CARRY add_2495_14 (.CI(n15525), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n15526));
    SB_LUT4 i15_4_lut_adj_460 (.I0(n25), .I1(n27_adj_2196), .I2(n26_adj_2184), 
            .I3(n28_adj_2183), .O(n15846));   // coms.v(513[9:61])
    defparam i15_4_lut_adj_460.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter2_2353_add_4_2_lut (.I0(GND_net), .I1(tx2_transmit_N_1997), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY byte_transmit_counter2_2353_add_4_2 (.CI(GND_net), .I0(tx2_transmit_N_1997), 
            .I1(byte_transmit_counter2[0]), .CO(n15615));
    SB_LUT4 select_238_Select_14_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [14]), .I3(GND_net), .O(n2_adj_2204));
    defparam select_238_Select_14_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_adj_461 (.I0(delay_counter[11]), .I1(delay_counter[10]), 
            .I2(GND_net), .I3(GND_net), .O(n12993));   // coms.v(280[12] 380[6])
    defparam i1_2_lut_adj_461.LUT_INIT = 16'heeee;
    SB_DFF \data_in_0[[1__2280  (.Q(\data_in[0] [1]), .C(CLK_c), .D(n10659));   // coms.v(426[12] 547[6])
    SB_DFF \data_in_0[[0__2281  (.Q(\data_in[0] [0]), .C(CLK_c), .D(n10658));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_462 (.I0(delay_counter[3]), .I1(delay_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n13298));   // coms.v(280[12] 380[6])
    defparam i1_2_lut_adj_462.LUT_INIT = 16'heeee;
    SB_LUT4 i8_4_lut_adj_463 (.I0(\data_out_frame2[14] [3]), .I1(\data_out_frame2[16] [0]), 
            .I2(\data_out_frame2[9] [2]), .I3(n9892), .O(n20_adj_2205));   // coms.v(237[17:221])
    defparam i8_4_lut_adj_463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_464 (.I0(delay_counter[9]), .I1(delay_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n12991));   // coms.v(280[12] 380[6])
    defparam i1_2_lut_adj_464.LUT_INIT = 16'heeee;
    SB_LUT4 select_238_Select_15_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [15]), .I3(GND_net), .O(n2_adj_2206));
    defparam select_238_Select_15_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF byte_transmit_counter__i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
           .D(n16247));   // coms.v(280[12] 380[6])
    SB_LUT4 i10_4_lut_adj_465 (.I0(n9859), .I1(n20_adj_2205), .I2(\data_out_frame2[9] [0]), 
            .I3(n9555), .O(n22_adj_2207));   // coms.v(237[17:221])
    defparam i10_4_lut_adj_465.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15552 (.I0(byte_transmit_counter[1]), 
            .I1(n17543), .I2(n5_adj_2208), .I3(\byte_transmit_counter[2] ), 
            .O(n18011));
    defparam byte_transmit_counter_1__bdd_4_lut_15552.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_2209), .S(n3_adj_2210));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_16_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [16]), .I3(GND_net), .O(n2_adj_2211));
    defparam select_238_Select_16_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_adj_466 (.I0(\FRAME_MATCHER.state_c [22]), .I1(\FRAME_MATCHER.state_c [21]), 
            .I2(GND_net), .I3(GND_net), .O(n61));   // coms.v(426[12] 547[6])
    defparam i1_2_lut_adj_466.LUT_INIT = 16'heeee;
    SB_LUT4 select_238_Select_17_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [17]), .I3(GND_net), .O(n2_adj_2212));
    defparam select_238_Select_17_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_adj_467 (.I0(\FRAME_MATCHER.state_c [6]), .I1(\FRAME_MATCHER.state_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2213));   // coms.v(448[5:27])
    defparam i1_2_lut_adj_467.LUT_INIT = 16'heeee;
    SB_LUT4 i14914_3_lut (.I0(\data_out_frame2[0] [0]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17352));
    defparam i14914_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_2214), .S(n3_adj_2215));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_2216), .S(n3_adj_2217));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_2218), .S(n3_adj_2219));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_2220), .S(n3_adj_2221));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_2222), .S(n3_adj_2223));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_2224), .S(n3_adj_2225));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_2226), .S(n3_adj_2227));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_2228), .S(n3_adj_2229));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_2230), .S(n3_adj_2231));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_2232), .S(n3_adj_2233));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_2234), .S(n3_adj_2235));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_2236), .S(n3_adj_2237));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_2238), .S(n3_adj_2239));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_2212), .S(n3_adj_2240));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_2211), .S(n3_adj_2241));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_2206), .S(n3_adj_2242));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_2204), .S(n3_adj_2243));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_2195), .S(n3_adj_2244));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_2192), .S(n3_adj_2245));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_2190), .S(n3_adj_2246));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_2186), .S(n3_adj_2247));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_2185), .S(n3_adj_2248));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_2182), .S(n3_adj_2249));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_2181), .S(n3_adj_2250));   // coms.v(426[12] 547[6])
    SB_LUT4 i4_4_lut_adj_468 (.I0(\FRAME_MATCHER.state_c [12]), .I1(\FRAME_MATCHER.state_c [10]), 
            .I2(\FRAME_MATCHER.state_c [9]), .I3(n6_adj_2213), .O(n16869));   // coms.v(448[5:27])
    defparam i4_4_lut_adj_468.LUT_INIT = 16'hfffe;
    SB_LUT4 i14916_4_lut (.I0(n17352), .I1(n15846), .I2(n5543), .I3(n5545), 
            .O(n17354));
    defparam i14916_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i11_4_lut_adj_469 (.I0(n16946), .I1(n22_adj_2207), .I2(n18_adj_2251), 
            .I3(n17040), .O(n17123));   // coms.v(237[17:221])
    defparam i11_4_lut_adj_469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_470 (.I0(\data_out_frame2[7] [2]), .I1(\data_out_frame2[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17121));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_470.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1522_i1_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n3071[0]));   // coms.v(283[4] 379[11])
    defparam mux_1522_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15636 (.I0(byte_transmit_counter2[2]), 
            .I1(n17924), .I2(n17918), .I3(byte_transmit_counter2[3]), 
            .O(n18107));
    defparam byte_transmit_counter2_2__bdd_4_lut_15636.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_471 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n16869), 
            .I2(GND_net), .I3(GND_net), .O(n16871));   // coms.v(448[5:27])
    defparam i1_2_lut_adj_471.LUT_INIT = 16'heeee;
    SB_LUT4 select_238_Select_18_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [18]), .I3(GND_net), .O(n2_adj_2238));
    defparam select_238_Select_18_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 n18041_bdd_4_lut (.I0(n18041), .I1(n2_adj_2137), .I2(n17585), 
            .I3(\byte_transmit_counter[2] ), .O(n18044));
    defparam n18041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_472 (.I0(\data_out_frame2[11] [4]), .I1(\data_out_frame2[9] [5]), 
            .I2(n9678), .I3(n16940), .O(n20_adj_2252));   // coms.v(230[16:237])
    defparam i8_4_lut_adj_472.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_2180), .S(n3_adj_2253));   // coms.v(426[12] 547[6])
    SB_LUT4 add_2495_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n15524), .O(n6517[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_473 (.I0(\data_out_frame2[0] [2]), .I1(n9901), 
            .I2(n9754), .I3(\data_out_frame2[9] [1]), .O(n19_adj_2254));   // coms.v(230[16:237])
    defparam i7_4_lut_adj_473.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_474 (.I0(n16994), .I1(n17082), .I2(n17052), .I3(n17121), 
            .O(n21_adj_2255));   // coms.v(230[16:237])
    defparam i9_4_lut_adj_474.LUT_INIT = 16'h6996;
    SB_DFF \data_out_2[[0__2228  (.Q(\data_out[2][0] ), .C(CLK_c), .D(n10365));   // coms.v(280[12] 380[6])
    SB_LUT4 n18107_bdd_4_lut (.I0(n18107), .I1(n6_c), .I2(n17579), .I3(byte_transmit_counter2[3]), 
            .O(n18110));
    defparam n18107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1080_i1_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\rand_setpoint[25] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(\UART_TRANSMITTER.state[0] ), 
            .O(n2476[0]));   // coms.v(283[4] 379[11])
    defparam mux_1080_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_3_lut (.I0(n21_adj_2255), .I1(n19_adj_2254), .I2(n20_adj_2252), 
            .I3(GND_net), .O(n17122));   // coms.v(230[16:237])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_475 (.I0(\data_out_frame2[11] [0]), .I1(\data_out_frame2[10] [7]), 
            .I2(\data_out_frame2[11] [3]), .I3(n16908), .O(n17022));   // coms.v(232[16:229])
    defparam i3_4_lut_adj_475.LUT_INIT = 16'h6996;
    SB_LUT4 select_238_Select_19_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [19]), .I3(GND_net), .O(n2_adj_2236));
    defparam select_238_Select_19_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_20_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [20]), .I3(GND_net), .O(n2_adj_2234));
    defparam select_238_Select_20_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_2179), .S(n3_adj_2256));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_2175), .S(n3_adj_2257));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [0]), .I2(\data_out_frame2[19] [0]), 
            .I3(byte_transmit_counter2[1]), .O(n18101));
    defparam byte_transmit_counter2_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_2173), .S(n3_adj_2258));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_21_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [21]), .I3(GND_net), .O(n2_adj_2232));
    defparam select_238_Select_21_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_2172), .S(n3_adj_2259));   // coms.v(426[12] 547[6])
    SB_LUT4 n18101_bdd_4_lut (.I0(n18101), .I1(\data_out_frame2[17] [0]), 
            .I2(\data_out_frame2[16] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n18104));
    defparam n18101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_2168), .S(n3_adj_2260));   // coms.v(426[12] 547[6])
    SB_DFFSR tx2_transmit_2249 (.Q(r_SM_Main_2__N_2036_adj_2400[0]), .C(CLK_c), 
            .D(n4130[0]), .R(n13496));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_4_lut_adj_476 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n16898), 
            .I2(n59), .I3(n16772), .O(n5_adj_2262));   // coms.v(457[5:29])
    defparam i1_4_lut_adj_476.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_477 (.I0(n16966), .I1(\data_out[8][5] ), .I2(n9728), 
            .I3(GND_net), .O(data_out_9__0__N_389));   // coms.v(21[11:19])
    defparam i2_3_lut_adj_477.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_478 (.I0(\data_out_frame2[10] [6]), .I1(n17022), 
            .I2(GND_net), .I3(GND_net), .O(n9555));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_478.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15606 (.I0(byte_transmit_counter2[2]), 
            .I1(n17393), .I2(n17894), .I3(byte_transmit_counter2[3]), 
            .O(n17963));
    defparam byte_transmit_counter2_2__bdd_4_lut_15606.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_479 (.I0(n5_adj_2262), .I1(n52), .I2(\FRAME_MATCHER.state_c [26]), 
            .I3(\FRAME_MATCHER.state_c [25]), .O(n16876));   // coms.v(457[5:29])
    defparam i3_4_lut_adj_479.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_480 (.I0(\data_out_frame2[14] [1]), .I1(n9555), 
            .I2(\data_out_frame2[0] [1]), .I3(n9763), .O(n17052));   // coms.v(229[16:299])
    defparam i3_4_lut_adj_480.LUT_INIT = 16'h6996;
    SB_LUT4 i15246_2_lut (.I0(\rand_setpoint[17] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17506));   // coms.v(283[4] 379[11])
    defparam i15246_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS \data_out_5[[0__2204  (.Q(data_out_6__1__N_537), .C(CLK_c), 
            .E(n10055), .D(n2502[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 select_238_Select_22_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [22]), .I3(GND_net), .O(n2_adj_2230));
    defparam select_238_Select_22_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i5_4_lut_adj_481 (.I0(\data_out_frame2[7] [0]), .I1(\data_out_frame2[9] [0]), 
            .I2(n9853), .I3(n16960), .O(n12_adj_2263));   // coms.v(229[16:299])
    defparam i5_4_lut_adj_481.LUT_INIT = 16'h6996;
    SB_LUT4 select_238_Select_23_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [23]), .I3(GND_net), .O(n2_adj_2228));
    defparam select_238_Select_23_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_24_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [24]), .I3(GND_net), .O(n2_adj_2226));
    defparam select_238_Select_24_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_25_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [25]), .I3(GND_net), .O(n2_adj_2224));
    defparam select_238_Select_25_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFF \data_out_2[[2__2226  (.Q(\data_out[2][2] ), .C(CLK_c), .D(n10364));   // coms.v(280[12] 380[6])
    SB_LUT4 i6_4_lut_adj_482 (.I0(n17052), .I1(n12_adj_2263), .I2(\data_out_frame2[7] [4]), 
            .I3(n9886), .O(n17053));   // coms.v(229[16:299])
    defparam i6_4_lut_adj_482.LUT_INIT = 16'h9669;
    SB_LUT4 add_2495_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n15517), .O(n6517[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_872_i1_4_lut (.I0(data_out_6__1__N_537), .I1(n17506), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n2196[0]));   // coms.v(283[4] 379[11])
    defparam mux_872_i1_4_lut.LUT_INIT = 16'hcacf;
    SB_LUT4 select_238_Select_26_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [26]), .I3(GND_net), .O(n2_adj_2222));
    defparam select_238_Select_26_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i5_3_lut (.I0(n17103), .I1(n9919), .I2(\data_out_frame2[5] [4]), 
            .I3(GND_net), .O(n14_adj_2264));   // coms.v(228[16:596])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_238_Select_27_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [27]), .I3(GND_net), .O(n2_adj_2220));
    defparam select_238_Select_27_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 select_238_Select_28_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [28]), .I3(GND_net), .O(n2_adj_2218));
    defparam select_238_Select_28_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n17632), .I2(n5_adj_2265), .I3(\byte_transmit_counter[2] ), 
            .O(n18095));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18095_bdd_4_lut (.I0(n18095), .I1(n2_adj_2266), .I2(n17581), 
            .I3(\byte_transmit_counter[2] ), .O(n18098));
    defparam n18095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS \data_out_5[[2__2202  (.Q(\data_out[5] [2]), .C(CLK_c), .E(n10055), 
            .D(n2432[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 i8_4_lut_adj_483 (.I0(delay_counter[4]), .I1(delay_counter[14]), 
            .I2(delay_counter[13]), .I3(delay_counter[0]), .O(n20_adj_2267));   // coms.v(272[12:25])
    defparam i8_4_lut_adj_483.LUT_INIT = 16'hfffe;
    SB_DFFESS \data_out_5[[3__2201  (.Q(\data_out[5] [3]), .C(CLK_c), .E(n10055), 
            .D(n2397[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 select_238_Select_29_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [29]), .I3(GND_net), .O(n2_adj_2216));
    defparam select_238_Select_29_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i4_4_lut_adj_484 (.I0(n9496), .I1(\data_out[6] [5]), .I2(n9716), 
            .I3(\data_out[6] [7]), .O(n10_adj_2268));   // coms.v(179[16:84])
    defparam i4_4_lut_adj_484.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_485 (.I0(\data_out[8]_c [3]), .I1(n10_adj_2268), 
            .I2(\data_out[8][4] ), .I3(GND_net), .O(data_out_9__1__N_378));   // coms.v(179[16:84])
    defparam i5_3_lut_adj_485.LUT_INIT = 16'h9696;
    SB_LUT4 i15245_3_lut (.I0(\data_out[5] [1]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(data_out_6__1__N_537), .I3(GND_net), .O(n17507));   // coms.v(283[4] 379[11])
    defparam i15245_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i6_4_lut_adj_486 (.I0(\data_out_frame2[9] [2]), .I1(\data_out_frame2[11] [0]), 
            .I2(\data_out_frame2[12] [4]), .I3(n16957), .O(n15_adj_2269));   // coms.v(228[16:596])
    defparam i6_4_lut_adj_486.LUT_INIT = 16'h6996;
    SB_LUT4 select_238_Select_31_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [31]), .I3(GND_net), .O(n2_adj_2209));
    defparam select_238_Select_31_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i8_4_lut_adj_487 (.I0(n15_adj_2269), .I1(n17046), .I2(n14_adj_2264), 
            .I3(n17097), .O(n17105));   // coms.v(228[16:596])
    defparam i8_4_lut_adj_487.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_488 (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[13] [7]), 
            .I2(n9758), .I3(\data_out_frame2[15] [5]), .O(n17073));   // coms.v(234[16:291])
    defparam i3_4_lut_adj_488.LUT_INIT = 16'h6996;
    SB_LUT4 mux_846_i1_4_lut (.I0(n17507), .I1(\rand_setpoint[18] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2161[0]));   // coms.v(283[4] 379[11])
    defparam mux_846_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7_4_lut_adj_489 (.I0(n12991), .I1(delay_counter[8]), .I2(delay_counter[5]), 
            .I3(delay_counter[2]), .O(n19_adj_2270));   // coms.v(272[12:25])
    defparam i7_4_lut_adj_489.LUT_INIT = 16'hfffe;
    SB_LUT4 i15249_3_lut (.I0(\data_out[5] [2]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [1]), .I3(GND_net), .O(n17514));   // coms.v(283[4] 379[11])
    defparam i15249_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_adj_490 (.I0(\data_out_frame2[6] [2]), .I1(\data_out_frame2[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17031));   // coms.v(233[16:291])
    defparam i1_2_lut_adj_490.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_491 (.I0(delay_counter[7]), .I1(n13298), .I2(n12993), 
            .I3(delay_counter[12]), .O(n21_adj_2271));   // coms.v(272[12:25])
    defparam i9_4_lut_adj_491.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_492 (.I0(\data_out_frame2[5] [6]), .I1(\data_out_frame2[6] [7]), 
            .I2(\data_out_frame2[5] [7]), .I3(n9678), .O(n24_adj_2272));   // coms.v(239[17:230])
    defparam i9_4_lut_adj_492.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_493 (.I0(n17031), .I1(n17073), .I2(n17049), 
            .I3(n17091), .O(n26_adj_2273));   // coms.v(239[17:230])
    defparam i11_4_lut_adj_493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_494 (.I0(\data_out[8][6] ), .I1(\data_out[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2274));   // coms.v(182[17:86])
    defparam i1_2_lut_adj_494.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_495 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state_c [28]), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(\FRAME_MATCHER.state_c [17]), 
            .O(n16761));   // coms.v(457[5:29])
    defparam i3_4_lut_adj_495.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_820_i1_4_lut (.I0(n17514), .I1(\rand_setpoint[19] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2126[0]));   // coms.v(283[4] 379[11])
    defparam mux_820_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i5_4_lut_adj_496 (.I0(n16761), .I1(n16876), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(n16871), .O(n12_adj_2189));   // coms.v(492[5:16])
    defparam i5_4_lut_adj_496.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut_adj_497 (.I0(\data_out[7] [0]), .I1(n17058), .I2(n16969), 
            .I3(n6_adj_2274), .O(data_out_9__4__N_345));   // coms.v(182[17:86])
    defparam i4_4_lut_adj_497.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_498 (.I0(\data_out_frame2[8] [1]), .I1(n16987), 
            .I2(n9814), .I3(n17010), .O(n25_adj_2275));   // coms.v(239[17:230])
    defparam i10_4_lut_adj_498.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_499 (.I0(\data_out[5] [3]), .I1(\data_out[8][7] ), 
            .I2(\data_out[9] [1]), .I3(\data_out[9] [0]), .O(n16969));   // coms.v(182[17:86])
    defparam i3_4_lut_adj_499.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_500 (.I0(\data_out[10] [5]), .I1(n16969), .I2(\data_out[7] [1]), 
            .I3(n17055), .O(data_out_9__5__N_334));   // coms.v(182[17:86])
    defparam i3_4_lut_adj_500.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_501 (.I0(n9530), .I1(\data_out[9] [0]), .I2(\data_out[10] [6]), 
            .I3(\data_out[7] [4]), .O(n10_adj_2276));   // coms.v(184[17:86])
    defparam i4_4_lut_adj_501.LUT_INIT = 16'h6996;
    SB_LUT4 select_238_Select_30_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [30]), .I3(GND_net), .O(n2_adj_2214));
    defparam select_238_Select_30_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15626 (.I0(byte_transmit_counter2[2]), 
            .I1(n18074), .I2(n18068), .I3(byte_transmit_counter2[3]), 
            .O(n18089));
    defparam byte_transmit_counter2_2__bdd_4_lut_15626.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_502 (.I0(n17133), .I1(n24_adj_2272), .I2(\data_out_frame2[13] [2]), 
            .I3(n9859), .O(n27_adj_2277));   // coms.v(239[17:230])
    defparam i12_4_lut_adj_502.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_503 (.I0(\data_out_frame2[0] [5]), .I1(n27_adj_2277), 
            .I2(n25_adj_2275), .I3(n26_adj_2273), .O(n17103));   // coms.v(227[16:31])
    defparam i1_4_lut_adj_503.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_504 (.I0(\data_out[9] [3]), .I1(n10_adj_2276), 
            .I2(n16981), .I3(GND_net), .O(data_out_9__6__N_324));   // coms.v(184[17:86])
    defparam i5_3_lut_adj_504.LUT_INIT = 16'h6969;
    SB_LUT4 n18089_bdd_4_lut (.I0(n18089), .I1(n6_adj_2278), .I2(n17561), 
            .I3(byte_transmit_counter2[3]), .O(n18092));
    defparam n18089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \UART_TRANSMITTER.state_i0_i2  (.Q(\UART_TRANSMITTER.state[2] ), 
           .C(CLK_c), .D(n33));   // coms.v(280[12] 380[6])
    SB_LUT4 n17963_bdd_4_lut (.I0(n17963), .I1(n6_adj_2280), .I2(n17571), 
            .I3(byte_transmit_counter2[3]), .O(n17966));
    defparam n17963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_505 (.I0(\data_out_frame2[11] [2]), .I1(\data_out_frame2[15] [0]), 
            .I2(\data_out_frame2[0] [0]), .I3(n16972), .O(n10_adj_2281));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_505.LUT_INIT = 16'h6996;
    SB_LUT4 i15210_3_lut (.I0(\data_out[5] [3]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [2]), .I3(GND_net), .O(n17518));   // coms.v(283[4] 379[11])
    defparam i15210_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_adj_506 (.I0(\data_out[7] [2]), .I1(\data_out[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17058));   // coms.v(182[17:86])
    defparam i1_2_lut_adj_506.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15514 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [3]), .I2(\data_out_frame2[11] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n17957));
    defparam byte_transmit_counter2_0__bdd_4_lut_15514.LUT_INIT = 16'he4aa;
    SB_LUT4 n17957_bdd_4_lut (.I0(n17957), .I1(\data_out_frame2[9] [3]), 
            .I2(\data_out_frame2[8] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n17960));
    defparam n17957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_794_i1_4_lut (.I0(n17518), .I1(\rand_setpoint[20] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2091[0]));   // coms.v(283[4] 379[11])
    defparam mux_794_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15505 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [3]), .I2(\data_out_frame2[15] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n17951));
    defparam byte_transmit_counter2_0__bdd_4_lut_15505.LUT_INIT = 16'he4aa;
    SB_LUT4 add_2495_2_lut (.I0(n53), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n17637)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 select_238_Select_0_i2_2_lut_3_lut (.I0(n9452), .I1(n12933), 
            .I2(\FRAME_MATCHER.i_31__N_1280 [0]), .I3(GND_net), .O(n2_adj_2159));
    defparam select_238_Select_0_i2_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 n17951_bdd_4_lut (.I0(n17951), .I1(\data_out_frame2[13] [3]), 
            .I2(\data_out_frame2[12] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n17954));
    defparam n17951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_507 (.I0(n16912), .I1(n16978), .I2(n16975), .I3(n16998), 
            .O(n20_adj_2282));   // coms.v(182[17:86])
    defparam i8_4_lut_adj_507.LUT_INIT = 16'h6996;
    SB_LUT4 i15395_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), .I2(n9460), 
            .I3(n491), .O(n17452));
    defparam i15395_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i15211_3_lut (.I0(\data_out[5] [4]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [3]), .I3(GND_net), .O(n17522));   // coms.v(283[4] 379[11])
    defparam i15211_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i5_3_lut_adj_508 (.I0(n17061), .I1(n10_adj_2281), .I2(n17103), 
            .I3(GND_net), .O(n17104));   // coms.v(227[16:31])
    defparam i5_3_lut_adj_508.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15500 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [3]), .I2(\data_out_frame2[19] [3]), 
            .I3(byte_transmit_counter2[1]), .O(n17945));
    defparam byte_transmit_counter2_0__bdd_4_lut_15500.LUT_INIT = 16'he4aa;
    SB_LUT4 n17945_bdd_4_lut (.I0(n17945), .I1(\data_out_frame2[17] [3]), 
            .I2(\data_out_frame2[16] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n17948));
    defparam n17945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_509 (.I0(\data_out[9] [5]), .I1(\data_out[5] [4]), 
            .I2(\data_out[5] [3]), .I3(n9522), .O(n19_adj_2283));   // coms.v(182[17:86])
    defparam i7_4_lut_adj_509.LUT_INIT = 16'h6996;
    SB_LUT4 mux_768_i1_4_lut (.I0(n17522), .I1(\rand_setpoint[21] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2056[0]));   // coms.v(283[4] 379[11])
    defparam mux_768_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_510 (.I0(\data_out_frame2[15] [1]), .I1(\data_out_frame2[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9678));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_510.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15495 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [2]), .I2(\data_out_frame2[11] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n17939));
    defparam byte_transmit_counter2_0__bdd_4_lut_15495.LUT_INIT = 16'he4aa;
    SB_LUT4 n17939_bdd_4_lut (.I0(n17939), .I1(\data_out_frame2[9] [2]), 
            .I2(\data_out_frame2[8] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n17942));
    defparam n17939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \data_out_2[[3__2225  (.Q(\data_out[2] [3]), .C(CLK_c), .D(n10363));   // coms.v(280[12] 380[6])
    SB_LUT4 i15256_3_lut (.I0(\data_out[5] [5]), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [4]), .I3(GND_net), .O(n17528));   // coms.v(283[4] 379[11])
    defparam i15256_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15490 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [2]), .I2(\data_out_frame2[15] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n17933));
    defparam byte_transmit_counter2_0__bdd_4_lut_15490.LUT_INIT = 16'he4aa;
    SB_LUT4 i9_4_lut_adj_511 (.I0(n17007), .I1(n17058), .I2(n17028), .I3(n17094), 
            .O(n21_adj_2284));   // coms.v(182[17:86])
    defparam i9_4_lut_adj_511.LUT_INIT = 16'h6996;
    SB_LUT4 n17933_bdd_4_lut (.I0(n17933), .I1(\data_out_frame2[13] [2]), 
            .I2(\data_out_frame2[12] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n17936));
    defparam n17933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_742_i1_4_lut (.I0(n17528), .I1(\rand_setpoint[22] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n2021[0]));   // coms.v(283[4] 379[11])
    defparam mux_742_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15485 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [2]), .I2(\data_out_frame2[19] [2]), 
            .I3(byte_transmit_counter2[1]), .O(n17927));
    defparam byte_transmit_counter2_0__bdd_4_lut_15485.LUT_INIT = 16'he4aa;
    SB_LUT4 i11_3_lut_adj_512 (.I0(n21_adj_2284), .I1(n19_adj_2283), .I2(n20_adj_2282), 
            .I3(GND_net), .O(data_out_9__7__N_272));   // coms.v(182[17:86])
    defparam i11_3_lut_adj_512.LUT_INIT = 16'h6969;
    SB_LUT4 n17927_bdd_4_lut (.I0(n17927), .I1(\data_out_frame2[17] [2]), 
            .I2(\data_out_frame2[16] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n17930));
    defparam n17927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_513 (.I0(data_out_7__2__N_447), .I1(data_out_7__3__N_441), 
            .I2(GND_net), .I3(GND_net), .O(n16912));   // coms.v(130[17:68])
    defparam i1_2_lut_adj_513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_514 (.I0(\data_out_frame2[6] [1]), .I1(\data_out_frame2[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17115));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_514.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15480 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[10] [1]), .I2(\data_out_frame2[11] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n17921));
    defparam byte_transmit_counter2_0__bdd_4_lut_15480.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_4_lut_adj_515 (.I0(n9783), .I1(n17070), .I2(n9737), .I3(n17076), 
            .O(n12_adj_2285));   // coms.v(173[16:77])
    defparam i5_4_lut_adj_515.LUT_INIT = 16'h6996;
    SB_LUT4 n17921_bdd_4_lut (.I0(n17921), .I1(\data_out_frame2[9] [1]), 
            .I2(\data_out_frame2[8] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n17924));
    defparam n17921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15475 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [1]), .I2(\data_out_frame2[15] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n17915));
    defparam byte_transmit_counter2_0__bdd_4_lut_15475.LUT_INIT = 16'he4aa;
    SB_LUT4 n17915_bdd_4_lut (.I0(n17915), .I1(\data_out_frame2[13] [1]), 
            .I2(\data_out_frame2[12] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n17918));
    defparam n17915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_516 (.I0(\data_out_frame2[7] [6]), .I1(\data_out_frame2[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16994));   // coms.v(234[16:291])
    defparam i1_2_lut_adj_516.LUT_INIT = 16'h6666;
    SB_LUT4 mux_716_i1_4_lut (.I0(n17532), .I1(\rand_setpoint[23] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1986[0]));   // coms.v(283[4] 379[11])
    defparam mux_716_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15470 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [1]), .I2(\data_out_frame2[19] [1]), 
            .I3(byte_transmit_counter2[1]), .O(n17909));
    defparam byte_transmit_counter2_0__bdd_4_lut_15470.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_517 (.I0(n17109), .I1(n12_adj_2285), .I2(\data_out[7] [3]), 
            .I3(\data_out[7] [6]), .O(data_out_10__0__N_219));   // coms.v(173[16:77])
    defparam i6_4_lut_adj_517.LUT_INIT = 16'h6996;
    SB_LUT4 n17909_bdd_4_lut (.I0(n17909), .I1(\data_out_frame2[17] [1]), 
            .I2(\data_out_frame2[16] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n17912));
    defparam n17909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_690_i1_4_lut (.I0(n17534), .I1(\rand_setpoint[8] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1951[0]));   // coms.v(283[4] 379[11])
    defparam mux_690_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_15611 (.I0(byte_transmit_counter2[2]), 
            .I1(n18050), .I2(n18008), .I3(byte_transmit_counter2[3]), 
            .O(n18083));
    defparam byte_transmit_counter2_2__bdd_4_lut_15611.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_518 (.I0(\data_out_frame2[6] [4]), .I1(\data_out_frame2[13] [6]), 
            .I2(n9707), .I3(n6_adj_2286), .O(n17133));   // coms.v(239[17:230])
    defparam i4_4_lut_adj_518.LUT_INIT = 16'h6996;
    SB_LUT4 i15417_2_lut_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n4445), .I3(\UART_TRANSMITTER.state[0] ), .O(n10054));
    defparam i15417_2_lut_3_lut_4_lut.LUT_INIT = 16'h0e00;
    SB_LUT4 i21_2_lut (.I0(\data_out[9][2] ), .I1(\data_out[5] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n9530));   // coms.v(21[11:19])
    defparam i21_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \data_out_7[[4__2184  (.Q(\data_out[7] [4]), .C(CLK_c), .E(VCC_net), 
            .D(n10839));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_519 (.I0(\FRAME_MATCHER.state [2]), .I1(n9460), 
            .I2(GND_net), .I3(GND_net), .O(n9462));   // coms.v(524[5:25])
    defparam i1_2_lut_adj_519.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_520 (.I0(\data_out_frame2[9] [2]), .I1(\data_out_frame2[5] [6]), 
            .I2(\data_out_frame2[9] [4]), .I3(GND_net), .O(n9819));   // coms.v(231[16:291])
    defparam i2_3_lut_adj_520.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_521 (.I0(\data_out[5] [2]), .I1(\data_out[6] [7]), 
            .I2(\data_out[7] [1]), .I3(\data_out[9] [0]), .O(n9522));   // coms.v(181[17:93])
    defparam i3_4_lut_adj_521.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_522 (.I0(\data_out[5] [5]), .I1(\data_out[7] [2]), 
            .I2(\data_out[9] [1]), .I3(GND_net), .O(n16981));   // coms.v(184[17:86])
    defparam i2_3_lut_adj_522.LUT_INIT = 16'h9696;
    SB_LUT4 i15441_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(data_out_10__7__N_110));   // coms.v(316[5:21])
    defparam i15441_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i3_4_lut_adj_523 (.I0(\data_out[6] [4]), .I1(n28_adj_2287), 
            .I2(\data_out[10] [4]), .I3(\data_out[10] [0]), .O(n16966));   // coms.v(21[11:19])
    defparam i3_4_lut_adj_523.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_524 (.I0(\data_out[10] [1]), .I1(\data_out[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9496));   // coms.v(171[16:93])
    defparam i1_2_lut_adj_524.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_525 (.I0(\data_out_frame2[11] [2]), .I1(\data_out_frame2[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16908));   // coms.v(235[16:291])
    defparam i1_2_lut_adj_525.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_526 (.I0(\data_out_frame2[8] [1]), .I1(n9695), 
            .I2(\data_out_frame2[0] [5]), .I3(n16908), .O(n9692));   // coms.v(235[16:291])
    defparam i3_4_lut_adj_526.LUT_INIT = 16'h6996;
    SB_LUT4 i10244_3_lut_4_lut (.I0(\data_out[8]_c [2]), .I1(\rand_setpoint[2] ), 
            .I2(\UART_TRANSMITTER.state[2] ), .I3(n2546[0]), .O(n10696));   // coms.v(21[11:19])
    defparam i10244_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i10246_3_lut_4_lut (.I0(\data_out[8]_c [3]), .I1(\rand_setpoint[3] ), 
            .I2(\UART_TRANSMITTER.state[2] ), .I3(n2546[0]), .O(n10694));   // coms.v(21[11:19])
    defparam i10246_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i4924_2_lut (.I0(n127_adj_2136), .I1(n127_adj_4), .I2(GND_net), 
            .I3(GND_net), .O(n7198));   // coms.v(437[13] 443[7])
    defparam i4924_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_527 (.I0(\data_out_frame2[0] [3]), .I1(\data_out_frame2[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16946));
    defparam i1_2_lut_adj_527.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_528 (.I0(\FRAME_MATCHER.state [2]), .I1(n9451), 
            .I2(GND_net), .I3(GND_net), .O(n9452));   // coms.v(448[5:27])
    defparam i1_2_lut_adj_528.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_529 (.I0(\data_out[10] [7]), .I1(\data_out[10] [3]), 
            .I2(n9522), .I3(GND_net), .O(n17043));   // coms.v(181[17:93])
    defparam i2_3_lut_adj_529.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_530 (.I0(\data_out[9] [7]), .I1(n16966), .I2(\data_out[9] [6]), 
            .I3(n16981), .O(n10_adj_2288));   // coms.v(178[16:77])
    defparam i4_4_lut_adj_530.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_531 (.I0(n16918), .I1(n17043), .I2(n10_adj_2288), 
            .I3(n17094), .O(n17109));   // coms.v(171[16:355])
    defparam i1_4_lut_adj_531.LUT_INIT = 16'h6996;
    SB_DFFESS \data_out_5[[4__2200  (.Q(\data_out[5] [4]), .C(CLK_c), .E(n10055), 
            .D(n2362[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_532 (.I0(\data_out_frame2[9] [3]), .I1(\data_out_frame2[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9901));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_532.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n10625));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n10624));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n10623));   // coms.v(426[12] 547[6])
    SB_LUT4 i5_4_lut_adj_533 (.I0(\data_out[5] [3]), .I1(n17055), .I2(n16990), 
            .I3(n17064), .O(n12_adj_2289));   // coms.v(171[16:355])
    defparam i5_4_lut_adj_533.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_534 (.I0(\data_out_frame2[7] [4]), .I1(\data_out_frame2[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9913));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_534.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_535 (.I0(\data_out_frame2[15] [3]), .I1(\data_out_frame2[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9916));   // coms.v(242[17:884])
    defparam i1_2_lut_adj_535.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n10622));   // coms.v(426[12] 547[6])
    SB_LUT4 i6_4_lut_adj_536 (.I0(n17109), .I1(n12_adj_2289), .I2(\data_out[6] [2]), 
            .I3(\data_out[9] [4]), .O(data_out_10__1__N_168));   // coms.v(171[16:355])
    defparam i6_4_lut_adj_536.LUT_INIT = 16'h6996;
    SB_LUT4 n18083_bdd_4_lut (.I0(n18083), .I1(n6_adj_2290), .I2(n17563), 
            .I3(byte_transmit_counter2[3]), .O(n18086));
    defparam n18083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n10621));   // coms.v(426[12] 547[6])
    SB_DFF \data_out_2[[5__2223  (.Q(\data_out[2][5] ), .C(CLK_c), .D(n10362));   // coms.v(280[12] 380[6])
    SB_LUT4 i2_3_lut_adj_537 (.I0(\data_out[6][0] ), .I1(data_out_7__2__N_447), 
            .I2(\data_out[7] [4]), .I3(GND_net), .O(n17064));   // coms.v(172[16:77])
    defparam i2_3_lut_adj_537.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut (.I0(data_out_6__1__N_537), .I1(\data_out[8][5] ), 
            .I2(\data_out[8][6] ), .I3(GND_net), .O(n9716));   // coms.v(181[17:93])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15411_2_lut_3_lut (.I0(n4445), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(GND_net), .O(n10259));
    defparam i15411_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 n18011_bdd_4_lut (.I0(n18011), .I1(n2_adj_2291), .I2(n17594), 
            .I3(\byte_transmit_counter[2] ), .O(n18014));
    defparam n18011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_538 (.I0(\data_out[5] [3]), .I1(\data_out[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9737));   // coms.v(115[16:67])
    defparam i1_2_lut_adj_538.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_539 (.I0(n9505), .I1(\data_out[9] [6]), .I2(\data_out[9][2] ), 
            .I3(GND_net), .O(n16978));   // coms.v(172[16:77])
    defparam i2_3_lut_adj_539.LUT_INIT = 16'h9696;
    SB_LUT4 i11_3_lut_adj_540 (.I0(n21_adj_2271), .I1(n19_adj_2270), .I2(n20_adj_2267), 
            .I3(GND_net), .O(n29));   // coms.v(272[12:25])
    defparam i11_3_lut_adj_540.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_541 (.I0(n9814), .I1(n9839), .I2(n9916), .I3(\data_out_frame2[5] [4]), 
            .O(n17040));   // coms.v(237[17:221])
    defparam i3_4_lut_adj_541.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_542 (.I0(\data_out_frame2[10] [6]), .I1(n9901), 
            .I2(n9919), .I3(n9589), .O(n10_adj_2292));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_542.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_543 (.I0(data_out_7__3__N_441), .I1(\data_out[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17076));   // coms.v(173[16:77])
    defparam i1_2_lut_adj_543.LUT_INIT = 16'h6666;
    SB_DFF \data_out_2[[7__2221  (.Q(\data_out[2][7] ), .C(CLK_c), .D(n10361));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_3[[0__2220  (.Q(\data_out[3][0] ), .C(CLK_c), .D(n10360));   // coms.v(280[12] 380[6])
    SB_LUT4 i2_3_lut_adj_544 (.I0(\data_out[7] [5]), .I1(\data_out[7] [6]), 
            .I2(\data_out[7] [7]), .I3(GND_net), .O(n9505));   // coms.v(172[16:77])
    defparam i2_3_lut_adj_544.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n10620));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_545 (.I0(\data_out[9] [7]), .I1(\data_out[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17007));   // coms.v(173[16:77])
    defparam i1_2_lut_adj_545.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n10619));   // coms.v(426[12] 547[6])
    SB_LUT4 i3_4_lut_adj_546 (.I0(\data_out[8] [0]), .I1(n17007), .I2(n9505), 
            .I3(n17076), .O(data_out_10__3__N_146));   // coms.v(173[16:77])
    defparam i3_4_lut_adj_546.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_547 (.I0(\data_out[6] [2]), .I1(\data_out[6][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n9783));   // coms.v(170[16:355])
    defparam i1_2_lut_adj_547.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_548 (.I0(n9678), .I1(n17016), .I2(n9671), .I3(n6_adj_2293), 
            .O(n16960));   // coms.v(229[16:299])
    defparam i4_4_lut_adj_548.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_549 (.I0(n16975), .I1(\data_out[7] [6]), .I2(n9509), 
            .I3(GND_net), .O(data_out_10__4__N_135));   // coms.v(174[16:77])
    defparam i2_3_lut_adj_549.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_550 (.I0(\data_out[7] [7]), .I1(\data_out[8] [1]), 
            .I2(\data_out[8] [0]), .I3(GND_net), .O(n9509));   // coms.v(174[16:77])
    defparam i2_3_lut_adj_550.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_551 (.I0(n9692), .I1(\data_out_frame2[6] [5]), 
            .I2(\data_out_frame2[13] [0]), .I3(n9749), .O(n28_adj_2294));   // coms.v(237[17:221])
    defparam i10_4_lut_adj_551.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(n17127), .I1(n28_adj_2294), .I2(n17133), .I3(GND_net), 
            .O(n32));   // coms.v(237[17:221])
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_552 (.I0(\data_out[9] [5]), .I1(n16990), .I2(GND_net), 
            .I3(GND_net), .O(n17070));   // coms.v(175[16:77])
    defparam i1_2_lut_adj_552.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_553 (.I0(n9737), .I1(data_out_6__1__N_537), .I2(\data_out[5] [1]), 
            .I3(\data_out[5] [2]), .O(n17025));   // coms.v(130[17:68])
    defparam i1_4_lut_adj_553.LUT_INIT = 16'h6996;
    SB_DFF \data_out_3[[2__2218  (.Q(\data_out[3][2] ), .C(CLK_c), .D(n10359));   // coms.v(280[12] 380[6])
    SB_LUT4 i3_4_lut_adj_554 (.I0(\data_out[10] [1]), .I1(\data_out[6] [3]), 
            .I2(\data_out[8]_c [2]), .I3(n17070), .O(data_out_10__5__N_124));   // coms.v(175[16:77])
    defparam i3_4_lut_adj_554.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_555 (.I0(n16960), .I1(n17034), .I2(n16972), 
            .I3(n17040), .O(n30_adj_2295));   // coms.v(237[17:221])
    defparam i12_4_lut_adj_555.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n17067), .I1(n17115), .I2(n17100), .I3(n17118), 
            .O(n31_c));   // coms.v(237[17:221])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_556 (.I0(\data_out[10] [2]), .I1(\data_out[9] [6]), 
            .I2(\data_out[6] [2]), .I3(n16998), .O(data_out_10__6__N_113));   // coms.v(176[16:77])
    defparam i3_4_lut_adj_556.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_557 (.I0(\data_out[8]_c [2]), .I1(\data_out[8]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28_adj_2287));   // coms.v(21[11:19])
    defparam i1_2_lut_adj_557.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_558 (.I0(\data_out[6] [3]), .I1(\data_out[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16918));   // coms.v(179[16:84])
    defparam i1_2_lut_adj_558.LUT_INIT = 16'h6666;
    SB_LUT4 i152_2_lut_4_lut (.I0(tx_transmit_N_1949[3]), .I1(n8938), .I2(tx_active), 
            .I3(r_SM_Main_2__N_2036[0]), .O(n456));   // coms.v(365[6] 377[9])
    defparam i152_2_lut_4_lut.LUT_INIT = 16'hfff1;
    SB_LUT4 i11_4_lut_adj_559 (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[5] [0]), 
            .I2(\data_out_frame2[6] [6]), .I3(\data_out_frame2[6] [2]), 
            .O(n29_adj_2296));   // coms.v(237[17:221])
    defparam i11_4_lut_adj_559.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n10618));   // coms.v(426[12] 547[6])
    SB_LUT4 i17_4_lut_adj_560 (.I0(n29_adj_2296), .I1(n31_c), .I2(n30_adj_2295), 
            .I3(n32), .O(n17135));   // coms.v(237[17:221])
    defparam i17_4_lut_adj_560.LUT_INIT = 16'h6996;
    SB_CARRY add_2495_13 (.CI(n15524), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n15525));
    SB_DFF delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .D(n10464));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_3[[4__2216  (.Q(\data_out[3][4] ), .C(CLK_c), .D(n10358));   // coms.v(280[12] 380[6])
    SB_LUT4 i3_4_lut_adj_561 (.I0(n32_adj_2297), .I1(\data_out[8][4] ), 
            .I2(\data_out[9] [7]), .I3(n17028), .O(data_out_10__7__N_101));   // coms.v(179[16:84])
    defparam i3_4_lut_adj_561.LUT_INIT = 16'h6996;
    SB_LUT4 i15337_2_lut (.I0(\data_out[0][5] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17589));
    defparam i15337_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_562 (.I0(\data_out_frame2[5] [2]), .I1(\data_out_frame2[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9886));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_562.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i2_3_lut (.I0(\data_out[2][5] ), 
            .I1(\data_out[3][5] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2298));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_563 (.I0(\data_out_frame2[15] [5]), .I1(\data_out_frame2[11] [0]), 
            .I2(\data_out_frame2[13] [6]), .I3(GND_net), .O(n16923));   // coms.v(233[16:291])
    defparam i2_3_lut_adj_563.LUT_INIT = 16'h9696;
    SB_DFF \data_out_3[[5__2215  (.Q(\data_out[3][5] ), .C(CLK_c), .D(n10357));   // coms.v(280[12] 380[6])
    SB_DFF \data_out_3[[6__2214  (.Q(\data_out[3] [6]), .C(CLK_c), .D(n10356));   // coms.v(280[12] 380[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n10617));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_564 (.I0(\data_out_frame2[12] [3]), .I1(\data_out_frame2[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9754));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_564.LUT_INIT = 16'h6666;
    SB_LUT4 i10601_2_lut (.I0(\rand_setpoint[30] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2292[0]));   // coms.v(283[4] 379[11])
    defparam i10601_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14792_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[0] ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_2036[0]), .I3(GND_net), .O(n17230));
    defparam i14792_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out[6] [5]), 
            .I1(\data_out[7] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2299));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut_adj_565 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state_c [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n8603));
    defparam i1_4_lut_4_lut_adj_565.LUT_INIT = 16'h0504;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15572 (.I0(byte_transmit_counter[1]), 
            .I1(n17555), .I2(n5_adj_2300), .I3(\byte_transmit_counter[2] ), 
            .O(n18035));
    defparam byte_transmit_counter_1__bdd_4_lut_15572.LUT_INIT = 16'he4aa;
    SB_LUT4 i15345_2_lut (.I0(\data_out[5] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17548));
    defparam i15345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_3_lut_4_lut_adj_566 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[2] [7]), .O(n22_adj_2301));
    defparam i6_3_lut_4_lut_adj_566.LUT_INIT = 16'h9f6f;
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n10616));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n10615));   // coms.v(426[12] 547[6])
    SB_LUT4 i2_3_lut_adj_567 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // coms.v(450[7:23])
    defparam i2_3_lut_adj_567.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out[6] [2]), 
            .I1(\data_out[7] [2]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2208));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n10614));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n10613));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n10612));   // coms.v(426[12] 547[6])
    SB_DFFE delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(VCC_net), 
            .D(n10851));   // coms.v(280[12] 380[6])
    SB_LUT4 i8_4_lut_adj_568 (.I0(\data_out_frame2[7] [2]), .I1(n16923), 
            .I2(n16915), .I3(n16933), .O(n20_adj_2302));   // coms.v(230[16:237])
    defparam i8_4_lut_adj_568.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n10611));   // coms.v(426[12] 547[6])
    SB_LUT4 i7_4_lut_adj_569 (.I0(n9749), .I1(\data_out_frame2[12] [0]), 
            .I2(\data_out_frame2[16] [5]), .I3(\data_out_frame2[5] [1]), 
            .O(n19_adj_2303));   // coms.v(230[16:237])
    defparam i7_4_lut_adj_569.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_570 (.I0(n16957), .I1(n17061), .I2(n17049), .I3(n17106), 
            .O(n21_adj_2304));   // coms.v(230[16:237])
    defparam i9_4_lut_adj_570.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i1_3_lut (.I0(\data_out[0] [6]), 
            .I1(\data_out[1][6] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n1_c));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_adj_571 (.I0(n21_adj_2304), .I1(n19_adj_2303), .I2(n20_adj_2302), 
            .I3(GND_net), .O(n17107));   // coms.v(230[16:237])
    defparam i11_3_lut_adj_571.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_572 (.I0(\data_out_frame2[16] [4]), .I1(\data_out_frame2[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9810));   // coms.v(240[17:239])
    defparam i1_2_lut_adj_572.LUT_INIT = 16'h6666;
    SB_LUT4 i15297_2_lut (.I0(\data_out[3] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17588));
    defparam i15297_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10596_2_lut (.I0(\rand_setpoint[29] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2327[0]));   // coms.v(283[4] 379[11])
    defparam i10596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15370_2_lut (.I0(\data_out[5] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17543));
    defparam i15370_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_573 (.I0(\data_out_frame2[9] [6]), .I1(\data_out_frame2[6] [0]), 
            .I2(n9826), .I3(GND_net), .O(n17100));   // coms.v(241[17:248])
    defparam i1_2_lut_3_lut_adj_573.LUT_INIT = 16'h9696;
    SB_DFF \data_out_3[[7__2213  (.Q(\data_out[3][7] ), .C(CLK_c), .D(n10355));   // coms.v(280[12] 380[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut (.I0(\data_out_frame2[14] [4]), 
            .I1(\data_out_frame2[15] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n12_adj_2305));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut (.I0(\data_out_frame2[12] [4]), 
            .I1(\data_out_frame2[13] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n11));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_574 (.I0(\data_out_frame2[10] [5]), .I1(\data_out_frame2[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9763));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_574.LUT_INIT = 16'h6666;
    SB_LUT4 i14798_2_lut (.I0(delay_counter[8]), .I1(delay_counter[13]), 
            .I2(GND_net), .I3(GND_net), .O(n17236));
    defparam i14798_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_575 (.I0(\data_out_frame2[9] [0]), .I1(\data_out_frame2[15] [4]), 
            .I2(\data_out_frame2[8] [4]), .I3(GND_net), .O(n9749));   // coms.v(241[17:248])
    defparam i2_3_lut_adj_575.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_576 (.I0(n9749), .I1(n9865), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_2306));   // coms.v(240[17:239])
    defparam i1_2_lut_adj_576.LUT_INIT = 16'h6666;
    SB_LUT4 i12728_3_lut (.I0(delay_counter[0]), .I1(n17637), .I2(n1419), 
            .I3(GND_net), .O(n10851));
    defparam i12728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14838_4_lut (.I0(delay_counter[7]), .I1(n12993), .I2(delay_counter[5]), 
            .I3(delay_counter[12]), .O(n17276));
    defparam i14838_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_577 (.I0(\data_out_frame2[13] [5]), .I1(n9843), 
            .I2(\data_out_frame2[10] [7]), .I3(n6_adj_2306), .O(n16987));   // coms.v(240[17:239])
    defparam i4_4_lut_adj_577.LUT_INIT = 16'h6996;
    SB_LUT4 n17987_bdd_4_lut_4_lut (.I0(byte_transmit_counter2[0]), .I1(\data_out_frame2[0] [4]), 
            .I2(byte_transmit_counter2[2]), .I3(n17987), .O(n17990));
    defparam n17987_bdd_4_lut_4_lut.LUT_INIT = 16'hfa04;
    SB_LUT4 i14840_4_lut (.I0(delay_counter[0]), .I1(n12991), .I2(delay_counter[14]), 
            .I3(n13298), .O(n17278));
    defparam i14840_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_578 (.I0(\data_out_frame2[13] [1]), .I1(\data_out_frame2[16] [7]), 
            .I2(\data_out_frame2[15] [7]), .I3(GND_net), .O(n9910));   // coms.v(227[16:31])
    defparam i1_2_lut_3_lut_adj_578.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[10] [1]), 
            .I2(\data_out_frame2[9] [7]), .I3(\data_out_frame2[9] [5]), 
            .O(n17034));   // coms.v(232[16:229])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_579 (.I0(n9579), .I1(\data_out_frame2[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_2307));   // coms.v(240[17:239])
    defparam i2_2_lut_adj_579.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_580 (.I0(\data_out_frame2[12] [4]), .I1(n17067), 
            .I2(n16987), .I3(n17112), .O(n14_adj_2308));   // coms.v(240[17:239])
    defparam i6_4_lut_adj_580.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15543 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [6]), .I2(\data_out_frame2[19] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n17999));
    defparam byte_transmit_counter2_0__bdd_4_lut_15543.LUT_INIT = 16'he4aa;
    SB_LUT4 i10_4_lut_adj_581 (.I0(delay_counter[2]), .I1(n42_adj_2165), 
            .I2(delay_counter[4]), .I3(n17236), .O(n23_adj_2309));
    defparam i10_4_lut_adj_581.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_582 (.I0(n23_adj_2309), .I1(n17230), .I2(n17278), 
            .I3(n17276), .O(n16839));
    defparam i1_4_lut_adj_582.LUT_INIT = 16'h0002;
    SB_LUT4 i8020_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n10380));
    defparam i8020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8021_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n10381));
    defparam i8021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_583 (.I0(\data_out_frame2[10] [1]), .I1(n14_adj_2308), 
            .I2(n10_adj_2307), .I3(n9763), .O(n17113));   // coms.v(240[17:239])
    defparam i7_4_lut_adj_583.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter2_1__bdd_4_lut_15528 (.I0(byte_transmit_counter2[1]), 
            .I1(n11), .I2(n12_adj_2305), .I3(byte_transmit_counter2[2]), 
            .O(n17897));
    defparam byte_transmit_counter2_1__bdd_4_lut_15528.LUT_INIT = 16'he4aa;
    SB_DFFESS \data_out_5[[5__2199  (.Q(\data_out[5] [5]), .C(CLK_c), .E(n10055), 
            .D(n2327[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 n18035_bdd_4_lut (.I0(n18035), .I1(n17588), .I2(n1_c), .I3(\byte_transmit_counter[2] ), 
            .O(n18038));
    defparam n18035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n10610));   // coms.v(426[12] 547[6])
    SB_LUT4 i8024_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n10384));
    defparam i8024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15567 (.I0(byte_transmit_counter[1]), 
            .I1(n17548), .I2(n5_adj_2299), .I3(\byte_transmit_counter[2] ), 
            .O(n18029));
    defparam byte_transmit_counter_1__bdd_4_lut_15567.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_664_i1_4_lut (.I0(n17445), .I1(\rand_setpoint[9] ), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n1916[0]));   // coms.v(283[4] 379[11])
    defparam mux_664_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i142_2_lut_4_lut (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(n9357), .I3(n445), .O(n446));   // coms.v(302[6] 314[9])
    defparam i142_2_lut_4_lut.LUT_INIT = 16'hff07;
    SB_LUT4 i8025_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n10385));
    defparam i8025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11084_2_lut (.I0(tx_transmit_N_1949[3]), .I1(n8938), .I2(GND_net), 
            .I3(GND_net), .O(n9357));
    defparam i11084_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15324_2_lut_3_lut (.I0(\data_out_frame2[0] [2]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17578));
    defparam i15324_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i15206_2_lut (.I0(\rand_setpoint[10] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17450));   // coms.v(283[4] 379[11])
    defparam i15206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_584 (.I0(\data_out_frame2[7] [0]), .I1(\data_out_frame2[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17097));   // coms.v(228[16:596])
    defparam i1_2_lut_adj_584.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_585 (.I0(n13272), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [3]), .O(n16891));
    defparam i1_2_lut_4_lut_adj_585.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_586 (.I0(\data_out_frame2[10] [6]), .I1(\data_out_frame2[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16933));   // coms.v(239[17:230])
    defparam i1_2_lut_adj_586.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_587 (.I0(byte_transmit_counter[0]), .I1(tx_transmit_N_1949[0]), 
            .I2(n10181), .I3(n16839), .O(n16247));   // coms.v(19[11:32])
    defparam i12_4_lut_adj_587.LUT_INIT = 16'h0aca;
    SB_LUT4 i8022_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n10382));
    defparam i8022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_588 (.I0(\data_out_frame2[5] [0]), .I1(\data_out_frame2[8] [3]), 
            .I2(\data_out_frame2[15] [3]), .I3(\data_out_frame2[5] [1]), 
            .O(n9865));   // coms.v(239[17:230])
    defparam i3_4_lut_adj_588.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_589 (.I0(\data_out_frame2[15] [2]), .I1(\data_out_frame2[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9814));   // coms.v(231[16:291])
    defparam i1_2_lut_adj_589.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_590 (.I0(\data_out_frame2[16] [2]), .I1(\data_out_frame2[14] [4]), 
            .I2(n9814), .I3(n9865), .O(n16_adj_2312));   // coms.v(239[17:230])
    defparam i6_4_lut_adj_590.LUT_INIT = 16'h6996;
    SB_LUT4 add_2494_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n15659), .O(tx_transmit_N_1949[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2494_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n15658), .O(tx_transmit_N_1949[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2494_8 (.CI(n15658), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n15659));
    SB_LUT4 add_2494_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n15657), .O(tx_transmit_N_1949[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2494_7 (.CI(n15657), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n15658));
    SB_LUT4 i8026_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n10386));
    defparam i8026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_2494_6_lut (.I0(GND_net), .I1(\byte_transmit_counter[4] ), 
            .I2(GND_net), .I3(n15656), .O(tx_transmit_N_1949[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 select_238_Select_7_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_2250));
    defparam select_238_Select_7_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_6_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_2253));
    defparam select_238_Select_6_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFFESS \data_out_5[[6__2198  (.Q(data_out_7__2__N_447), .C(CLK_c), 
            .E(n10055), .D(n2292[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_CARRY add_2494_6 (.CI(n15656), .I0(\byte_transmit_counter[4] ), .I1(GND_net), 
            .CO(n15657));
    SB_LUT4 i7_4_lut_adj_591 (.I0(\data_out_frame2[11] [6]), .I1(n17037), 
            .I2(n16933), .I3(n17088), .O(n17_adj_2313));   // coms.v(239[17:230])
    defparam i7_4_lut_adj_591.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_592 (.I0(n17_adj_2313), .I1(n17097), .I2(n16_adj_2312), 
            .I3(n17112), .O(n17114));   // coms.v(239[17:230])
    defparam i9_4_lut_adj_592.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out[6] [6]), 
            .I1(\data_out[7] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2300));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2494_5_lut (.I0(GND_net), .I1(\byte_transmit_counter[3] ), 
            .I2(GND_net), .I3(n15655), .O(tx_transmit_N_1949[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_593 (.I0(\data_out_frame2[16] [2]), .I1(\data_out_frame2[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9839));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_593.LUT_INIT = 16'h6666;
    SB_CARRY add_2494_5 (.CI(n15655), .I0(\byte_transmit_counter[3] ), .I1(GND_net), 
            .CO(n15656));
    SB_LUT4 select_238_Select_8_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_2249));
    defparam select_238_Select_8_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_2494_4_lut (.I0(GND_net), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n15654), .O(tx_transmit_N_1949[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_594 (.I0(\data_out_frame2[12] [2]), .I1(\data_out_frame2[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9671));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_594.LUT_INIT = 16'h6666;
    SB_LUT4 i15362_2_lut (.I0(data_out_7__2__N_447), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17555));
    defparam i15362_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_595 (.I0(\data_out_frame2[8] [2]), .I1(\data_out_frame2[6] [3]), 
            .I2(\data_out_frame2[10] [5]), .I3(GND_net), .O(n17118));   // coms.v(238[17:230])
    defparam i1_2_lut_3_lut_adj_595.LUT_INIT = 16'h9696;
    SB_LUT4 i10568_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [0]), .O(\FRAME_MATCHER.i_31__N_1312 [0]));
    defparam i10568_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_596 (.I0(\data_out_frame2[8] [2]), .I1(\data_out_frame2[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9758));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_596.LUT_INIT = 16'h6666;
    SB_LUT4 i10733_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [31]), .O(\FRAME_MATCHER.i_31__N_1312 [31]));
    defparam i10733_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_9_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_2248));
    defparam select_238_Select_9_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_adj_597 (.I0(\data_out_frame2[16] [1]), .I1(\data_out_frame2[13] [3]), 
            .I2(\data_out_frame2[15] [2]), .I3(GND_net), .O(n17082));   // coms.v(238[17:230])
    defparam i2_3_lut_adj_597.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_598 (.I0(\data_out_frame2[12] [1]), .I1(\data_out_frame2[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16915));   // coms.v(238[17:230])
    defparam i1_2_lut_adj_598.LUT_INIT = 16'h6666;
    SB_LUT4 select_238_Select_10_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_2247));
    defparam select_238_Select_10_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10736_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [30]), .O(\FRAME_MATCHER.i_31__N_1312 [30]));
    defparam i10736_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10741_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [29]), .O(\FRAME_MATCHER.i_31__N_1312 [29]));
    defparam i10741_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_11_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_2246));
    defparam select_238_Select_11_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10742_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [28]), .O(\FRAME_MATCHER.i_31__N_1312 [28]));
    defparam i10742_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_4_lut_adj_599 (.I0(n16915), .I1(n17082), .I2(n17019), 
            .I3(n17118), .O(n26_adj_2314));   // coms.v(238[17:230])
    defparam i11_4_lut_adj_599.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_600 (.I0(\data_out_frame2[10] [3]), .I1(\data_out_frame2[12] [3]), 
            .I2(\data_out_frame2[8] [5]), .I3(\data_out_frame2[16] [7]), 
            .O(n24_adj_2315));   // coms.v(238[17:230])
    defparam i9_4_lut_adj_600.LUT_INIT = 16'h6996;
    SB_LUT4 i10743_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [27]), .O(\FRAME_MATCHER.i_31__N_1312 [27]));
    defparam i10743_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_601 (.I0(n9671), .I1(n9839), .I2(\data_out_frame2[9] [7]), 
            .I3(\data_out_frame2[6] [7]), .O(n25_adj_2316));   // coms.v(238[17:230])
    defparam i10_4_lut_adj_601.LUT_INIT = 16'h6996;
    SB_LUT4 i8027_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n10387));
    defparam i8027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10744_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [26]), .O(\FRAME_MATCHER.i_31__N_1312 [26]));
    defparam i10744_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10745_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [25]), .O(\FRAME_MATCHER.i_31__N_1312 [25]));
    defparam i10745_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6319_2_lut (.I0(byte_transmit_counter2[0]), .I1(byte_transmit_counter2[1]), 
            .I2(GND_net), .I3(GND_net), .O(n8621));   // coms.v(413[36:58])
    defparam i6319_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame2[6] [2]), 
            .I1(\data_out_frame2[7] [2]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2317));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_602 (.I0(n23_adj_2318), .I1(n25_adj_2316), .I2(n24_adj_2315), 
            .I3(n26_adj_2314), .O(n17132));   // coms.v(238[17:230])
    defparam i14_4_lut_adj_602.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame2[5] [2]), 
            .I1(n5_adj_2317), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2201));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 select_238_Select_12_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_2245));
    defparam select_238_Select_12_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_603 (.I0(\data_out_frame2[11] [4]), .I1(\data_out_frame2[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9892));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_603.LUT_INIT = 16'h6666;
    SB_LUT4 i15336_3_lut_4_lut (.I0(\data_out[5] [5]), .I1(n17025), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(data_out_7__2__N_447), .O(n17445));   // coms.v(283[4] 379[11])
    defparam i15336_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i10746_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [24]), .O(\FRAME_MATCHER.i_31__N_1312 [24]));
    defparam i10746_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10747_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [23]), .O(\FRAME_MATCHER.i_31__N_1312 [23]));
    defparam i10747_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10748_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [22]), .O(\FRAME_MATCHER.i_31__N_1312 [22]));
    defparam i10748_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_2494_4 (.CI(n15654), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n15655));
    SB_LUT4 add_2494_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n15653), .O(tx_transmit_N_1949[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 select_238_Select_13_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_2244));
    defparam select_238_Select_13_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out[6] [7]), 
            .I1(\data_out[7] [7]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2188));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8028_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n10388));
    defparam i8028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_238_Select_14_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_2243));
    defparam select_238_Select_14_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_15_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_2242));
    defparam select_238_Select_15_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_16_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_2241));
    defparam select_238_Select_16_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_17_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_2240));
    defparam select_238_Select_17_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_604 (.I0(tx_transmit_N_1949[0]), .I1(tx_transmit_N_1949[1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2311));
    defparam i1_2_lut_adj_604.LUT_INIT = 16'h8888;
    SB_CARRY add_2494_3 (.CI(n15653), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n15654));
    SB_LUT4 add_2494_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(n65), .I3(GND_net), .O(tx_transmit_N_1949[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2494_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2494_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(n65), 
            .CO(n15653));
    SB_LUT4 i1_2_lut_adj_605 (.I0(\data_out_frame2[10] [0]), .I1(\data_out_frame2[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n9707));   // coms.v(239[17:230])
    defparam i1_2_lut_adj_605.LUT_INIT = 16'h6666;
    SB_LUT4 select_238_Select_18_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_2239));
    defparam select_238_Select_18_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_997_33_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [31]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17889), .I3(n15652), .O(\FRAME_MATCHER.i_31__N_1280 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_33_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut_adj_606 (.I0(\data_out_frame2[12] [3]), .I1(\data_out_frame2[12] [2]), 
            .I2(\data_out_frame2[11] [7]), .I3(n16963), .O(n9579));   // coms.v(227[16:31])
    defparam i3_4_lut_adj_606.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_607 (.I0(n9579), .I1(n9707), .I2(\data_out_frame2[10] [4]), 
            .I3(GND_net), .O(n17088));   // coms.v(239[17:230])
    defparam i2_3_lut_adj_607.LUT_INIT = 16'h9696;
    SB_LUT4 i10749_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [21]), .O(\FRAME_MATCHER.i_31__N_1312 [21]));
    defparam i10749_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10750_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [20]), .O(\FRAME_MATCHER.i_31__N_1312 [20]));
    defparam i10750_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 n18029_bdd_4_lut (.I0(n18029), .I1(n2_adj_2298), .I2(n17589), 
            .I3(\byte_transmit_counter[2] ), .O(n18032));
    defparam n18029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_608 (.I0(\data_out_frame2[13] [2]), .I1(\data_out_frame2[16] [0]), 
            .I2(\data_out_frame2[16] [6]), .I3(\data_out_frame2[15] [0]), 
            .O(n17016));   // coms.v(237[17:221])
    defparam i2_4_lut_adj_608.LUT_INIT = 16'h6996;
    SB_LUT4 add_997_32_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [30]), .I1(\FRAME_MATCHER.i [30]), 
            .I2(n17889), .I3(n15651), .O(\FRAME_MATCHER.i_31__N_1280 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_32_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15347_2_lut (.I0(\data_out[1] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17594));
    defparam i15347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_609 (.I0(\data_out_frame2[6] [6]), .I1(\data_out_frame2[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9776));   // coms.v(237[17:221])
    defparam i1_2_lut_adj_609.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i2_3_lut (.I0(\data_out[2][2] ), 
            .I1(\data_out[3][2] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2291));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_2_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_997_32 (.CI(n15651), .I0(\FRAME_MATCHER.i [30]), .I1(n17889), 
            .CO(n15652));
    SB_LUT4 add_2495_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n15523), .O(n6517[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_997_31_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [29]), .I1(\FRAME_MATCHER.i [29]), 
            .I2(n17889), .I3(n15650), .O(\FRAME_MATCHER.i_31__N_1280 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_31_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_31 (.CI(n15650), .I0(\FRAME_MATCHER.i [29]), .I1(n17889), 
            .CO(n15651));
    SB_DFFE \data_out_10[[7__2157  (.Q(\data_out[10] [7]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__7__N_101));   // coms.v(280[12] 380[6])
    SB_LUT4 add_997_30_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [28]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(n17889), .I3(n15649), .O(\FRAME_MATCHER.i_31__N_1280 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_30_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15281_2_lut (.I0(data_out_7__3__N_441), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17569));
    defparam i15281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10751_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [19]), .O(\FRAME_MATCHER.i_31__N_1312 [19]));
    defparam i10751_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15284_3_lut (.I0(\data_out_frame2[0] [3]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17576));
    defparam i15284_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 select_238_Select_19_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_2237));
    defparam select_238_Select_19_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFFE \data_out_10[[6__2158  (.Q(\data_out[10] [6]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__6__N_113));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_10[[5__2159  (.Q(\data_out[10] [5]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__5__N_124));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_10[[4__2160  (.Q(\data_out[10] [4]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__4__N_135));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_10[[3__2161  (.Q(\data_out[10] [3]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__3__N_146));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_10[[2__2162  (.Q(\data_out[10] [2]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__2__N_157));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_10[[1__2163  (.Q(\data_out[10] [1]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__1__N_168));   // coms.v(280[12] 380[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n10609));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_10[[0__2164  (.Q(\data_out[10] [0]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_10__0__N_219));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_9[[7__2165  (.Q(\data_out[9] [7]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__7__N_272));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_9[[6__2166  (.Q(\data_out[9] [6]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__6__N_324));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_9[[5__2167  (.Q(\data_out[9] [5]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__5__N_334));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_9[[4__2168  (.Q(\data_out[9] [4]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__4__N_345));   // coms.v(280[12] 380[6])
    SB_DFFE \data_out_9[[3__2169  (.Q(\data_out[9] [3]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__3__N_356));   // coms.v(280[12] 380[6])
    SB_LUT4 i10752_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [18]), .O(\FRAME_MATCHER.i_31__N_1312 [18]));
    defparam i10752_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10753_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [17]), .O(\FRAME_MATCHER.i_31__N_1312 [17]));
    defparam i10753_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFFE \data_out_9[[1__2171  (.Q(\data_out[9] [1]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__1__N_378));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_610 (.I0(tx_transmit_N_1949[7]), .I1(tx_transmit_N_1949[5]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_2319));   // coms.v(336[10:53])
    defparam i1_2_lut_adj_610.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_611 (.I0(n9776), .I1(\data_out_frame2[6] [2]), 
            .I2(\data_out_frame2[14] [2]), .I3(n17016), .O(n15_adj_2320));   // coms.v(237[17:221])
    defparam i6_4_lut_adj_611.LUT_INIT = 16'h6996;
    SB_LUT4 i10754_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [16]), .O(\FRAME_MATCHER.i_31__N_1312 [16]));
    defparam i10754_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15313_3_lut (.I0(\data_out_frame2[0] [6]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17563));
    defparam i15313_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 select_238_Select_20_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_2235));
    defparam select_238_Select_20_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n10608));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_9[[0__2172  (.Q(\data_out[9] [0]), .C(CLK_c), .E(data_out_10__7__N_110), 
            .D(data_out_9__0__N_389));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i1 (.Q(\data_out_frame2[0] [0]), .C(CLK_c), 
           .D(n17354));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame2[6] [6]), 
            .I1(\data_out_frame2[7] [6]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2321));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame2[6] [3]), 
            .I1(\data_out_frame2[7] [3]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2322));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame2[5] [3]), 
            .I1(n5_adj_2322), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2187));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_out_frame2_0___i140 (.Q(\data_out_frame2[17] [3]), .C(CLK_c), 
           .D(n10824));   // coms.v(426[12] 547[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut (.I0(\data_out_frame2[5] [6]), 
            .I1(n5_adj_2321), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2290));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_CARRY add_997_30 (.CI(n15649), .I0(\FRAME_MATCHER.i [28]), .I1(n17889), 
            .CO(n15650));
    SB_DFF data_out_frame2_0___i139 (.Q(\data_out_frame2[17] [2]), .C(CLK_c), 
           .D(n10823));   // coms.v(426[12] 547[6])
    SB_LUT4 i8_4_lut_adj_612 (.I0(n15_adj_2320), .I1(n17079), .I2(n14_adj_2323), 
            .I3(n17088), .O(n17131));   // coms.v(237[17:221])
    defparam i8_4_lut_adj_612.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n10604));   // coms.v(426[12] 547[6])
    SB_LUT4 mux_638_i1_4_lut (.I0(data_out_7__2__N_447), .I1(n17450), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1881[0]));   // coms.v(283[4] 379[11])
    defparam mux_638_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_2_lut_adj_613 (.I0(\data_out_frame2[9] [7]), .I1(\data_out_frame2[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16926));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_613.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n10603));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n10602));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n10601));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n10600));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n10599));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n10598));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n10597));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n10596));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n10592));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_21_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_2233));
    defparam select_238_Select_21_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n10591));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n10590));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n10589));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n10588));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n10584));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n10583));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n10582));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n10577));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n10576));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n10575));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n10574));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(CLK_c), 
            .D(n16383), .S(n16377));   // coms.v(426[12] 547[6])
    SB_DFF \UART_TRANSMITTER.state_i0_i0  (.Q(\UART_TRANSMITTER.state[0] ), 
           .C(CLK_c), .D(n16259));   // coms.v(280[12] 380[6])
    SB_LUT4 add_997_29_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [27]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(n17889), .I3(n15648), .O(\FRAME_MATCHER.i_31__N_1280 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_29_lut.LUT_INIT = 16'hA3AC;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(CLK_c), 
            .D(n16385), .S(n16379));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(CLK_c), 
            .D(n16387), .S(n16381));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(CLK_c), 
            .D(n16389), .S(n16353));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(CLK_c), 
            .D(n16391), .S(n16355));   // coms.v(426[12] 547[6])
    SB_LUT4 select_238_Select_22_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_2231));
    defparam select_238_Select_22_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_614 (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9895));   // coms.v(234[16:291])
    defparam i1_2_lut_adj_614.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(CLK_c), 
            .D(n16393), .S(n16357));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(CLK_c), 
            .D(n16395), .S(n16359));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(CLK_c), 
            .D(n16397), .S(n16361));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_615 (.I0(\data_out_frame2[16] [5]), .I1(n17034), 
            .I2(GND_net), .I3(GND_net), .O(n9688));   // coms.v(232[16:229])
    defparam i1_2_lut_adj_615.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(CLK_c), 
            .D(n16399), .S(n16363));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(CLK_c), 
            .D(n16401), .S(n16365));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(CLK_c), 
            .D(n16403), .S(n16367));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(CLK_c), 
            .D(n16405), .S(n16369));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(CLK_c), 
            .D(n16407), .S(n16371));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(CLK_c), 
            .D(n16409), .S(n16343));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(CLK_c), 
            .D(n16411), .S(n16345));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(CLK_c), 
            .D(n16413), .S(n16347));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(CLK_c), 
            .D(n16415), .S(n16349));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(CLK_c), 
            .D(n16417), .S(n16351));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(CLK_c), 
            .D(n16419), .S(n16447));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(CLK_c), 
            .D(n16421), .S(n16449));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(CLK_c), 
            .D(n16423), .S(n16451));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(CLK_c), 
            .D(n16425), .S(n16453));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(CLK_c), 
            .D(n16427), .S(n16455));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(CLK_c), 
            .D(n16429), .S(n16445));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(CLK_c), 
            .D(n16431), .S(n16443));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(CLK_c), 
            .D(n16433), .S(n16441));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(CLK_c), 
            .D(n16435), .S(n16335));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(CLK_c), 
            .D(n16437), .S(n16339));   // coms.v(426[12] 547[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state_c [3]), .C(CLK_c), 
            .D(n16439), .S(n16331));   // coms.v(426[12] 547[6])
    SB_DFFESS \data_out_5[[7__2197  (.Q(data_out_7__3__N_441), .C(CLK_c), 
            .E(n10055), .D(n2257[0]), .S(n10259));   // coms.v(280[12] 380[6])
    SB_LUT4 select_238_Select_23_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_2229));
    defparam select_238_Select_23_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10755_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [15]), .O(\FRAME_MATCHER.i_31__N_1312 [15]));
    defparam i10755_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15216_3_lut (.I0(n17254), .I1(n445), .I2(n8938), .I3(GND_net), 
            .O(n17460));
    defparam i15216_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i43_4_lut (.I0(n446), .I1(n17460), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(\UART_TRANSMITTER.state[1] ), .O(n25_adj_2324));
    defparam i43_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_3_lut_adj_616 (.I0(n10181), .I1(n25_adj_2324), .I2(\UART_TRANSMITTER.state[0] ), 
            .I3(GND_net), .O(n1419));
    defparam i1_3_lut_adj_616.LUT_INIT = 16'h5d5d;
    SB_LUT4 select_238_Select_24_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_2227));
    defparam select_238_Select_24_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_617 (.I0(\data_out_frame2[6] [1]), .I1(n9695), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2325));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_617.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_618 (.I0(\data_out_frame2[16] [0]), .I1(\data_out_frame2[12] [1]), 
            .I2(n9688), .I3(n6_adj_2325), .O(n17010));   // coms.v(227[16:31])
    defparam i4_4_lut_adj_618.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_619 (.I0(\data_out_frame2[16] [7]), .I1(\data_out_frame2[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16940));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_619.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_620 (.I0(\data_out_frame2[16] [4]), .I1(\data_out_frame2[12] [6]), 
            .I2(\data_out_frame2[5] [2]), .I3(GND_net), .O(n17067));   // coms.v(240[17:239])
    defparam i1_2_lut_3_lut_adj_620.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_621 (.I0(\data_out_frame2[6] [5]), .I1(\data_out_frame2[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9843));   // coms.v(240[17:239])
    defparam i1_2_lut_adj_621.LUT_INIT = 16'h6666;
    SB_LUT4 select_238_Select_25_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_2225));
    defparam select_238_Select_25_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_out_frame2_0___i138 (.Q(\data_out_frame2[17] [1]), .C(CLK_c), 
           .D(n10822));   // coms.v(426[12] 547[6])
    SB_CARRY add_997_29 (.CI(n15648), .I0(\FRAME_MATCHER.i [27]), .I1(n17889), 
            .CO(n15649));
    SB_LUT4 i10756_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [14]), .O(\FRAME_MATCHER.i_31__N_1312 [14]));
    defparam i10756_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_26_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_2223));
    defparam select_238_Select_26_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15208_2_lut (.I0(\rand_setpoint[11] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17456));   // coms.v(283[4] 379[11])
    defparam i15208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15562 (.I0(byte_transmit_counter[1]), 
            .I1(n17547), .I2(n5_adj_2326), .I3(\byte_transmit_counter[2] ), 
            .O(n18023));
    defparam byte_transmit_counter_1__bdd_4_lut_15562.LUT_INIT = 16'he4aa;
    SB_CARRY add_2495_12 (.CI(n15523), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n15524));
    SB_LUT4 i10757_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [13]), .O(\FRAME_MATCHER.i_31__N_1312 [13]));
    defparam i10757_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_622 (.I0(\data_out_frame2[0] [7]), .I1(n9843), 
            .I2(n9910), .I3(n9826), .O(n16_adj_2327));   // coms.v(227[16:31])
    defparam i6_4_lut_adj_622.LUT_INIT = 16'h6996;
    SB_LUT4 i12714_3_lut (.I0(delay_counter[14]), .I1(n17635), .I2(n1419), 
            .I3(GND_net), .O(n10858));
    defparam i12714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 select_238_Select_27_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_2221));
    defparam select_238_Select_27_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10758_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [12]), .O(\FRAME_MATCHER.i_31__N_1312 [12]));
    defparam i10758_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_28_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_2219));
    defparam select_238_Select_28_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7_4_lut_adj_623 (.I0(\data_out_frame2[8] [4]), .I1(\data_out_frame2[8] [0]), 
            .I2(\data_out_frame2[14] [1]), .I3(\data_out_frame2[15] [0]), 
            .O(n17_adj_2328));   // coms.v(227[16:31])
    defparam i7_4_lut_adj_623.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_624 (.I0(\data_out_frame2[12] [6]), .I1(\data_out_frame2[12] [2]), 
            .I2(\data_out_frame2[5] [2]), .I3(\data_out_frame2[10] [4]), 
            .O(n16957));   // coms.v(228[16:596])
    defparam i2_3_lut_4_lut_adj_624.LUT_INIT = 16'h6996;
    SB_LUT4 add_997_28_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [26]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(n17889), .I3(n15647), .O(\FRAME_MATCHER.i_31__N_1280 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_28_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i9_4_lut_adj_625 (.I0(n17_adj_2328), .I1(\data_out_frame2[12] [2]), 
            .I2(n16_adj_2327), .I3(n17010), .O(n17011));   // coms.v(227[16:31])
    defparam i9_4_lut_adj_625.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_626 (.I0(\data_out_frame2[12] [5]), .I1(\data_out_frame2[12] [7]), 
            .I2(\data_out_frame2[12] [3]), .I3(\data_out_frame2[5] [3]), 
            .O(n17061));   // coms.v(227[16:31])
    defparam i2_3_lut_4_lut_adj_626.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_627 (.I0(n13272), .I1(\FRAME_MATCHER.i [0]), .I2(n10_adj_2329), 
            .I3(GND_net), .O(n16895));
    defparam i1_3_lut_adj_627.LUT_INIT = 16'hfdfd;
    SB_LUT4 select_238_Select_29_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_2217));
    defparam select_238_Select_29_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_adj_628 (.I0(\data_out_frame2[7] [7]), .I1(\data_out_frame2[14] [7]), 
            .I2(\data_out_frame2[8] [3]), .I3(GND_net), .O(n9826));   // coms.v(227[16:31])
    defparam i2_3_lut_adj_628.LUT_INIT = 16'h9696;
    SB_LUT4 select_238_Select_30_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_2215));
    defparam select_238_Select_30_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_4_lut_adj_629 (.I0(\data_out_frame2[16] [4]), .I1(\data_out_frame2[9] [1]), 
            .I2(\data_out_frame2[6] [6]), .I3(\data_out_frame2[8] [5]), 
            .O(n17049));   // coms.v(230[16:237])
    defparam i2_3_lut_4_lut_adj_629.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_630 (.I0(\data_out_frame2[9] [6]), .I1(\data_out_frame2[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9859));   // coms.v(235[16:291])
    defparam i1_2_lut_adj_630.LUT_INIT = 16'h6666;
    SB_LUT4 mux_612_i1_4_lut (.I0(data_out_7__3__N_441), .I1(n17456), .I2(\UART_TRANSMITTER.state[1] ), 
            .I3(\UART_TRANSMITTER.state[2] ), .O(n1846[0]));   // coms.v(283[4] 379[11])
    defparam mux_612_i1_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 select_238_Select_31_i3_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n7212), 
            .I2(n1439), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_2210));
    defparam select_238_Select_31_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10759_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [11]), .O(\FRAME_MATCHER.i_31__N_1312 [11]));
    defparam i10759_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8029_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n10389));
    defparam i8029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_631 (.I0(\data_out_frame2[0] [6]), .I1(\data_out_frame2[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9589));
    defparam i1_2_lut_adj_631.LUT_INIT = 16'h6666;
    SB_LUT4 i10760_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [10]), .O(\FRAME_MATCHER.i_31__N_1312 [10]));
    defparam i10760_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11148_2_lut_3_lut (.I0(n62), .I1(n13464), .I2(\FRAME_MATCHER.state_c [3]), 
            .I3(GND_net), .O(n13496));
    defparam i11148_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_632 (.I0(\data_out_frame2[15] [6]), .I1(\data_out_frame2[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9853));   // coms.v(229[16:299])
    defparam i1_2_lut_adj_632.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame2_0___i137 (.Q(\data_out_frame2[17] [0]), .C(CLK_c), 
           .D(n10821));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_7[[7__2181  (.Q(\data_out[7] [7]), .C(CLK_c), .E(VCC_net), 
            .D(n10849));   // coms.v(280[12] 380[6])
    SB_LUT4 i3112_3_lut_4_lut (.I0(n62), .I1(n13464), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(n8603), .O(n5543));
    defparam i3112_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_DFF data_out_frame2_0___i136 (.Q(\data_out_frame2[16] [7]), .C(CLK_c), 
           .D(n10820));   // coms.v(426[12] 547[6])
    SB_LUT4 i3_4_lut_adj_633 (.I0(\data_out_frame2[13] [0]), .I1(\data_out_frame2[16] [6]), 
            .I2(n9853), .I3(n9589), .O(n17046));   // coms.v(228[16:596])
    defparam i3_4_lut_adj_633.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_634 (.I0(\data_out_frame2[11] [5]), .I1(\data_out_frame2[11] [6]), 
            .I2(\data_out_frame2[11] [7]), .I3(GND_net), .O(n17019));   // coms.v(238[17:230])
    defparam i2_3_lut_adj_634.LUT_INIT = 16'h9696;
    SB_LUT4 n18023_bdd_4_lut (.I0(n18023), .I1(n17591), .I2(n17590), .I3(\byte_transmit_counter[2] ), 
            .O(n18026));
    defparam n18023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_997_28 (.CI(n15647), .I0(\FRAME_MATCHER.i [26]), .I1(n17889), 
            .CO(n15648));
    SB_LUT4 i1_2_lut_adj_635 (.I0(\FRAME_MATCHER.state_c [23]), .I1(\FRAME_MATCHER.state_c [30]), 
            .I2(GND_net), .I3(GND_net), .O(n16898));   // coms.v(457[5:29])
    defparam i1_2_lut_adj_635.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_636 (.I0(n62), .I1(n13464), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n2_adj_2330), .O(n5545));
    defparam i2_3_lut_4_lut_adj_636.LUT_INIT = 16'h0100;
    SB_LUT4 i8030_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n10390));
    defparam i8030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame2_0___i135 (.Q(\data_out_frame2[16] [6]), .C(CLK_c), 
           .D(n10819));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i134 (.Q(\data_out_frame2[16] [5]), .C(CLK_c), 
           .D(n10818));   // coms.v(426[12] 547[6])
    SB_LUT4 i10595_2_lut (.I0(\rand_setpoint[28] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2362[0]));   // coms.v(283[4] 379[11])
    defparam i10595_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_997_27_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [25]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(n17889), .I3(n15646), .O(\FRAME_MATCHER.i_31__N_1280 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_27_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_637 (.I0(\data_out_frame2[7] [6]), .I1(\data_out_frame2[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16936));   // coms.v(237[17:221])
    defparam i1_2_lut_adj_637.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_638 (.I0(n17019), .I1(\data_out_frame2[11] [4]), 
            .I2(\data_out_frame2[11] [3]), .I3(GND_net), .O(n9695));   // coms.v(238[17:230])
    defparam i2_3_lut_adj_638.LUT_INIT = 16'h9696;
    SB_LUT4 i10657_3_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n127), 
            .I2(n2275), .I3(n7198), .O(\FRAME_MATCHER.state_31__N_1440[1] ));   // coms.v(453[6] 455[9])
    defparam i10657_3_lut_4_lut.LUT_INIT = 16'hfbf0;
    SB_CARRY add_997_27 (.CI(n15646), .I0(\FRAME_MATCHER.i [25]), .I1(n17889), 
            .CO(n15647));
    SB_LUT4 add_997_26_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [24]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(n17889), .I3(n15645), .O(\FRAME_MATCHER.i_31__N_1280 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_26_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_26 (.CI(n15645), .I0(\FRAME_MATCHER.i [24]), .I1(n17889), 
            .CO(n15646));
    SB_LUT4 add_997_25_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [23]), .I1(\FRAME_MATCHER.i [23]), 
            .I2(n17889), .I3(n15644), .O(\FRAME_MATCHER.i_31__N_1280 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_25_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_25 (.CI(n15644), .I0(\FRAME_MATCHER.i [23]), .I1(n17889), 
            .CO(n15645));
    SB_LUT4 add_997_24_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [22]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(n17889), .I3(n15643), .O(\FRAME_MATCHER.i_31__N_1280 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_24_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_24 (.CI(n15643), .I0(\FRAME_MATCHER.i [22]), .I1(n17889), 
            .CO(n15644));
    SB_LUT4 i1_2_lut_adj_639 (.I0(\data_out_frame2[6] [4]), .I1(\data_out_frame2[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17037));   // coms.v(239[17:230])
    defparam i1_2_lut_adj_639.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_640 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n16871), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(n16772), .O(n13464));
    defparam i3_4_lut_adj_640.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame2_0___i133 (.Q(\data_out_frame2[16] [4]), .C(CLK_c), 
           .D(n10817));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_7[[6__2182  (.Q(\data_out[7] [6]), .C(CLK_c), .E(VCC_net), 
            .D(n10846));   // coms.v(280[12] 380[6])
    SB_LUT4 i8031_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16882), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n10391));
    defparam i8031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10761_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [9]), .O(\FRAME_MATCHER.i_31__N_1312 [9]));
    defparam i10761_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 n18005_bdd_4_lut (.I0(n18005), .I1(\data_out_frame2[13] [6]), 
            .I2(\data_out_frame2[12] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n18008));
    defparam n18005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .D(n10467));   // coms.v(280[12] 380[6])
    SB_LUT4 i1_2_lut_adj_641 (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16963));   // coms.v(227[16:31])
    defparam i1_2_lut_adj_641.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_642 (.I0(\data_out_frame2[14] [6]), .I1(\data_out_frame2[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17106));   // coms.v(230[16:237])
    defparam i1_2_lut_adj_642.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_643 (.I0(\data_out[8] [1]), .I1(\data_out[8]_c [2]), 
            .I2(\data_out[8]_c [3]), .I3(GND_net), .O(n32_adj_2297));   // coms.v(21[11:19])
    defparam i1_2_lut_3_lut_adj_643.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame2_0___i2 (.Q(\data_out_frame2[0] [1]), .C(CLK_c), 
           .D(n17351));   // coms.v(426[12] 547[6])
    SB_DFFE \data_out_7[[5__2183  (.Q(\data_out[7] [5]), .C(CLK_c), .E(VCC_net), 
            .D(n10843));   // coms.v(280[12] 380[6])
    SB_LUT4 i7_4_lut_adj_644 (.I0(\data_out_frame2[15] [7]), .I1(\data_out_frame2[16] [4]), 
            .I2(n9695), .I3(n16936), .O(n18_adj_2331));   // coms.v(241[17:248])
    defparam i7_4_lut_adj_644.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(n17046), .I1(n17100), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_2332));   // coms.v(241[17:248])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_645 (.I0(n17106), .I1(n18_adj_2331), .I2(\data_out_frame2[10] [0]), 
            .I3(\data_out_frame2[11] [2]), .O(n20_adj_2333));   // coms.v(241[17:248])
    defparam i9_4_lut_adj_645.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_646 (.I0(n16963), .I1(n20_adj_2333), .I2(n16_adj_2332), 
            .I3(n17037), .O(n17108));   // coms.v(241[17:248])
    defparam i10_4_lut_adj_646.LUT_INIT = 16'h6996;
    SB_LUT4 i14890_3_lut (.I0(\data_out_frame2[0] [7]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17328));
    defparam i14890_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_2_lut_3_lut_adj_647 (.I0(\data_out[10] [3]), .I1(\data_out[6] [3]), 
            .I2(\data_out[6] [5]), .I3(GND_net), .O(n17028));   // coms.v(179[16:84])
    defparam i1_2_lut_3_lut_adj_647.LUT_INIT = 16'h9696;
    SB_LUT4 i14892_4_lut (.I0(n17328), .I1(n15846), .I2(n5543), .I3(n5545), 
            .O(n17330));
    defparam i14892_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14893_3_lut (.I0(\data_out_frame2[0] [6]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17331));
    defparam i14893_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8483_4_lut_4_lut (.I0(n10054), .I1(n2546[0]), .I2(\rand_setpoint[13] ), 
            .I3(\data_out[7] [5]), .O(n10843));
    defparam i8483_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 add_997_23_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [21]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(n17889), .I3(n15642), .O(\FRAME_MATCHER.i_31__N_1280 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_23_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame2[6] [0]), 
            .I1(\data_out_frame2[7] [0]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2334));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14895_4_lut (.I0(n17331), .I1(n15846), .I2(n5543), .I3(n5545), 
            .O(n17333));
    defparam i14895_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame2[5] [0]), 
            .I1(n5_adj_2334), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2335));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i8023_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n10383));
    defparam i8023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_648 (.I0(\data_out[8] [1]), .I1(n28_adj_2287), 
            .I2(\data_out[6] [4]), .I3(\data_out[8] [0]), .O(n16998));   // coms.v(176[16:77])
    defparam i2_3_lut_4_lut_adj_648.LUT_INIT = 16'h6996;
    SB_LUT4 i7942_2_lut (.I0(n10052), .I1(\FRAME_MATCHER.state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n10297));   // coms.v(493[6] 500[9])
    defparam i7942_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8486_4_lut_4_lut (.I0(n10054), .I1(n2546[0]), .I2(\rand_setpoint[14] ), 
            .I3(\data_out[7] [6]), .O(n10846));
    defparam i8486_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i8489_4_lut_4_lut (.I0(n10054), .I1(n2546[0]), .I2(\rand_setpoint[15] ), 
            .I3(\data_out[7] [7]), .O(n10849));
    defparam i8489_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i15294_2_lut (.I0(\data_out_frame2[0] [0]), .I1(byte_transmit_counter2[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17560));
    defparam i15294_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_997_23 (.CI(n15642), .I0(\FRAME_MATCHER.i [21]), .I1(n17889), 
            .CO(n15643));
    SB_CARRY add_2495_6 (.CI(n15517), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n15518));
    SB_LUT4 add_2495_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n15522), .O(n6517[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_649 (.I0(\FRAME_MATCHER.state_c [19]), .I1(\FRAME_MATCHER.state_c [26]), 
            .I2(\FRAME_MATCHER.state_c [25]), .I3(n16761), .O(n10_adj_2336));
    defparam i4_4_lut_adj_649.LUT_INIT = 16'hfffe;
    SB_LUT4 i14863_4_lut (.I0(n17560), .I1(n6_adj_2335), .I2(byte_transmit_counter2[2]), 
            .I3(byte_transmit_counter2[1]), .O(n17301));
    defparam i14863_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i14896_3_lut (.I0(\data_out_frame2[0] [5]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17334));
    defparam i14896_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14898_4_lut (.I0(n17334), .I1(n15846), .I2(n5543), .I3(n5545), 
            .O(n17336));
    defparam i14898_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut (.I0(n18104), .I1(\data_out_frame2[20] [0]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2337));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14865_3_lut (.I0(n17301), .I1(n18056), .I2(byte_transmit_counter2[3]), 
            .I3(GND_net), .O(n17303));
    defparam i14865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8479_4_lut_4_lut (.I0(n10054), .I1(n2546[0]), .I2(\rand_setpoint[12] ), 
            .I3(\data_out[7] [4]), .O(n10839));
    defparam i8479_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_DFF byte_transmit_counter__i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
           .D(n16269));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
           .D(n16283));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
           .D(n16261));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i4 (.Q(\byte_transmit_counter[4] ), .C(CLK_c), 
           .D(n16267));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i3 (.Q(\byte_transmit_counter[3] ), .C(CLK_c), 
           .D(n16285));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i2 (.Q(\byte_transmit_counter[2] ), .C(CLK_c), 
           .D(n16281));   // coms.v(280[12] 380[6])
    SB_DFF byte_transmit_counter__i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
           .D(n16257));   // coms.v(280[12] 380[6])
    SB_DFF data_out_frame2_0___i3 (.Q(\data_out_frame2[0] [2]), .C(CLK_c), 
           .D(n17345));   // coms.v(426[12] 547[6])
    SB_LUT4 i10762_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [8]), .O(\FRAME_MATCHER.i_31__N_1312 [8]));
    defparam i10762_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 equal_40_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_2310));   // coms.v(450[7:23])
    defparam equal_40_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_650 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n16133), 
            .I2(n10_adj_2336), .I3(n16898), .O(n62));
    defparam i1_4_lut_adj_650.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_651 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n16895), .I3(GND_net), .O(n16897));   // coms.v(450[7:23])
    defparam i1_2_lut_3_lut_adj_651.LUT_INIT = 16'hfefe;
    SB_LUT4 i10763_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [7]), .O(\FRAME_MATCHER.i_31__N_1312 [7]));
    defparam i10763_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10764_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [6]), .O(\FRAME_MATCHER.i_31__N_1312 [6]));
    defparam i10764_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8107_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[2]), .I3(delay_counter[2]), 
            .O(n10467));
    defparam i8107_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i1_2_lut_adj_652 (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_2330));
    defparam i1_2_lut_adj_652.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_653 (.I0(n13464), .I1(n62), .I2(n31), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n5_adj_2339));
    defparam i1_4_lut_adj_653.LUT_INIT = 16'h1101;
    SB_LUT4 i1_2_lut_adj_654 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16814));
    defparam i1_2_lut_adj_654.LUT_INIT = 16'h2222;
    SB_LUT4 i8104_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[1]), .I3(delay_counter[1]), 
            .O(n10464));
    defparam i8104_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i4_4_lut_adj_655 (.I0(\data_in_frame[2] [3]), .I1(n2336), .I2(n9541), 
            .I3(\data_in_frame[2] [5]), .O(n20_adj_2340));
    defparam i4_4_lut_adj_655.LUT_INIT = 16'h7bde;
    SB_LUT4 i8134_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[11]), .I3(delay_counter[11]), 
            .O(n10494));
    defparam i8134_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i7_4_lut_adj_656 (.I0(\data_in_frame[0] [7]), .I1(n2352), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[1] [7]), .O(n23_adj_2341));
    defparam i7_4_lut_adj_656.LUT_INIT = 16'hde7b;
    SB_LUT4 i11_4_lut_adj_657 (.I0(\data_in_frame[1] [2]), .I1(n22_adj_2301), 
            .I2(\data_in_frame[2] [2]), .I3(n9585), .O(n27_adj_2342));
    defparam i11_4_lut_adj_657.LUT_INIT = 16'hdffd;
    SB_LUT4 i8131_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[10]), .I3(delay_counter[10]), 
            .O(n10491));
    defparam i8131_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i2_4_lut_adj_658 (.I0(n2351), .I1(n2334), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[2] [4]), .O(n18_adj_2343));
    defparam i2_4_lut_adj_658.LUT_INIT = 16'hb7ed;
    SB_LUT4 i10_4_lut_adj_659 (.I0(n2342), .I1(n20_adj_2340), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[1] [0]), .O(n26_adj_2344));
    defparam i10_4_lut_adj_659.LUT_INIT = 16'hefdf;
    SB_LUT4 i14_4_lut_adj_660 (.I0(n27_adj_2342), .I1(n23_adj_2341), .I2(\data_in_frame[1] [3]), 
            .I3(\data_in_frame[1] [4]), .O(n30_adj_2345));
    defparam i14_4_lut_adj_660.LUT_INIT = 16'hefff;
    SB_LUT4 i1_4_lut_adj_661 (.I0(n2352), .I1(n2338), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[2] [6]), .O(n17_adj_2346));
    defparam i1_4_lut_adj_661.LUT_INIT = 16'h7bde;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut (.I0(n17303), .I1(n22_adj_2337), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[0]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15_4_lut_adj_662 (.I0(n17_adj_2346), .I1(n30_adj_2345), .I2(n26_adj_2344), 
            .I3(n18_adj_2343), .O(n31));
    defparam i15_4_lut_adj_662.LUT_INIT = 16'hfffe;
    SB_LUT4 i15387_3_lut (.I0(\data_out_frame2[0] [5]), .I1(byte_transmit_counter2[1]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17571));
    defparam i15387_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i14899_3_lut (.I0(\data_out_frame2[0] [4]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17337));
    defparam i14899_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14901_3_lut (.I0(n17337), .I1(n17769), .I2(n5543), .I3(GND_net), 
            .O(n17339));
    defparam i14901_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8128_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[9]), .I3(delay_counter[9]), 
            .O(n10488));
    defparam i8128_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i8125_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[8]), .I3(delay_counter[8]), 
            .O(n10485));
    defparam i8125_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i14903_3_lut (.I0(n31), .I1(n15846), .I2(n5545), .I3(GND_net), 
            .O(n17769));
    defparam i14903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8119_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[6]), .I3(delay_counter[6]), 
            .O(n10479));
    defparam i8119_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 add_2495_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n15516), .O(n6517[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8113_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[4]), .I3(delay_counter[4]), 
            .O(n10473));
    defparam i8113_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i12754_3_lut (.I0(delay_counter[13]), .I1(n17639), .I2(n1419), 
            .I3(GND_net), .O(n10859));
    defparam i12754_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_997_22_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [20]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(n17889), .I3(n15641), .O(\FRAME_MATCHER.i_31__N_1280 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_22_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_2495_5 (.CI(n15516), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n15517));
    SB_CARRY add_2495_11 (.CI(n15522), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n15523));
    SB_LUT4 add_2495_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n15521), .O(n6517[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14902_3_lut (.I0(\data_out_frame2[0] [3]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17340));
    defparam i14902_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10765_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [5]), .O(\FRAME_MATCHER.i_31__N_1312 [5]));
    defparam i10765_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_997_22 (.CI(n15641), .I0(\FRAME_MATCHER.i [20]), .I1(n17889), 
            .CO(n15642));
    SB_LUT4 i3_4_lut_adj_663 (.I0(n5_adj_2339), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n16814), .I3(\FRAME_MATCHER.state[0] ), .O(n10052));
    defparam i3_4_lut_adj_663.LUT_INIT = 16'h8020;
    SB_LUT4 i1_2_lut_4_lut_adj_664 (.I0(\data_out[6] [1]), .I1(\data_out[7] [7]), 
            .I2(\data_out[8] [1]), .I3(\data_out[8] [0]), .O(n16990));   // coms.v(175[16:77])
    defparam i1_2_lut_4_lut_adj_664.LUT_INIT = 16'h6996;
    SB_LUT4 i8110_4_lut_4_lut (.I0(n1419), .I1(n29), .I2(n6517[3]), .I3(delay_counter[3]), 
            .O(n10470));
    defparam i8110_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i1_2_lut_4_lut_adj_665 (.I0(\data_out_frame2[9] [2]), .I1(\data_out_frame2[5] [6]), 
            .I2(\data_out_frame2[9] [4]), .I3(\data_out_frame2[0] [0]), 
            .O(n6_adj_2293));   // coms.v(229[16:299])
    defparam i1_2_lut_4_lut_adj_665.LUT_INIT = 16'h6996;
    SB_LUT4 i14904_3_lut (.I0(n17340), .I1(n17769), .I2(n5543), .I3(GND_net), 
            .O(n17342));
    defparam i14904_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 n17897_bdd_4_lut (.I0(n17897), .I1(n9_adj_2347), .I2(n8_adj_2348), 
            .I3(byte_transmit_counter2[2]), .O(n17900));
    defparam n17897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame2[6] [5]), 
            .I1(\data_out_frame2[7] [5]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2349));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17993_bdd_4_lut (.I0(n17993), .I1(\data_out_frame2[9] [5]), 
            .I2(\data_out_frame2[8] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n17393));
    defparam n17993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out[6] [3]), 
            .I1(\data_out[7] [3]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2350));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_666 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n13272), .O(n16882));   // coms.v(450[7:23])
    defparam i1_3_lut_4_lut_adj_666.LUT_INIT = 16'hefff;
    SB_LUT4 equal_42_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_2329));   // coms.v(450[7:23])
    defparam equal_42_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15261_2_lut (.I0(\data_out[5] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17546));
    defparam i15261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut (.I0(\data_out_frame2[8] [4]), 
            .I1(\data_out_frame2[9] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n8_adj_2348));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_15557 (.I0(byte_transmit_counter[1]), 
            .I1(n17546), .I2(n5_adj_2350), .I3(\byte_transmit_counter[2] ), 
            .O(n18017));
    defparam byte_transmit_counter_1__bdd_4_lut_15557.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_667 (.I0(\data_out[9] [4]), .I1(\data_out[10] [0]), 
            .I2(\data_out[6] [2]), .I3(\data_out[6][0] ), .O(n16975));   // coms.v(174[16:77])
    defparam i2_3_lut_4_lut_adj_667.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut (.I0(\data_out_frame2[10] [4]), 
            .I1(\data_out_frame2[11] [4]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n9_adj_2347));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_997_21_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [19]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(n17889), .I3(n15640), .O(\FRAME_MATCHER.i_31__N_1280 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_21_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i14905_3_lut (.I0(\data_out_frame2[0] [2]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17343));
    defparam i14905_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14907_3_lut (.I0(n17343), .I1(n17769), .I2(n5543), .I3(GND_net), 
            .O(n17345));
    defparam i14907_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12_4_lut_adj_668 (.I0(byte_transmit_counter[1]), .I1(tx_transmit_N_1949[1]), 
            .I2(n10181), .I3(n16839), .O(n16257));   // coms.v(19[11:32])
    defparam i12_4_lut_adj_668.LUT_INIT = 16'h0aca;
    SB_CARRY add_2495_10 (.CI(n15521), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n15522));
    SB_LUT4 add_2495_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n15515), .O(n6517[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_669 (.I0(\byte_transmit_counter[2] ), .I1(tx_transmit_N_1949[2]), 
            .I2(n10181), .I3(n16839), .O(n16281));
    defparam i12_4_lut_adj_669.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut (.I0(\data_out_frame2[5] [5]), 
            .I1(n5_adj_2349), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2280));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i12_4_lut_adj_670 (.I0(\byte_transmit_counter[3] ), .I1(tx_transmit_N_1949[3]), 
            .I2(n10181), .I3(n16839), .O(n16285));
    defparam i12_4_lut_adj_670.LUT_INIT = 16'h0aca;
    SB_DFF data_out_frame2_0___i4 (.Q(\data_out_frame2[0] [3]), .C(CLK_c), 
           .D(n17342));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i5 (.Q(\data_out_frame2[0] [4]), .C(CLK_c), 
           .D(n17339));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i6 (.Q(\data_out_frame2[0] [5]), .C(CLK_c), 
           .D(n17336));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i7 (.Q(\data_out_frame2[0] [6]), .C(CLK_c), 
           .D(n17333));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i8 (.Q(\data_out_frame2[0] [7]), .C(CLK_c), 
           .D(n17330));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i153 (.Q(\data_out_frame2[19] [0]), .C(CLK_c), 
            .E(n10197), .D(n17108));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i154 (.Q(\data_out_frame2[19] [1]), .C(CLK_c), 
            .E(n10197), .D(n17011));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i155 (.Q(\data_out_frame2[19] [2]), .C(CLK_c), 
            .E(n10197), .D(n17131));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i156 (.Q(\data_out_frame2[19] [3]), .C(CLK_c), 
            .E(n10197), .D(n17132));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i157 (.Q(\data_out_frame2[19] [4]), .C(CLK_c), 
            .E(n10197), .D(n17114));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i158 (.Q(\data_out_frame2[19] [5]), .C(CLK_c), 
            .E(n10197), .D(n17113));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i159 (.Q(\data_out_frame2[19] [6]), .C(CLK_c), 
            .E(n10197), .D(n17107));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i160 (.Q(\data_out_frame2[19] [7]), .C(CLK_c), 
            .E(n10197), .D(n17135));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i161 (.Q(\data_out_frame2[20] [0]), .C(CLK_c), 
            .E(n10197), .D(n17104));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i162 (.Q(\data_out_frame2[20] [1]), .C(CLK_c), 
            .E(n10197), .D(n17105));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i163 (.Q(\data_out_frame2[20] [2]), .C(CLK_c), 
            .E(n10197), .D(n17053));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i164 (.Q(\data_out_frame2[20] [3]), .C(CLK_c), 
            .E(n10197), .D(n17122));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i165 (.Q(\data_out_frame2[20] [4]), .C(CLK_c), 
            .E(n10197), .D(n17123));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i166 (.Q(\data_out_frame2[20] [5]), .C(CLK_c), 
            .E(n10197), .D(n17126));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i167 (.Q(\data_out_frame2[20] [6]), .C(CLK_c), 
            .E(n10197), .D(n17125));   // coms.v(426[12] 547[6])
    SB_DFFE data_out_frame2_0___i168 (.Q(\data_out_frame2[20] [7]), .C(CLK_c), 
            .E(n10197), .D(n17128));   // coms.v(426[12] 547[6])
    SB_DFF data_out_frame2_0___i111 (.Q(\data_out_frame2[13] [6]), .C(CLK_c), 
           .D(n10795));   // coms.v(426[12] 547[6])
    SB_LUT4 i12_4_lut_adj_671 (.I0(\byte_transmit_counter[4] ), .I1(tx_transmit_N_1949[4]), 
            .I2(n10181), .I3(n16839), .O(n16267));
    defparam i12_4_lut_adj_671.LUT_INIT = 16'h0aca;
    SB_LUT4 i14852_3_lut_4_lut (.I0(tx_transmit_N_1949[6]), .I1(tx_transmit_N_1949[4]), 
            .I2(n5_adj_2319), .I3(n17254), .O(n17290));
    defparam i14852_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_3_lut (.I0(tx_transmit_N_1949[6]), .I1(tx_transmit_N_1949[4]), 
            .I2(n5_adj_2319), .I3(GND_net), .O(n8938));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_672 (.I0(byte_transmit_counter[5]), .I1(tx_transmit_N_1949[5]), 
            .I2(n10181), .I3(n16839), .O(n16261));
    defparam i12_4_lut_adj_672.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_3_lut_4_lut_adj_673 (.I0(\data_out_frame2[7] [4]), .I1(\data_out_frame2[5] [5]), 
            .I2(n10_adj_2292), .I3(n9910), .O(n16972));   // coms.v(227[16:31])
    defparam i5_3_lut_4_lut_adj_673.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_4_lut (.I0(\data_out_frame2[8] [1]), .I1(\data_out_frame2[15] [1]), 
            .I2(n9895), .I3(\data_out_frame2[14] [3]), .O(n23_adj_2318));   // coms.v(237[17:221])
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_674 (.I0(\data_out_frame2[8] [1]), .I1(\data_out_frame2[15] [1]), 
            .I2(\data_out_frame2[9] [6]), .I3(\data_out_frame2[8] [4]), 
            .O(n14_adj_2323));   // coms.v(237[17:221])
    defparam i5_3_lut_4_lut_adj_674.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_675 (.I0(byte_transmit_counter[6]), .I1(tx_transmit_N_1949[6]), 
            .I2(n10181), .I3(n16839), .O(n16283));
    defparam i12_4_lut_adj_675.LUT_INIT = 16'h0aca;
    SB_LUT4 i14816_3_lut_4_lut (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(tx_transmit_N_1949[3]), 
            .O(n17254));
    defparam i14816_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i12_4_lut_adj_676 (.I0(byte_transmit_counter[7]), .I1(tx_transmit_N_1949[7]), 
            .I2(n10181), .I3(n16839), .O(n16269));
    defparam i12_4_lut_adj_676.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_4_lut_adj_677 (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(tx_transmit_N_1949[3]), .I3(n8938), .O(n22_adj_2164));
    defparam i1_3_lut_4_lut_adj_677.LUT_INIT = 16'hffe0;
    SB_LUT4 i2_3_lut_4_lut_adj_678 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n16891), .O(n16893));
    defparam i2_3_lut_4_lut_adj_678.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_4_lut_adj_679 (.I0(n9505), .I1(\data_out[9] [6]), .I2(\data_out[9][2] ), 
            .I3(n17064), .O(data_out_10__2__N_157));   // coms.v(172[16:77])
    defparam i1_2_lut_4_lut_adj_679.LUT_INIT = 16'h6996;
    SB_LUT4 i10766_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [4]), .O(\FRAME_MATCHER.i_31__N_1312 [4]));
    defparam i10766_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15224_3_lut (.I0(\data_out_frame2[0] [7]), .I1(byte_transmit_counter2[0]), 
            .I2(byte_transmit_counter2[1]), .I3(GND_net), .O(n17561));
    defparam i15224_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_4_lut_adj_680 (.I0(n17475), .I1(n17230), .I2(n17290), .I3(\UART_TRANSMITTER.state[2] ), 
            .O(n16838));   // coms.v(283[4] 379[11])
    defparam i1_4_lut_adj_680.LUT_INIT = 16'h0322;
    SB_CARRY add_997_21 (.CI(n15640), .I0(\FRAME_MATCHER.i [19]), .I1(n17889), 
            .CO(n15641));
    SB_LUT4 i14911_3_lut (.I0(\data_out_frame2[0] [1]), .I1(n16148), .I2(n5545), 
            .I3(GND_net), .O(n17349));
    defparam i14911_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame2[6] [7]), 
            .I1(\data_out_frame2[7] [7]), .I2(byte_transmit_counter2[0]), 
            .I3(GND_net), .O(n5_adj_2351));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut (.I0(\data_out_frame2[5] [7]), 
            .I1(n5_adj_2351), .I2(byte_transmit_counter2[1]), .I3(byte_transmit_counter2[0]), 
            .O(n6_adj_2278));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i14913_4_lut (.I0(n17349), .I1(n15846), .I2(n5543), .I3(n5545), 
            .O(n17351));
    defparam i14913_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_3_lut_adj_681 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n16895), .I3(GND_net), .O(n16896));
    defparam i1_2_lut_3_lut_adj_681.LUT_INIT = 16'hf7f7;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15577 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [6]), .I2(\data_out_frame2[15] [6]), 
            .I3(byte_transmit_counter2[1]), .O(n18005));
    defparam byte_transmit_counter2_0__bdd_4_lut_15577.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_682 (.I0(\data_out_frame2[8] [0]), .I1(\data_out_frame2[16] [1]), 
            .I2(n9892), .I3(\data_out_frame2[11] [6]), .O(n17079));   // coms.v(237[17:221])
    defparam i2_3_lut_4_lut_adj_682.LUT_INIT = 16'h6996;
    SB_LUT4 i10565_2_lut (.I0(\rand_setpoint[27] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2397[0]));   // coms.v(283[4] 379[11])
    defparam i10565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_997_20_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [18]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(n17889), .I3(n15639), .O(\FRAME_MATCHER.i_31__N_1280 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_20_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_20 (.CI(n15639), .I0(\FRAME_MATCHER.i [18]), .I1(n17889), 
            .CO(n15640));
    SB_LUT4 i10561_2_lut (.I0(\rand_setpoint[26] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2432[0]));   // coms.v(283[4] 379[11])
    defparam i10561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15331_2_lut (.I0(\data_out[0][0] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17581));
    defparam i15331_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_683 (.I0(\data_out[7] [3]), .I1(\data_out[9][2] ), 
            .I2(\data_out[5] [4]), .I3(GND_net), .O(n17055));   // coms.v(182[17:86])
    defparam i1_2_lut_3_lut_adj_683.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_684 (.I0(\data_out_frame2[8] [0]), .I1(\data_out_frame2[16] [1]), 
            .I2(\data_out_frame2[13] [3]), .I3(GND_net), .O(n6_adj_2286));   // coms.v(237[17:221])
    defparam i1_2_lut_3_lut_adj_684.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i2_3_lut (.I0(\data_out[2][0] ), 
            .I1(\data_out[3][0] ), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n2_adj_2266));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8251_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n10611));
    defparam i8251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out[6][0] ), 
            .I1(\data_out[7] [0]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2265));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut (.I0(n18062), .I1(\data_out_frame2[20] [7]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2352));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut (.I0(n18092), .I1(n22_adj_2352), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[7]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i4944_2_lut (.I0(n127), .I1(n127_adj_2136), .I2(GND_net), 
            .I3(GND_net), .O(n7212));   // coms.v(440[13] 443[7])
    defparam i4944_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut (.I0(n18002), .I1(\data_out_frame2[20] [6]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2353));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10767_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [3]), .O(\FRAME_MATCHER.i_31__N_1312 [3]));
    defparam i10767_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_4_lut_adj_685 (.I0(\data_out_frame2[0] [3]), .I1(\data_out_frame2[0] [2]), 
            .I2(\data_out_frame2[0] [4]), .I3(\data_out_frame2[0] [1]), 
            .O(n9919));
    defparam i2_3_lut_4_lut_adj_685.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_686 (.I0(\data_out[10] [1]), .I1(\data_out[10] [5]), 
            .I2(data_out_9__2__N_367), .I3(GND_net), .O(n17094));   // coms.v(178[16:77])
    defparam i1_2_lut_3_lut_adj_686.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut (.I0(n18086), .I1(n22_adj_2353), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[6]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15367_2_lut (.I0(data_out_6__1__N_537), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17632));
    defparam i15367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10768_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [2]), .O(\FRAME_MATCHER.i_31__N_1312 [2]));
    defparam i10768_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8252_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n10612));
    defparam i8252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10769_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(\FRAME_MATCHER.i [1]), .O(\FRAME_MATCHER.i_31__N_1312 [1]));
    defparam i10769_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_238_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [0]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_c));
    defparam select_238_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_687 (.I0(\data_out_frame2[15] [6]), .I1(\data_out_frame2[7] [6]), 
            .I2(\data_out_frame2[5] [7]), .I3(GND_net), .O(n17127));   // coms.v(234[16:291])
    defparam i1_2_lut_3_lut_adj_687.LUT_INIT = 16'h9696;
    SB_LUT4 i15255_3_lut_4_lut (.I0(data_out_7__3__N_441), .I1(\UART_TRANSMITTER.state[2] ), 
            .I2(\data_out[5] [5]), .I3(n17025), .O(n17534));   // coms.v(283[4] 379[11])
    defparam i15255_3_lut_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i8253_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n10613));
    defparam i8253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8254_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n10614));
    defparam i8254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15401_4_lut (.I0(n446), .I1(n456), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n10031));
    defparam i15401_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i8255_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n10615));
    defparam i8255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15213_3_lut_4_lut (.I0(data_out_7__2__N_447), .I1(data_out_7__3__N_441), 
            .I2(\UART_TRANSMITTER.state[2] ), .I3(n17025), .O(n17532));   // coms.v(283[4] 379[11])
    defparam i15213_3_lut_4_lut.LUT_INIT = 16'h6090;
    SB_LUT4 i8256_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n10616));
    defparam i8256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut (.I0(n17984), .I1(\data_out_frame2[20] [5]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2354));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut (.I0(n17966), .I1(n22_adj_2354), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[5]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8257_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n10617));
    defparam i8257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8258_3_lut_4_lut (.I0(n8_adj_2310), .I1(n16891), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n10618));
    defparam i8258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_997_19_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [17]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(n17889), .I3(n15638), .O(\FRAME_MATCHER.i_31__N_1280 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10624_2_lut (.I0(\rand_setpoint[24] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2502[0]));   // coms.v(283[4] 379[11])
    defparam i10624_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_997_19 (.CI(n15638), .I0(\FRAME_MATCHER.i [17]), .I1(n17889), 
            .CO(n15639));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut (.I0(n17972), .I1(\data_out_frame2[20] [4]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2355));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_997_18_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [16]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(n17889), .I3(n15637), .O(\FRAME_MATCHER.i_31__N_1280 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_18_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15414_3_lut (.I0(n5545), .I1(n5543), .I2(n31), .I3(GND_net), 
            .O(n10197));
    defparam i15414_3_lut.LUT_INIT = 16'h0404;
    SB_CARRY add_997_18 (.CI(n15637), .I0(\FRAME_MATCHER.i [16]), .I1(n17889), 
            .CO(n15638));
    SB_LUT4 i15357_2_lut_3_lut_4_lut (.I0(n127_adj_4), .I1(n127), .I2(n127_adj_2136), 
            .I3(n2275), .O(n17454));
    defparam i15357_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_adj_688 (.I0(\data_out[8][5] ), .I1(\data_out[8][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n16949));   // coms.v(181[17:93])
    defparam i1_2_lut_adj_688.LUT_INIT = 16'h6666;
    SB_LUT4 i11219217_i1_3_lut (.I0(n17990), .I1(n17900), .I2(byte_transmit_counter2[3]), 
            .I3(GND_net), .O(n15_adj_2356));
    defparam i11219217_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut (.I0(n15_adj_2356), 
            .I1(n22_adj_2355), .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[4]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_997_17_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [15]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(n17889), .I3(n15636), .O(\FRAME_MATCHER.i_31__N_1280 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_17_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_689 (.I0(\data_out[8][4] ), .I1(\data_out[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9728));   // coms.v(178[16:77])
    defparam i1_2_lut_adj_689.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_690 (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(n9357), .I3(\UART_TRANSMITTER.state[2] ), .O(n44_adj_2163));
    defparam i1_3_lut_4_lut_adj_690.LUT_INIT = 16'hf0f8;
    SB_CARRY add_997_17 (.CI(n15636), .I0(\FRAME_MATCHER.i [15]), .I1(n17889), 
            .CO(n15637));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut (.I0(n17948), .I1(\data_out_frame2[20] [3]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2357));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut (.I0(n18128), .I1(n22_adj_2357), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[3]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_691 (.I0(n127_adj_2136), .I1(n127_adj_4), 
            .I2(n9346), .I3(\FRAME_MATCHER.i [31]), .O(n9435));   // coms.v(529[6] 531[9])
    defparam i1_2_lut_4_lut_adj_691.LUT_INIT = 16'h8808;
    SB_LUT4 i1_2_lut_3_lut_adj_692 (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(n9357), .I3(GND_net), .O(n9358));
    defparam i1_2_lut_3_lut_adj_692.LUT_INIT = 16'hf8f8;
    SB_LUT4 n17981_bdd_4_lut (.I0(n17981), .I1(\data_out_frame2[17] [5]), 
            .I2(\data_out_frame2[16] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n17984));
    defparam n17981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_2495_9_lut (.I0(n29), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n15520), .O(n17638)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2495_9 (.CI(n15520), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n15521));
    SB_LUT4 add_997_16_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [14]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(n17889), .I3(n15635), .O(\FRAME_MATCHER.i_31__N_1280 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_16_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15533 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [5]), .I2(\data_out_frame2[19] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n17981));
    defparam byte_transmit_counter2_0__bdd_4_lut_15533.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1820_i1_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(tx2_transmit_N_1997), .O(n4130[0]));   // coms.v(444[4] 546[11])
    defparam mux_1820_i1_4_lut.LUT_INIT = 16'hd454;
    SB_LUT4 i4_4_lut_adj_693 (.I0(\data_out[10] [2]), .I1(n9728), .I2(\data_out[7] [0]), 
            .I3(n9716), .O(n10_adj_2162));   // coms.v(171[16:93])
    defparam i4_4_lut_adj_693.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_694 (.I0(\data_out_frame2[7] [7]), .I1(\data_out_frame2[7] [6]), 
            .I2(\data_out_frame2[9] [4]), .I3(GND_net), .O(n17091));   // coms.v(237[17:221])
    defparam i1_2_lut_3_lut_adj_694.LUT_INIT = 16'h9696;
    SB_LUT4 i15277_3_lut_4_lut (.I0(tx_transmit_N_1949[2]), .I1(n4_adj_2311), 
            .I2(\UART_TRANSMITTER.state[1] ), .I3(n9357), .O(n17475));
    defparam i15277_3_lut_4_lut.LUT_INIT = 16'h0070;
    SB_CARRY add_997_16 (.CI(n15635), .I0(\FRAME_MATCHER.i [14]), .I1(n17889), 
            .CO(n15636));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut (.I0(n17930), .I1(\data_out_frame2[20] [2]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2358));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11115_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n9451), 
            .I2(n12933), .I3(n9488), .O(n1439));
    defparam i11115_2_lut_3_lut_4_lut.LUT_INIT = 16'he000;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut (.I0(n18122), .I1(n22_adj_2358), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[2]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_1__bdd_4_lut_15582 (.I0(byte_transmit_counter2[1]), 
            .I1(n17495), .I2(n5_adj_2141), .I3(byte_transmit_counter2[2]), 
            .O(n17987));
    defparam byte_transmit_counter2_1__bdd_4_lut_15582.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_695 (.I0(\FRAME_MATCHER.state_c [14]), .I1(\FRAME_MATCHER.state_c [22]), 
            .I2(\FRAME_MATCHER.state_c [21]), .I3(\FRAME_MATCHER.state_c [19]), 
            .O(n52));   // coms.v(457[5:29])
    defparam i2_3_lut_4_lut_adj_695.LUT_INIT = 16'hfffe;
    SB_LUT4 add_997_15_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [13]), .I1(\FRAME_MATCHER.i [13]), 
            .I2(n17889), .I3(n15634), .O(\FRAME_MATCHER.i_31__N_1280 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[12] [5]), 
            .I2(\data_out_frame2[0] [3]), .I3(n17124), .O(n20_adj_2202));   // coms.v(232[16:229])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_696 (.I0(\data_out_frame2[16] [3]), .I1(\data_out_frame2[12] [5]), 
            .I2(\data_out_frame2[8] [7]), .I3(GND_net), .O(n17112));   // coms.v(232[16:229])
    defparam i1_2_lut_3_lut_adj_696.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut (.I0(n17912), .I1(\data_out_frame2[20] [1]), 
            .I2(byte_transmit_counter2[2]), .I3(n8621), .O(n22_adj_2359));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_997_15 (.CI(n15634), .I0(\FRAME_MATCHER.i [13]), .I1(n17889), 
            .CO(n15635));
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut (.I0(n18110), .I1(n22_adj_2359), 
            .I2(byte_transmit_counter2[4]), .I3(byte_transmit_counter2[3]), 
            .O(tx2_data[1]));   // coms.v(413[36:58])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8240_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n10600));
    defparam i8240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_238_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [1]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_adj_2260));
    defparam select_238_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8241_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n10601));
    defparam i8241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_2495_4 (.CI(n15515), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n15516));
    SB_LUT4 i6_2_lut_4_lut (.I0(\data_out_frame2[7] [7]), .I1(n16936), .I2(\data_out_frame2[7] [2]), 
            .I3(\data_out_frame2[14] [2]), .O(n18_adj_2251));   // coms.v(237[17:221])
    defparam i6_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_997_14_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [12]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(n17889), .I3(n15633), .O(\FRAME_MATCHER.i_31__N_1280 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_14_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i8242_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n10602));
    defparam i8242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n18017_bdd_4_lut (.I0(n18017), .I1(n17593), .I2(n17592), .I3(\byte_transmit_counter[2] ), 
            .O(n18020));
    defparam n18017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_997_14 (.CI(n15633), .I0(\FRAME_MATCHER.i [12]), .I1(n17889), 
            .CO(n15634));
    SB_LUT4 i2_4_lut_adj_697 (.I0(n4445), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n9361), .I3(n10031), .O(n15868));
    defparam i2_4_lut_adj_697.LUT_INIT = 16'hfefa;
    SB_LUT4 i6219_4_lut (.I0(n446), .I1(n456), .I2(\UART_TRANSMITTER.state[2] ), 
            .I3(\UART_TRANSMITTER.state[0] ), .O(n8631));   // coms.v(283[4] 379[11])
    defparam i6219_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i1_2_lut_4_lut_adj_698 (.I0(\data_in[2] [7]), .I1(\data_in[1] [2]), 
            .I2(\data_in[1] [1]), .I3(\data_in[3] [6]), .O(n12_adj_2200));
    defparam i1_2_lut_4_lut_adj_698.LUT_INIT = 16'hffef;
    SB_DFFESR byte_transmit_counter2_2353__i0 (.Q(byte_transmit_counter2[0]), 
            .C(CLK_c), .E(n10052), .D(n37[0]), .R(n10297));   // coms.v(493[6] 500[9])
    SB_LUT4 select_238_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [2]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_adj_2259));
    defparam select_238_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_2_lut_3_lut_adj_699 (.I0(\data_out_frame2[15] [3]), .I1(\data_out_frame2[7] [3]), 
            .I2(\data_out_frame2[9] [1]), .I3(GND_net), .O(n16_adj_2197));   // coms.v(232[16:229])
    defparam i3_2_lut_3_lut_adj_699.LUT_INIT = 16'h9696;
    SB_LUT4 i15288_2_lut (.I0(\data_out[1] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17590));
    defparam i15288_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 add_2495_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n15519), .O(n6517[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15289_2_lut (.I0(\data_out[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17591));
    defparam i15289_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_700 (.I0(n127_adj_4), .I1(n9346), .I2(\FRAME_MATCHER.i [31]), 
            .I3(GND_net), .O(n9393));   // coms.v(529[6] 531[9])
    defparam i1_2_lut_3_lut_adj_700.LUT_INIT = 16'ha2a2;
    SB_LUT4 i8243_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n10603));
    defparam i8243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_2495_8 (.CI(n15519), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n15520));
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15465 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[14] [5]), .I2(\data_out_frame2[15] [5]), 
            .I3(byte_transmit_counter2[1]), .O(n17891));
    defparam byte_transmit_counter2_0__bdd_4_lut_15465.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out[6] [4]), 
            .I1(\data_out[7] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n5_adj_2326));   // coms.v(257[28:49])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10929_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n9451), 
            .I2(n12933), .I3(rx_data_ready), .O(n13272));
    defparam i10929_2_lut_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_4_lut_adj_701 (.I0(n8631), .I1(n15868), .I2(n29), .I3(\UART_TRANSMITTER.state[1] ), 
            .O(n10141));
    defparam i1_4_lut_adj_701.LUT_INIT = 16'h2333;
    SB_LUT4 i14908_3_lut (.I0(\data_out_frame2[8] [0]), .I1(\data_out_frame2[9] [0]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17346));
    defparam i14908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14909_3_lut (.I0(\data_out_frame2[10] [0]), .I1(\data_out_frame2[11] [0]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17347));
    defparam i14909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15348_2_lut (.I0(\data_out[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17547));
    defparam i15348_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_238_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [3]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_adj_2258));
    defparam select_238_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10603_2_lut (.I0(\rand_setpoint[31] ), .I1(\UART_TRANSMITTER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n2257[0]));   // coms.v(283[4] 379[11])
    defparam i10603_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_702 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[10] [2]), .O(n15930));
    defparam i2_3_lut_4_lut_adj_702.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_703 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16331));
    defparam i1_2_lut_adj_703.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_704 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16439));
    defparam i1_2_lut_adj_704.LUT_INIT = 16'h8888;
    SB_LUT4 i14885_3_lut (.I0(\data_out_frame2[14] [0]), .I1(\data_out_frame2[15] [0]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17323));
    defparam i14885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_705 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16339));
    defparam i1_2_lut_adj_705.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_706 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16437));
    defparam i1_2_lut_adj_706.LUT_INIT = 16'h8888;
    SB_LUT4 i8244_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n10604));
    defparam i8244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_707 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16335));
    defparam i1_2_lut_adj_707.LUT_INIT = 16'h8888;
    SB_LUT4 i8248_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n10608));
    defparam i8248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_997_13_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [11]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(n17889), .I3(n15632), .O(\FRAME_MATCHER.i_31__N_1280 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i8249_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n10609));
    defparam i8249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_2495_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n15514), .O(n6517[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_997_13 (.CI(n15632), .I0(\FRAME_MATCHER.i [11]), .I1(n17889), 
            .CO(n15633));
    SB_LUT4 add_2495_7_lut (.I0(n29), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n15518), .O(n17574)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_708 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16435));
    defparam i1_2_lut_adj_708.LUT_INIT = 16'h8888;
    SB_LUT4 add_997_12_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [10]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(n17889), .I3(n15631), .O(\FRAME_MATCHER.i_31__N_1280 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_12_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_12 (.CI(n15631), .I0(\FRAME_MATCHER.i [10]), .I1(n17889), 
            .CO(n15632));
    SB_CARRY add_2495_3 (.CI(n15514), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n15515));
    SB_LUT4 add_997_11_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [9]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(n17889), .I3(n15630), .O(\FRAME_MATCHER.i_31__N_1280 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_11_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_11 (.CI(n15630), .I0(\FRAME_MATCHER.i [9]), .I1(n17889), 
            .CO(n15631));
    SB_LUT4 n17891_bdd_4_lut (.I0(n17891), .I1(\data_out_frame2[13] [5]), 
            .I2(\data_out_frame2[12] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n17894));
    defparam n17891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_2495_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n15514));
    SB_LUT4 i1_2_lut_adj_709 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16441));
    defparam i1_2_lut_adj_709.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_710 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16433));
    defparam i1_2_lut_adj_710.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_711 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16443));
    defparam i1_2_lut_adj_711.LUT_INIT = 16'h8888;
    SB_LUT4 i8250_3_lut_4_lut (.I0(n8), .I1(n16891), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n10610));
    defparam i8250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_997_10_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [8]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(n17889), .I3(n15629), .O(\FRAME_MATCHER.i_31__N_1280 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_712 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16431));
    defparam i1_2_lut_adj_712.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_713 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16445));
    defparam i1_2_lut_adj_713.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_714 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16429));
    defparam i1_2_lut_adj_714.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_715 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[10] [3]), .O(n15929));
    defparam i2_3_lut_4_lut_adj_715.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut_4_lut_adj_716 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[7] [7]), .O(n22));
    defparam i6_3_lut_4_lut_adj_716.LUT_INIT = 16'h9f6f;
    SB_LUT4 i1_2_lut_adj_717 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16455));
    defparam i1_2_lut_adj_717.LUT_INIT = 16'h8888;
    SB_LUT4 i8003_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10055), .I3(\data_out[2] [3]), .O(n10363));
    defparam i8003_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_15523 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_out_frame2[18] [4]), .I2(\data_out_frame2[19] [4]), 
            .I3(byte_transmit_counter2[1]), .O(n17969));
    defparam byte_transmit_counter2_0__bdd_4_lut_15523.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_718 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16427));
    defparam i1_2_lut_adj_718.LUT_INIT = 16'h8888;
    SB_CARRY add_997_10 (.CI(n15629), .I0(\FRAME_MATCHER.i [8]), .I1(n17889), 
            .CO(n15630));
    SB_LUT4 add_997_9_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [7]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(n17889), .I3(n15628), .O(\FRAME_MATCHER.i_31__N_1280 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_719 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16453));
    defparam i1_2_lut_adj_719.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_720 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16425));
    defparam i1_2_lut_adj_720.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_721 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16451));
    defparam i1_2_lut_adj_721.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_722 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16423));
    defparam i1_2_lut_adj_722.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_723 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16449));
    defparam i1_2_lut_adj_723.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_724 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16421));
    defparam i1_2_lut_adj_724.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_725 (.I0(n2), .I1(n7212), .I2(n12933), .I3(n9393), 
            .O(n4_adj_2360));
    defparam i1_4_lut_adj_725.LUT_INIT = 16'haeaa;
    SB_LUT4 i8008_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10055), .I3(\data_out[1] [4]), .O(n10368));
    defparam i8008_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_CARRY add_997_9 (.CI(n15628), .I0(\FRAME_MATCHER.i [7]), .I1(n17889), 
            .CO(n15629));
    SB_LUT4 i14884_3_lut (.I0(\data_out_frame2[12] [0]), .I1(\data_out_frame2[13] [0]), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n17322));
    defparam i14884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_726 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n4_adj_2360), 
            .I2(GND_net), .I3(GND_net), .O(n16447));
    defparam i1_2_lut_adj_726.LUT_INIT = 16'h8888;
    SB_LUT4 select_238_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [4]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_adj_2257));
    defparam select_238_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_727 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16419));
    defparam i1_2_lut_adj_727.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_728 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16351));
    defparam i1_2_lut_adj_728.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_729 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16417));
    defparam i1_2_lut_adj_729.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_730 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16349));
    defparam i1_2_lut_adj_730.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_731 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16415));
    defparam i1_2_lut_adj_731.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_732 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16347));
    defparam i1_2_lut_adj_732.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_733 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16413));
    defparam i1_2_lut_adj_733.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_734 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16345));
    defparam i1_2_lut_adj_734.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_735 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16411));
    defparam i1_2_lut_adj_735.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_736 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16343));
    defparam i1_2_lut_adj_736.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_737 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16409));
    defparam i1_2_lut_adj_737.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_738 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16371));
    defparam i1_2_lut_adj_738.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_739 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16407));
    defparam i1_2_lut_adj_739.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_740 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16369));
    defparam i1_2_lut_adj_740.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_741 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16405));
    defparam i1_2_lut_adj_741.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_742 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16367));
    defparam i1_2_lut_adj_742.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_743 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16403));
    defparam i1_2_lut_adj_743.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_744 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16365));
    defparam i1_2_lut_adj_744.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_745 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16401));
    defparam i1_2_lut_adj_745.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_746 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(n16943), .I3(GND_net), .O(n2351));   // coms.v(76[16:62])
    defparam i1_2_lut_3_lut_adj_746.LUT_INIT = 16'h9696;
    SB_LUT4 add_997_8_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [6]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(n17889), .I3(n15627), .O(\FRAME_MATCHER.i_31__N_1280 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_8 (.CI(n15627), .I0(\FRAME_MATCHER.i [6]), .I1(n17889), 
            .CO(n15628));
    SB_LUT4 i1_2_lut_adj_747 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16363));
    defparam i1_2_lut_adj_747.LUT_INIT = 16'h8888;
    SB_LUT4 i8010_3_lut_4_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(n10055), .I3(\data_out[0] [6]), .O(n10370));
    defparam i8010_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 select_238_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [5]), 
            .I1(n1439), .I2(GND_net), .I3(GND_net), .O(n3_adj_2256));
    defparam select_238_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_2_lut_3_lut (.I0(\UART_TRANSMITTER.state[2] ), .I1(\UART_TRANSMITTER.state[1] ), 
            .I2(\UART_TRANSMITTER.state[0] ), .I3(GND_net), .O(n10181));
    defparam i6_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_adj_748 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16399));
    defparam i1_2_lut_adj_748.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_749 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16361));
    defparam i1_2_lut_adj_749.LUT_INIT = 16'h8888;
    SB_LUT4 add_2495_16_lut (.I0(n29), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n15527), .O(n17635)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_750 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16397));
    defparam i1_2_lut_adj_750.LUT_INIT = 16'h8888;
    SB_LUT4 add_997_7_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [5]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n17889), .I3(n15626), .O(\FRAME_MATCHER.i_31__N_1280 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_7 (.CI(n15626), .I0(\FRAME_MATCHER.i [5]), .I1(n17889), 
            .CO(n15627));
    SB_LUT4 add_2495_15_lut (.I0(n29), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n15526), .O(n17639)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2495_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_997_6_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [4]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n17889), .I3(n15625), .O(\FRAME_MATCHER.i_31__N_1280 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_6 (.CI(n15625), .I0(\FRAME_MATCHER.i [4]), .I1(n17889), 
            .CO(n15626));
    SB_LUT4 i10592_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n9460), 
            .I2(n9451), .I3(GND_net), .O(n12933));
    defparam i10592_2_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_997_5_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [3]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n17889), .I3(n15624), .O(\FRAME_MATCHER.i_31__N_1280 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_997_5 (.CI(n15624), .I0(\FRAME_MATCHER.i [3]), .I1(n17889), 
            .CO(n15625));
    SB_LUT4 add_997_4_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [2]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n17889), .I3(n15623), .O(\FRAME_MATCHER.i_31__N_1280 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_adj_751 (.I0(n127), .I1(n127_adj_2136), .I2(n127_adj_4), 
            .I3(n16795), .O(n2));
    defparam i1_2_lut_4_lut_adj_751.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_adj_752 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16359));
    defparam i1_2_lut_adj_752.LUT_INIT = 16'h8888;
    SB_LUT4 i8016_3_lut_4_lut (.I0(n8), .I1(n16882), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n10376));
    defparam i8016_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame2_0___i110 (.Q(\data_out_frame2[13] [5]), .C(CLK_c), 
           .D(n10794));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_753 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16395));
    defparam i1_2_lut_adj_753.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n10392));   // coms.v(426[12] 547[6])
    SB_CARRY add_997_4 (.CI(n15623), .I0(\FRAME_MATCHER.i [2]), .I1(n17889), 
            .CO(n15624));
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n10391));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n10390));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_754 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16357));
    defparam i1_2_lut_adj_754.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_755 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16393));
    defparam i1_2_lut_adj_755.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_756 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16355));
    defparam i1_2_lut_adj_756.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n10389));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n10388));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n10387));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n10386));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n10385));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n10384));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_757 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16391));
    defparam i1_2_lut_adj_757.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n10383));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n10382));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n10381));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n10380));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n10379));   // coms.v(426[12] 547[6])
    SB_CARRY add_2495_15 (.CI(n15526), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n15527));
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n10378));   // coms.v(426[12] 547[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n10377));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_758 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16353));
    defparam i1_2_lut_adj_758.LUT_INIT = 16'h8888;
    SB_LUT4 add_997_3_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [1]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n17889), .I3(n15622), .O(\FRAME_MATCHER.i_31__N_1280 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n10376));   // coms.v(426[12] 547[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(CLK_c), 
           .D(n16327));   // coms.v(426[12] 547[6])
    SB_LUT4 i1_2_lut_adj_759 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16389));
    defparam i1_2_lut_adj_759.LUT_INIT = 16'h8888;
    SB_DFF \data_out_0[[0__2244  (.Q(\data_out[0][0] ), .C(CLK_c), .D(n10374));   // coms.v(280[12] 380[6])
    SB_CARRY add_997_3 (.CI(n15622), .I0(\FRAME_MATCHER.i [1]), .I1(n17889), 
            .CO(n15623));
    SB_LUT4 add_997_2_lut (.I0(\FRAME_MATCHER.i_31__N_1312 [0]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n17889), .I3(VCC_net), .O(\FRAME_MATCHER.i_31__N_1280 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_997_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_760 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16381));
    defparam i1_2_lut_adj_760.LUT_INIT = 16'h8888;
    SB_CARRY add_997_2 (.CI(VCC_net), .I0(\FRAME_MATCHER.i [0]), .I1(n17889), 
            .CO(n15622));
    SB_LUT4 byte_transmit_counter2_2353_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[7]), .I3(n15621), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_761 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16387));
    defparam i1_2_lut_adj_761.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_762 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n4_c), 
            .I2(GND_net), .I3(GND_net), .O(n16379));
    defparam i1_2_lut_adj_762.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_2353_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[6]), .I3(n15620), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_763 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n7), 
            .I2(GND_net), .I3(GND_net), .O(n16385));
    defparam i1_2_lut_adj_763.LUT_INIT = 16'h8888;
    SB_CARRY byte_transmit_counter2_2353_add_4_8 (.CI(n15620), .I0(GND_net), 
            .I1(byte_transmit_counter2[6]), .CO(n15621));
    SB_LUT4 byte_transmit_counter2_2353_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[5]), .I3(n15619), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_2353_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY byte_transmit_counter2_2353_add_4_7 (.CI(n15619), .I0(GND_net), 
            .I1(byte_transmit_counter2[5]), .CO(n15620));
    SB_LUT4 i1_2_lut_3_lut_adj_764 (.I0(n127), .I1(n127_adj_2136), .I2(n127_adj_4), 
            .I3(GND_net), .O(n8828));
    defparam i1_2_lut_3_lut_adj_764.LUT_INIT = 16'h8080;
    uart_tx tx (.r_SM_Main({r_SM_Main}), .n3(n3), .GND_net(GND_net), .\r_Bit_Index[1] (\r_Bit_Index[1] ), 
            .n14060(n14060), .\r_SM_Main_2__N_2036[0] (r_SM_Main_2__N_2036[0]), 
            .n5(n5), .n13276(n13276), .n16671(n16671), .r_Clock_Count({r_Clock_Count}), 
            .CLK_c(CLK_c), .n16651(n16651), .n16649(n16649), .n16567(n16567), 
            .n16509(n16509), .n16477(n16477), .n16467(n16467), .n16459(n16459), 
            .n16595(n16595), .r_Tx_Data({r_Tx_Data}), .n16625(n16625), 
            .n17537(n17537), .n16844(n16844), .n17641(n17641), .n17636(n17636), 
            .n17631(n17631), .n16828(n16828), .tx_active(tx_active), .n29(n29), 
            .n22(n22_adj_2164), .n16886(n16886), .n17573(n17573), .n17494(n17494), 
            .n8730(n8730), .tx_active_prev(tx_active_prev), .n65(n65), 
            .n17484(n17484), .n17461(n17461), .n17542(n17542), .VCC_net(VCC_net), 
            .n15701(n15701), .n10580(n10580), .n10579(n10579), .n10578(n10578), 
            .tx_o(tx_o), .n445(n445), .n9406(n9406), .n4(n4), .n12(n12), 
            .n16627(n16627), .n16629(n16629), .n9937(n9937), .n16683(n16683), 
            .n16681(n16681), .n17395(n17395), .n17394(n17394), .n16679(n16679), 
            .n16639(n16639), .n16533(n16533), .n17397(n17397), .n17398(n17398), 
            .tx_enable(tx_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(259[10:70])
    uart_tx_U0 tx2 (.r_Bit_Index({r_Bit_Index}), .GND_net(GND_net), .r_SM_Main({r_SM_Main_adj_41}), 
            .n3(n3_adj_12), .\r_SM_Main_2__N_2036[0] (r_SM_Main_2__N_2036_adj_2400[0]), 
            .\r_SM_Main_2__N_2033[1] (\r_SM_Main_2__N_2033[1] ), .n7866(n7866), 
            .n16463(n16463), .r_Clock_Count({r_Clock_Count_adj_42}), .CLK_c(CLK_c), 
            .\byte_transmit_counter2[2] (byte_transmit_counter2[2]), .\byte_transmit_counter2[4] (byte_transmit_counter2[4]), 
            .\byte_transmit_counter2[3] (byte_transmit_counter2[3]), .\byte_transmit_counter2[7] (byte_transmit_counter2[7]), 
            .\byte_transmit_counter2[5] (byte_transmit_counter2[5]), .\byte_transmit_counter2[6] (byte_transmit_counter2[6]), 
            .n10714(n10714), .n10607(n10607), .tx2_data({tx2_data}), .n17458(n17458), 
            .n16824(n16824), .n17640(n17640), .n17634(n17634), .n17629(n17629), 
            .n16817(n16817), .n16677(n16677), .n17567(n17567), .n16623(n16623), 
            .VCC_net(VCC_net), .n17457(n17457), .n16675(n16675), .n17570(n17570), 
            .n17504(n17504), .n17544(n17544), .n16673(n16673), .n16577(n16577), 
            .n16517(n16517), .n9403(n9403), .n16483(n16483), .n10587(n10587), 
            .n10585(n10585), .tx2_o(tx2_o), .n15837(n15837), .n16473(n16473), 
            .n10396(n10396), .n10399(n10399), .n9929(n9929), .n12(n12_adj_22), 
            .tx2_transmit_N_1997(tx2_transmit_N_1997), .n491(n491), .n5029(n5029), 
            .n17194(n17194), .n10398(n10398), .n15689(n15689), .tx2_enable(tx2_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(414[10:77])
    uart_rx rx (.r_Rx_Data(r_Rx_Data), .r_SM_Main({r_SM_Main_adj_43}), .n1(n1), 
            .GND_net(GND_net), .r_Clock_Count({r_Clock_Count_adj_44}), .n16863(n16863), 
            .CLK_c(CLK_c), .n16575(n16575), .n17222(n17222), .n16573(n16573), 
            .n16571(n16571), .r_Bit_Index({r_Bit_Index_adj_45}), .n13082(n13082), 
            .n4(n4_adj_37), .n16569(n16569), .n4_adj_1(n4_adj_38), .n9472(n9472), 
            .n16515(n16515), .n16479(n16479), .n16469(n16469), .n13510(n13510), 
            .rx_i(rx_i), .n10631(n10631), .rx_data_ready(rx_data_ready), 
            .n16547(n16547), .VCC_net(VCC_net), .n16855(n16855), .n16852(n16852), 
            .n16856(n16856), .n16857(n16857), .n16854(n16854), .n16858(n16858), 
            .n16860(n16860), .n16853(n16853), .n10635(n10635), .rx_data({rx_data}), 
            .n16859(n16859), .n4_adj_2(n4_adj_39), .n17260(n17260), .n17889(n17889), 
            .n17602(n17602), .n17601(n17601), .n10581(n10581), .n9477(n9477), 
            .n4_adj_3(n4_adj_40), .n6(n6), .n10423(n10423), .n10426(n10426), 
            .n16867(n16867), .n10433(n10433), .n10432(n10432), .n10431(n10431), 
            .n10430(n10430), .n10429(n10429), .n10428(n10428), .n10427(n10427), 
            .n13440(n13440), .n10425(n10425)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(386[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_SM_Main, n3, GND_net, \r_Bit_Index[1] , n14060, 
            \r_SM_Main_2__N_2036[0] , n5, n13276, n16671, r_Clock_Count, 
            CLK_c, n16651, n16649, n16567, n16509, n16477, n16467, 
            n16459, n16595, r_Tx_Data, n16625, n17537, n16844, n17641, 
            n17636, n17631, n16828, tx_active, n29, n22, n16886, 
            n17573, n17494, n8730, tx_active_prev, n65, n17484, 
            n17461, n17542, VCC_net, n15701, n10580, n10579, n10578, 
            tx_o, n445, n9406, n4, n12, n16627, n16629, n9937, 
            n16683, n16681, n17395, n17394, n16679, n16639, n16533, 
            n17397, n17398, tx_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [2:0]r_SM_Main;
    output n3;
    input GND_net;
    output \r_Bit_Index[1] ;
    output n14060;
    input \r_SM_Main_2__N_2036[0] ;
    output n5;
    output n13276;
    input n16671;
    output [8:0]r_Clock_Count;
    input CLK_c;
    input n16651;
    input n16649;
    input n16567;
    input n16509;
    input n16477;
    input n16467;
    input n16459;
    input n16595;
    output [7:0]r_Tx_Data;
    input n16625;
    output n17537;
    input n16844;
    output n17641;
    output n17636;
    output n17631;
    input n16828;
    output tx_active;
    input n29;
    input n22;
    output n16886;
    output n17573;
    output n17494;
    output n8730;
    input tx_active_prev;
    output n65;
    output n17484;
    output n17461;
    output n17542;
    input VCC_net;
    output n15701;
    input n10580;
    input n10579;
    input n10578;
    output tx_o;
    output n445;
    output n9406;
    output n4;
    output n12;
    input n16627;
    input n16629;
    output n9937;
    input n16683;
    input n16681;
    input n17395;
    input n17394;
    input n16679;
    input n16639;
    input n16533;
    input n17397;
    input n17398;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire o_Tx_Serial_N_2064;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n17462, n14082, n16539, n10872, n15683, n10873, n10712, 
        n15667, n15666, n15665, n15664, n10434, n15663, n15662, 
        n15661, n15660, n10, n17975;
    
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2064), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i15371_4_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[0]), .I2(\r_Bit_Index[1] ), 
            .I3(n14060), .O(n17462));   // verilog/uart_tx.v(31[16:25])
    defparam i15371_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9_3_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(n17462), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n5));   // verilog/uart_tx.v(31[16:25])
    defparam i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14754_4_lut (.I0(n14060), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n14082));
    defparam i14754_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i12_3_lut (.I0(n14082), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n16539));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 i10933_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n13276));
    defparam i10933_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11808_4_lut (.I0(n14082), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(\r_Bit_Index[1] ), .O(n10872));   // verilog/uart_tx.v(31[16:25])
    defparam i11808_4_lut.LUT_INIT = 16'hba40;
    SB_LUT4 i13245_2_lut (.I0(r_Bit_Index[0]), .I1(\r_Bit_Index[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n15683));   // verilog/uart_tx.v(33[16:27])
    defparam i13245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11800_4_lut (.I0(n14082), .I1(r_SM_Main[1]), .I2(r_Bit_Index[2]), 
            .I3(n15683), .O(n10873));   // verilog/uart_tx.v(31[16:25])
    defparam i11800_4_lut.LUT_INIT = 16'ha4e0;
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n16671));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n10712));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n16651));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n16649));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n16567));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n16509));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .D(n16477));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n16467));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .D(n16459));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .D(n16595));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n16539));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .D(n16625));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(n16844), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n15667), .O(n17537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_59_9_lut (.I0(n16844), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n15666), .O(n17641)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_9 (.CI(n15666), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n15667));
    SB_LUT4 add_59_8_lut (.I0(n16844), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n15665), .O(n17636)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_8 (.CI(n15665), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n15666));
    SB_LUT4 add_59_7_lut (.I0(n16828), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n15664), .O(n17631)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_7 (.CI(n15664), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n15665));
    SB_LUT4 i1_3_lut_4_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_2036[0] ), 
            .I2(n29), .I3(n22), .O(n16886));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n14060), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n10434));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 add_59_6_lut (.I0(n16828), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n15663), .O(n17573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_6 (.CI(n15663), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n15664));
    SB_LUT4 add_59_5_lut (.I0(n16828), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n15662), .O(n17494)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n8730));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut (.I0(tx_active), .I1(tx_active_prev), .I2(GND_net), 
            .I3(GND_net), .O(n65));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_59_5 (.CI(n15662), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n15663));
    SB_LUT4 add_59_4_lut (.I0(n16828), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n15661), .O(n17484)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_4 (.CI(n15661), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n15662));
    SB_LUT4 add_59_3_lut (.I0(n16828), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n15660), .O(n17461)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_3 (.CI(n15660), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n15661));
    SB_LUT4 add_59_2_lut (.I0(n16828), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n17542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n15660));
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[4]), 
            .I3(r_Clock_Count[3]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n15701));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n10580));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n10579));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .D(n10578));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut_adj_400 (.I0(tx_active), .I1(\r_SM_Main_2__N_2036[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n445));
    defparam i1_2_lut_adj_400.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_401 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n9406));
    defparam i1_2_lut_adj_401.LUT_INIT = 16'h2222;
    SB_LUT4 i8352_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n14060), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n10712));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i8352_3_lut_4_lut.LUT_INIT = 16'h0078;
    SB_LUT4 i15400_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(n14060), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2036[0] ), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15400_3_lut_4_lut_4_lut.LUT_INIT = 16'h8580;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(n15701), .O(n14060));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_402 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n12));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_4_lut_adj_402.LUT_INIT = 16'h0100;
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .D(n16627));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .D(n16629));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_2_lut_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n9937));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .D(n16683));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .D(n16681));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 n17975_bdd_4_lut (.I0(n17975), .I1(n17395), .I2(n17394), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_2064));
    defparam n17975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .D(n16679));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .D(n16639));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .D(n16533));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n10873));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(\r_Bit_Index[1] ), .C(CLK_c), .D(n10872));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(n17397), 
            .I2(n17398), .I3(r_Bit_Index[2]), .O(n17975));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n10434));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_tx_U0
//

module uart_tx_U0 (r_Bit_Index, GND_net, r_SM_Main, n3, \r_SM_Main_2__N_2036[0] , 
            \r_SM_Main_2__N_2033[1] , n7866, n16463, r_Clock_Count, 
            CLK_c, \byte_transmit_counter2[2] , \byte_transmit_counter2[4] , 
            \byte_transmit_counter2[3] , \byte_transmit_counter2[7] , \byte_transmit_counter2[5] , 
            \byte_transmit_counter2[6] , n10714, n10607, tx2_data, n17458, 
            n16824, n17640, n17634, n17629, n16817, n16677, n17567, 
            n16623, VCC_net, n17457, n16675, n17570, n17504, n17544, 
            n16673, n16577, n16517, n9403, n16483, n10587, n10585, 
            tx2_o, n15837, n16473, n10396, n10399, n9929, n12, 
            tx2_transmit_N_1997, n491, n5029, n17194, n10398, n15689, 
            tx2_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [2:0]r_Bit_Index;
    input GND_net;
    output [2:0]r_SM_Main;
    output n3;
    input \r_SM_Main_2__N_2036[0] ;
    output \r_SM_Main_2__N_2033[1] ;
    output n7866;
    input n16463;
    output [8:0]r_Clock_Count;
    input CLK_c;
    input \byte_transmit_counter2[2] ;
    input \byte_transmit_counter2[4] ;
    input \byte_transmit_counter2[3] ;
    input \byte_transmit_counter2[7] ;
    input \byte_transmit_counter2[5] ;
    input \byte_transmit_counter2[6] ;
    input n10714;
    input n10607;
    input [7:0]tx2_data;
    output n17458;
    input n16824;
    output n17640;
    output n17634;
    output n17629;
    input n16817;
    input n16677;
    output n17567;
    input n16623;
    input VCC_net;
    output n17457;
    input n16675;
    output n17570;
    output n17504;
    output n17544;
    input n16673;
    input n16577;
    input n16517;
    output n9403;
    input n16483;
    input n10587;
    input n10585;
    output tx2_o;
    output n15837;
    input n16473;
    input n10396;
    input n10399;
    output n9929;
    output n12;
    output tx2_transmit_N_1997;
    output n491;
    output n5029;
    output n17194;
    output n10398;
    input n15689;
    output tx2_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n18116, n17906, o_Tx_Serial_N_2064, n6480, n1, n10101, 
        tx2_active, n10586, n13281, n89, n113, n8737;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n18113, n15682, n15681, n15680, n15679, n15678, n15677, 
        n15676, n15675, n17903, n10;
    
    SB_LUT4 i11207211_i1_3_lut (.I0(n18116), .I1(n17906), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_2064));
    defparam i11207211_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2064), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n6480), .I2(n1), .I3(r_SM_Main[1]), 
            .O(n10101));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i10194_3_lut (.I0(n10101), .I1(r_SM_Main[1]), .I2(tx2_active), 
            .I3(GND_net), .O(n10586));   // verilog/uart_tx.v(31[16:25])
    defparam i10194_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i5592_4_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(n13281), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2033[1] ), .O(n7866));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5592_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .D(n16463));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut (.I0(\byte_transmit_counter2[2] ), .I1(\byte_transmit_counter2[4] ), 
            .I2(\byte_transmit_counter2[3] ), .I3(GND_net), .O(n89));   // coms.v(409[12:34])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i3_4_lut (.I0(n89), .I1(\byte_transmit_counter2[7] ), .I2(\byte_transmit_counter2[5] ), 
            .I3(\byte_transmit_counter2[6] ), .O(n113));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n10714));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10607));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n8737), .D(tx2_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n18113));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n18113_bdd_4_lut (.I0(n18113), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n18116));
    defparam n18113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_59_10_lut (.I0(n16824), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n15682), .O(n17458)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_59_9_lut (.I0(n16824), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n15681), .O(n17640)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_9 (.CI(n15681), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n15682));
    SB_LUT4 add_59_8_lut (.I0(n16824), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n15680), .O(n17634)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_8 (.CI(n15680), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n15681));
    SB_LUT4 add_59_7_lut (.I0(n16817), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n15679), .O(n17629)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n16677));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_7 (.CI(n15679), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n15680));
    SB_LUT4 add_59_6_lut (.I0(n16817), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n15678), .O(n17567)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_6 (.CI(n15678), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n15679));
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(VCC_net), 
            .D(n16623));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_5_lut (.I0(n16817), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n15677), .O(n17457)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n16675));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_5 (.CI(n15677), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n15678));
    SB_LUT4 add_59_4_lut (.I0(n16817), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n15676), .O(n17570)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_4 (.CI(n15676), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n15677));
    SB_LUT4 add_59_3_lut (.I0(n16817), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n15675), .O(n17504)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_3 (.CI(n15675), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n15676));
    SB_LUT4 add_59_2_lut (.I0(n16817), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n17544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n16673));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n15675));
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_15631 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n17903));
    defparam r_Bit_Index_0__bdd_4_lut_15631.LUT_INIT = 16'he4aa;
    SB_LUT4 n17903_bdd_4_lut (.I0(n17903), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n17906));
    defparam n17903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n13281));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n16577));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n16517));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n9403));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .D(n16483));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n8737));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n10587));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx2_active), .C(CLK_c), .D(n10586));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx2_o), .C(CLK_c), .D(n10585));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[4]), 
            .I3(r_Clock_Count[3]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[1]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n15837));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10646_2_lut (.I0(\r_SM_Main_2__N_2033[1] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i10646_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4216_2_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6480));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i4216_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n8737), .D(tx2_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n8737), .D(tx2_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n8737), .D(tx2_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n8737), .D(tx2_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n8737), .D(tx2_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n8737), .D(tx2_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n8737), .D(tx2_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n16473));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n10396));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .D(n10399));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_2_lut_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n9929));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_SM_Main[0]), .O(n12));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_adj_399 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(n15837), .O(\r_SM_Main_2__N_2033[1] ));
    defparam i1_2_lut_4_lut_adj_399.LUT_INIT = 16'hfffe;
    SB_LUT4 i15437_2_lut_3_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(tx2_active), 
            .I2(n113), .I3(GND_net), .O(tx2_transmit_N_1997));
    defparam i15437_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main_2__N_2036[0] ), .I1(tx2_active), 
            .I2(n113), .I3(GND_net), .O(n491));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2595_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5029));   // verilog/uart_tx.v(98[36:51])
    defparam i2595_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14756_4_lut (.I0(\r_SM_Main_2__N_2033[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n17194));
    defparam i14756_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i14834_3_lut (.I0(n17194), .I1(n13281), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n10398));
    defparam i14834_3_lut.LUT_INIT = 16'hbaba;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n15689));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx2_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx2_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (r_Rx_Data, r_SM_Main, n1, GND_net, r_Clock_Count, 
            n16863, CLK_c, n16575, n17222, n16573, n16571, r_Bit_Index, 
            n13082, n4, n16569, n4_adj_1, n9472, n16515, n16479, 
            n16469, n13510, rx_i, n10631, rx_data_ready, n16547, 
            VCC_net, n16855, n16852, n16856, n16857, n16854, n16858, 
            n16860, n16853, n10635, rx_data, n16859, n4_adj_2, n17260, 
            n17889, n17602, n17601, n10581, n9477, n4_adj_3, n6, 
            n10423, n10426, n16867, n10433, n10432, n10431, n10430, 
            n10429, n10428, n10427, n13440, n10425) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output r_Rx_Data;
    output [2:0]r_SM_Main;
    output n1;
    input GND_net;
    output [7:0]r_Clock_Count;
    output n16863;
    input CLK_c;
    input n16575;
    output n17222;
    input n16573;
    input n16571;
    output [2:0]r_Bit_Index;
    output n13082;
    output n4;
    input n16569;
    output n4_adj_1;
    output n9472;
    input n16515;
    input n16479;
    input n16469;
    input n13510;
    input rx_i;
    input n10631;
    output rx_data_ready;
    input n16547;
    input VCC_net;
    output n16855;
    input n16852;
    output n16856;
    output n16857;
    output n16854;
    output n16858;
    output n16860;
    output n16853;
    input n10635;
    output [7:0]rx_data;
    output n16859;
    output n4_adj_2;
    output n17260;
    output n17889;
    output n17602;
    output n17601;
    input n10581;
    output n9477;
    output n4_adj_3;
    output n6;
    input n10423;
    input n10426;
    output n16867;
    input n10433;
    input n10432;
    input n10431;
    input n10430;
    input n10429;
    input n10428;
    input n10427;
    output n13440;
    output n10425;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_SM_Main_2__N_2096;
    
    wire n6_c;
    wire [2:0]r_SM_Main_2__N_2090;
    
    wire n16850, n13452, n9323, r_Rx_Data_R, n16501, n15674, n15673, 
        n15672, n15671, n15670, n15669, n15668, n10086;
    
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2096[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(n6_c), 
            .I3(r_Clock_Count[3]), .O(n16863));
    defparam i1_4_lut.LUT_INIT = 16'h8000;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(r_SM_Main_2__N_2090[2]), 
            .R(n16850));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n16575));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i14784_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17222));
    defparam i14784_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11107_2_lut (.I0(r_Clock_Count[5]), .I1(n16863), .I2(GND_net), 
            .I3(GND_net), .O(n13452));
    defparam i11107_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n16573));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n16571));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i10739_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n13082));
    defparam i10739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_52_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_52_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n16569));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_54_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_54_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n9323), .I1(r_Bit_Index[0]), .I2(GND_net), .I3(GND_net), 
            .O(n9472));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n16515));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .D(n16479));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n16469));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n13510));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(rx_i));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n10631));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n16501));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(VCC_net), 
            .D(n16547));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(n16852), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n15674), .O(n16855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n16852), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n15673), .O(n16856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n15673), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n15674));
    SB_LUT4 add_62_7_lut (.I0(n16852), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n15672), .O(n16857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n15672), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n15673));
    SB_LUT4 add_62_6_lut (.I0(n16852), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n15671), .O(n16854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n15671), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n15672));
    SB_LUT4 add_62_5_lut (.I0(n16852), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n15670), .O(n16858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n15670), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n15671));
    SB_LUT4 add_62_4_lut (.I0(n16852), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n15669), .O(n16860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n15669), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n15670));
    SB_LUT4 add_62_3_lut (.I0(n16852), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n15668), .O(n16853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n15668), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n15669));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n10635));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_2_lut (.I0(n16852), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n16859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n15668));
    SB_LUT4 i1_2_lut_adj_395 (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));
    defparam i1_2_lut_adj_395.LUT_INIT = 16'h8888;
    SB_LUT4 i14822_4_lut (.I0(r_SM_Main_2__N_2090[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n17260));
    defparam i14822_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(n16863), .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_2096[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i15448_1_lut (.I0(rx_data_ready), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17889));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15448_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15361_2_lut (.I0(r_SM_Main_2__N_2090[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n17602));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15303_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_2096[0]), 
            .I3(GND_net), .O(n17601));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i15303_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n10581));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_2090[2]), .O(n9323));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i2_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_396 (.I0(r_Bit_Index[0]), .I1(n9323), .I2(GND_net), 
            .I3(GND_net), .O(n9477));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_396.LUT_INIT = 16'heeee;
    SB_LUT4 equal_56_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3));   // verilog/uart_rx.v(97[17:39])
    defparam equal_56_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_397 (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2096[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_397.LUT_INIT = 16'h2222;
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .D(n10423));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .D(n10426));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut_4_lut_adj_398 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(n13452), .I3(n17222), .O(n16867));
    defparam i2_3_lut_4_lut_adj_398.LUT_INIT = 16'h0004;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_2090[2]), 
            .I3(r_SM_Main[0]), .O(n10086));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h4033;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n10086), 
            .I3(rx_data_ready), .O(n16501));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n10433));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n10432));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n10431));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n10430));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n10429));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n10428));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n10427));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i15447_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n16850));
    defparam i15447_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[5]), .I1(n16863), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(r_SM_Main_2__N_2090[2]));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff8;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut (.I0(r_Bit_Index[2]), 
            .I1(n4_adj_2), .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_2090[2]), 
            .O(n13440));
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut.LUT_INIT = 16'hf70f;
    SB_LUT4 i14832_3_lut_4_lut (.I0(r_Bit_Index[2]), .I1(n4_adj_2), .I2(r_SM_Main[1]), 
            .I3(n17260), .O(n10425));
    defparam i14832_3_lut_4_lut.LUT_INIT = 16'hff70;
    
endmodule
