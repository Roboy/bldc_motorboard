// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jun 29 2019 15:10:02

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    pin9,
    pin8,
    pin7,
    pin6,
    pin5,
    pin4,
    pin3_clk_16mhz,
    pin2_usb_dn,
    pin24,
    pin23,
    pin22,
    pin21,
    pin20,
    pin1_usb_dp,
    pin19,
    pin18,
    pin17_ss,
    pin16_sck,
    pin15_sdi,
    pin14_sdo,
    pin13,
    pin12,
    pin11,
    pin10);

    output pin9;
    output pin8;
    output pin7;
    input pin6;
    input pin5;
    input pin4;
    input pin3_clk_16mhz;
    output pin2_usb_dn;
    output pin24;
    output pin23;
    output pin22;
    output pin21;
    output pin20;
    output pin1_usb_dp;
    output pin19;
    output pin18;
    output pin17_ss;
    output pin16_sck;
    output pin15_sdi;
    output pin14_sdo;
    output pin13;
    output pin12;
    output pin11;
    output pin10;

    wire N__69497;
    wire N__69496;
    wire N__69495;
    wire N__69488;
    wire N__69487;
    wire N__69486;
    wire N__69479;
    wire N__69478;
    wire N__69477;
    wire N__69470;
    wire N__69469;
    wire N__69468;
    wire N__69461;
    wire N__69460;
    wire N__69459;
    wire N__69452;
    wire N__69451;
    wire N__69450;
    wire N__69443;
    wire N__69442;
    wire N__69441;
    wire N__69434;
    wire N__69433;
    wire N__69432;
    wire N__69425;
    wire N__69424;
    wire N__69423;
    wire N__69416;
    wire N__69415;
    wire N__69414;
    wire N__69407;
    wire N__69406;
    wire N__69405;
    wire N__69398;
    wire N__69397;
    wire N__69396;
    wire N__69389;
    wire N__69388;
    wire N__69387;
    wire N__69380;
    wire N__69379;
    wire N__69378;
    wire N__69371;
    wire N__69370;
    wire N__69369;
    wire N__69362;
    wire N__69361;
    wire N__69360;
    wire N__69353;
    wire N__69352;
    wire N__69351;
    wire N__69344;
    wire N__69343;
    wire N__69342;
    wire N__69335;
    wire N__69334;
    wire N__69333;
    wire N__69326;
    wire N__69325;
    wire N__69324;
    wire N__69317;
    wire N__69316;
    wire N__69315;
    wire N__69298;
    wire N__69295;
    wire N__69294;
    wire N__69293;
    wire N__69288;
    wire N__69285;
    wire N__69282;
    wire N__69279;
    wire N__69276;
    wire N__69273;
    wire N__69268;
    wire N__69265;
    wire N__69262;
    wire N__69259;
    wire N__69256;
    wire N__69253;
    wire N__69252;
    wire N__69251;
    wire N__69246;
    wire N__69243;
    wire N__69240;
    wire N__69237;
    wire N__69234;
    wire N__69231;
    wire N__69226;
    wire N__69223;
    wire N__69220;
    wire N__69217;
    wire N__69214;
    wire N__69211;
    wire N__69208;
    wire N__69205;
    wire N__69204;
    wire N__69203;
    wire N__69200;
    wire N__69197;
    wire N__69194;
    wire N__69191;
    wire N__69186;
    wire N__69183;
    wire N__69180;
    wire N__69175;
    wire N__69172;
    wire N__69169;
    wire N__69166;
    wire N__69163;
    wire N__69160;
    wire N__69157;
    wire N__69156;
    wire N__69155;
    wire N__69150;
    wire N__69147;
    wire N__69144;
    wire N__69141;
    wire N__69136;
    wire N__69133;
    wire N__69130;
    wire N__69127;
    wire N__69124;
    wire N__69121;
    wire N__69118;
    wire N__69115;
    wire N__69112;
    wire N__69109;
    wire N__69108;
    wire N__69107;
    wire N__69102;
    wire N__69099;
    wire N__69096;
    wire N__69093;
    wire N__69090;
    wire N__69087;
    wire N__69084;
    wire N__69081;
    wire N__69076;
    wire N__69073;
    wire N__69072;
    wire N__69071;
    wire N__69068;
    wire N__69067;
    wire N__69064;
    wire N__69063;
    wire N__69060;
    wire N__69059;
    wire N__69046;
    wire N__69045;
    wire N__69044;
    wire N__69043;
    wire N__69040;
    wire N__69037;
    wire N__69032;
    wire N__69025;
    wire N__69022;
    wire N__69019;
    wire N__69016;
    wire N__69013;
    wire N__69010;
    wire N__69007;
    wire N__69006;
    wire N__69003;
    wire N__69000;
    wire N__68997;
    wire N__68994;
    wire N__68991;
    wire N__68988;
    wire N__68983;
    wire N__68980;
    wire N__68977;
    wire N__68974;
    wire N__68971;
    wire N__68968;
    wire N__68965;
    wire N__68962;
    wire N__68961;
    wire N__68958;
    wire N__68955;
    wire N__68952;
    wire N__68949;
    wire N__68944;
    wire N__68943;
    wire N__68942;
    wire N__68937;
    wire N__68936;
    wire N__68933;
    wire N__68930;
    wire N__68927;
    wire N__68924;
    wire N__68919;
    wire N__68914;
    wire N__68911;
    wire N__68910;
    wire N__68907;
    wire N__68904;
    wire N__68901;
    wire N__68898;
    wire N__68895;
    wire N__68890;
    wire N__68887;
    wire N__68884;
    wire N__68881;
    wire N__68878;
    wire N__68875;
    wire N__68872;
    wire N__68871;
    wire N__68866;
    wire N__68863;
    wire N__68862;
    wire N__68861;
    wire N__68858;
    wire N__68855;
    wire N__68852;
    wire N__68845;
    wire N__68842;
    wire N__68839;
    wire N__68836;
    wire N__68833;
    wire N__68830;
    wire N__68829;
    wire N__68826;
    wire N__68823;
    wire N__68818;
    wire N__68815;
    wire N__68812;
    wire N__68809;
    wire N__68806;
    wire N__68803;
    wire N__68800;
    wire N__68799;
    wire N__68794;
    wire N__68793;
    wire N__68792;
    wire N__68789;
    wire N__68786;
    wire N__68783;
    wire N__68776;
    wire N__68773;
    wire N__68770;
    wire N__68769;
    wire N__68766;
    wire N__68763;
    wire N__68760;
    wire N__68757;
    wire N__68754;
    wire N__68751;
    wire N__68746;
    wire N__68743;
    wire N__68740;
    wire N__68737;
    wire N__68734;
    wire N__68731;
    wire N__68728;
    wire N__68727;
    wire N__68722;
    wire N__68721;
    wire N__68720;
    wire N__68717;
    wire N__68714;
    wire N__68711;
    wire N__68704;
    wire N__68701;
    wire N__68698;
    wire N__68697;
    wire N__68694;
    wire N__68691;
    wire N__68688;
    wire N__68685;
    wire N__68682;
    wire N__68679;
    wire N__68674;
    wire N__68671;
    wire N__68668;
    wire N__68665;
    wire N__68662;
    wire N__68659;
    wire N__68658;
    wire N__68653;
    wire N__68650;
    wire N__68649;
    wire N__68648;
    wire N__68645;
    wire N__68642;
    wire N__68639;
    wire N__68636;
    wire N__68631;
    wire N__68626;
    wire N__68623;
    wire N__68620;
    wire N__68617;
    wire N__68614;
    wire N__68611;
    wire N__68608;
    wire N__68607;
    wire N__68602;
    wire N__68601;
    wire N__68598;
    wire N__68595;
    wire N__68594;
    wire N__68591;
    wire N__68588;
    wire N__68585;
    wire N__68582;
    wire N__68577;
    wire N__68572;
    wire N__68569;
    wire N__68566;
    wire N__68563;
    wire N__68560;
    wire N__68557;
    wire N__68554;
    wire N__68551;
    wire N__68550;
    wire N__68549;
    wire N__68546;
    wire N__68543;
    wire N__68540;
    wire N__68537;
    wire N__68534;
    wire N__68531;
    wire N__68528;
    wire N__68523;
    wire N__68518;
    wire N__68515;
    wire N__68512;
    wire N__68509;
    wire N__68506;
    wire N__68503;
    wire N__68500;
    wire N__68497;
    wire N__68496;
    wire N__68493;
    wire N__68490;
    wire N__68487;
    wire N__68484;
    wire N__68479;
    wire N__68476;
    wire N__68473;
    wire N__68470;
    wire N__68467;
    wire N__68464;
    wire N__68461;
    wire N__68460;
    wire N__68459;
    wire N__68456;
    wire N__68453;
    wire N__68450;
    wire N__68445;
    wire N__68440;
    wire N__68437;
    wire N__68436;
    wire N__68435;
    wire N__68434;
    wire N__68429;
    wire N__68428;
    wire N__68427;
    wire N__68426;
    wire N__68423;
    wire N__68422;
    wire N__68419;
    wire N__68418;
    wire N__68415;
    wire N__68412;
    wire N__68411;
    wire N__68408;
    wire N__68407;
    wire N__68404;
    wire N__68403;
    wire N__68402;
    wire N__68401;
    wire N__68400;
    wire N__68399;
    wire N__68398;
    wire N__68397;
    wire N__68396;
    wire N__68395;
    wire N__68394;
    wire N__68393;
    wire N__68392;
    wire N__68391;
    wire N__68390;
    wire N__68387;
    wire N__68384;
    wire N__68379;
    wire N__68374;
    wire N__68365;
    wire N__68364;
    wire N__68361;
    wire N__68360;
    wire N__68357;
    wire N__68356;
    wire N__68353;
    wire N__68352;
    wire N__68349;
    wire N__68348;
    wire N__68345;
    wire N__68344;
    wire N__68341;
    wire N__68340;
    wire N__68337;
    wire N__68336;
    wire N__68333;
    wire N__68332;
    wire N__68329;
    wire N__68326;
    wire N__68323;
    wire N__68320;
    wire N__68317;
    wire N__68314;
    wire N__68311;
    wire N__68306;
    wire N__68303;
    wire N__68300;
    wire N__68283;
    wire N__68266;
    wire N__68257;
    wire N__68250;
    wire N__68247;
    wire N__68244;
    wire N__68231;
    wire N__68226;
    wire N__68223;
    wire N__68218;
    wire N__68215;
    wire N__68214;
    wire N__68211;
    wire N__68208;
    wire N__68203;
    wire N__68200;
    wire N__68197;
    wire N__68194;
    wire N__68191;
    wire N__68188;
    wire N__68187;
    wire N__68184;
    wire N__68181;
    wire N__68180;
    wire N__68179;
    wire N__68174;
    wire N__68171;
    wire N__68168;
    wire N__68165;
    wire N__68162;
    wire N__68159;
    wire N__68156;
    wire N__68151;
    wire N__68146;
    wire N__68143;
    wire N__68140;
    wire N__68137;
    wire N__68136;
    wire N__68133;
    wire N__68130;
    wire N__68125;
    wire N__68122;
    wire N__68119;
    wire N__68116;
    wire N__68113;
    wire N__68110;
    wire N__68107;
    wire N__68106;
    wire N__68101;
    wire N__68100;
    wire N__68099;
    wire N__68096;
    wire N__68091;
    wire N__68086;
    wire N__68083;
    wire N__68080;
    wire N__68077;
    wire N__68076;
    wire N__68073;
    wire N__68070;
    wire N__68065;
    wire N__68062;
    wire N__68059;
    wire N__68056;
    wire N__68053;
    wire N__68050;
    wire N__68049;
    wire N__68048;
    wire N__68047;
    wire N__68042;
    wire N__68037;
    wire N__68034;
    wire N__68031;
    wire N__68028;
    wire N__68025;
    wire N__68020;
    wire N__68017;
    wire N__68014;
    wire N__68013;
    wire N__68010;
    wire N__68007;
    wire N__68004;
    wire N__68001;
    wire N__67996;
    wire N__67993;
    wire N__67990;
    wire N__67987;
    wire N__67984;
    wire N__67981;
    wire N__67978;
    wire N__67977;
    wire N__67974;
    wire N__67971;
    wire N__67970;
    wire N__67965;
    wire N__67964;
    wire N__67961;
    wire N__67958;
    wire N__67955;
    wire N__67952;
    wire N__67949;
    wire N__67946;
    wire N__67943;
    wire N__67936;
    wire N__67933;
    wire N__67930;
    wire N__67929;
    wire N__67926;
    wire N__67923;
    wire N__67918;
    wire N__67915;
    wire N__67912;
    wire N__67909;
    wire N__67906;
    wire N__67903;
    wire N__67900;
    wire N__67899;
    wire N__67898;
    wire N__67895;
    wire N__67892;
    wire N__67889;
    wire N__67886;
    wire N__67885;
    wire N__67880;
    wire N__67877;
    wire N__67874;
    wire N__67867;
    wire N__67864;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67852;
    wire N__67849;
    wire N__67846;
    wire N__67843;
    wire N__67842;
    wire N__67839;
    wire N__67836;
    wire N__67833;
    wire N__67830;
    wire N__67825;
    wire N__67822;
    wire N__67819;
    wire N__67816;
    wire N__67813;
    wire N__67810;
    wire N__67809;
    wire N__67806;
    wire N__67803;
    wire N__67798;
    wire N__67795;
    wire N__67792;
    wire N__67789;
    wire N__67786;
    wire N__67783;
    wire N__67780;
    wire N__67779;
    wire N__67776;
    wire N__67773;
    wire N__67768;
    wire N__67765;
    wire N__67762;
    wire N__67759;
    wire N__67758;
    wire N__67755;
    wire N__67752;
    wire N__67747;
    wire N__67744;
    wire N__67741;
    wire N__67738;
    wire N__67735;
    wire N__67732;
    wire N__67729;
    wire N__67728;
    wire N__67725;
    wire N__67722;
    wire N__67717;
    wire N__67714;
    wire N__67711;
    wire N__67708;
    wire N__67705;
    wire N__67702;
    wire N__67699;
    wire N__67696;
    wire N__67695;
    wire N__67692;
    wire N__67689;
    wire N__67686;
    wire N__67683;
    wire N__67678;
    wire N__67677;
    wire N__67674;
    wire N__67673;
    wire N__67670;
    wire N__67667;
    wire N__67664;
    wire N__67661;
    wire N__67654;
    wire N__67651;
    wire N__67650;
    wire N__67647;
    wire N__67644;
    wire N__67641;
    wire N__67638;
    wire N__67633;
    wire N__67630;
    wire N__67627;
    wire N__67624;
    wire N__67621;
    wire N__67618;
    wire N__67617;
    wire N__67612;
    wire N__67611;
    wire N__67610;
    wire N__67607;
    wire N__67604;
    wire N__67601;
    wire N__67596;
    wire N__67591;
    wire N__67588;
    wire N__67585;
    wire N__67582;
    wire N__67581;
    wire N__67578;
    wire N__67575;
    wire N__67570;
    wire N__67567;
    wire N__67564;
    wire N__67561;
    wire N__67558;
    wire N__67555;
    wire N__67554;
    wire N__67549;
    wire N__67548;
    wire N__67547;
    wire N__67544;
    wire N__67541;
    wire N__67538;
    wire N__67535;
    wire N__67530;
    wire N__67525;
    wire N__67522;
    wire N__67519;
    wire N__67516;
    wire N__67513;
    wire N__67510;
    wire N__67507;
    wire N__67504;
    wire N__67503;
    wire N__67500;
    wire N__67497;
    wire N__67492;
    wire N__67489;
    wire N__67486;
    wire N__67485;
    wire N__67482;
    wire N__67479;
    wire N__67474;
    wire N__67471;
    wire N__67468;
    wire N__67467;
    wire N__67466;
    wire N__67465;
    wire N__67464;
    wire N__67463;
    wire N__67462;
    wire N__67461;
    wire N__67460;
    wire N__67459;
    wire N__67458;
    wire N__67457;
    wire N__67456;
    wire N__67455;
    wire N__67452;
    wire N__67449;
    wire N__67446;
    wire N__67443;
    wire N__67442;
    wire N__67439;
    wire N__67436;
    wire N__67433;
    wire N__67430;
    wire N__67427;
    wire N__67426;
    wire N__67425;
    wire N__67422;
    wire N__67421;
    wire N__67418;
    wire N__67417;
    wire N__67414;
    wire N__67413;
    wire N__67410;
    wire N__67409;
    wire N__67406;
    wire N__67405;
    wire N__67404;
    wire N__67401;
    wire N__67398;
    wire N__67397;
    wire N__67396;
    wire N__67395;
    wire N__67392;
    wire N__67389;
    wire N__67386;
    wire N__67381;
    wire N__67372;
    wire N__67355;
    wire N__67352;
    wire N__67351;
    wire N__67348;
    wire N__67345;
    wire N__67342;
    wire N__67337;
    wire N__67334;
    wire N__67331;
    wire N__67328;
    wire N__67323;
    wire N__67320;
    wire N__67315;
    wire N__67312;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67300;
    wire N__67297;
    wire N__67296;
    wire N__67293;
    wire N__67290;
    wire N__67287;
    wire N__67284;
    wire N__67279;
    wire N__67272;
    wire N__67269;
    wire N__67262;
    wire N__67259;
    wire N__67254;
    wire N__67243;
    wire N__67240;
    wire N__67237;
    wire N__67234;
    wire N__67227;
    wire N__67224;
    wire N__67221;
    wire N__67216;
    wire N__67213;
    wire N__67210;
    wire N__67207;
    wire N__67204;
    wire N__67203;
    wire N__67200;
    wire N__67197;
    wire N__67192;
    wire N__67189;
    wire N__67186;
    wire N__67183;
    wire N__67180;
    wire N__67177;
    wire N__67174;
    wire N__67171;
    wire N__67168;
    wire N__67165;
    wire N__67162;
    wire N__67161;
    wire N__67158;
    wire N__67155;
    wire N__67150;
    wire N__67147;
    wire N__67144;
    wire N__67141;
    wire N__67138;
    wire N__67135;
    wire N__67132;
    wire N__67129;
    wire N__67126;
    wire N__67123;
    wire N__67120;
    wire N__67117;
    wire N__67116;
    wire N__67113;
    wire N__67110;
    wire N__67105;
    wire N__67102;
    wire N__67099;
    wire N__67096;
    wire N__67093;
    wire N__67090;
    wire N__67087;
    wire N__67084;
    wire N__67081;
    wire N__67078;
    wire N__67077;
    wire N__67074;
    wire N__67071;
    wire N__67066;
    wire N__67063;
    wire N__67060;
    wire N__67057;
    wire N__67054;
    wire N__67051;
    wire N__67048;
    wire N__67045;
    wire N__67042;
    wire N__67039;
    wire N__67036;
    wire N__67033;
    wire N__67032;
    wire N__67029;
    wire N__67026;
    wire N__67021;
    wire N__67018;
    wire N__67015;
    wire N__67012;
    wire N__67009;
    wire N__67006;
    wire N__67003;
    wire N__67000;
    wire N__66997;
    wire N__66994;
    wire N__66991;
    wire N__66988;
    wire N__66985;
    wire N__66982;
    wire N__66979;
    wire N__66976;
    wire N__66973;
    wire N__66970;
    wire N__66967;
    wire N__66964;
    wire N__66961;
    wire N__66958;
    wire N__66955;
    wire N__66952;
    wire N__66949;
    wire N__66946;
    wire N__66943;
    wire N__66940;
    wire N__66937;
    wire N__66934;
    wire N__66931;
    wire N__66930;
    wire N__66929;
    wire N__66928;
    wire N__66927;
    wire N__66926;
    wire N__66925;
    wire N__66924;
    wire N__66923;
    wire N__66922;
    wire N__66921;
    wire N__66920;
    wire N__66917;
    wire N__66914;
    wire N__66913;
    wire N__66910;
    wire N__66907;
    wire N__66904;
    wire N__66901;
    wire N__66898;
    wire N__66895;
    wire N__66892;
    wire N__66891;
    wire N__66890;
    wire N__66889;
    wire N__66888;
    wire N__66885;
    wire N__66884;
    wire N__66881;
    wire N__66880;
    wire N__66877;
    wire N__66876;
    wire N__66875;
    wire N__66870;
    wire N__66861;
    wire N__66852;
    wire N__66849;
    wire N__66846;
    wire N__66843;
    wire N__66840;
    wire N__66837;
    wire N__66834;
    wire N__66831;
    wire N__66830;
    wire N__66829;
    wire N__66828;
    wire N__66825;
    wire N__66824;
    wire N__66823;
    wire N__66822;
    wire N__66819;
    wire N__66816;
    wire N__66813;
    wire N__66808;
    wire N__66805;
    wire N__66796;
    wire N__66789;
    wire N__66786;
    wire N__66783;
    wire N__66782;
    wire N__66779;
    wire N__66776;
    wire N__66773;
    wire N__66770;
    wire N__66767;
    wire N__66764;
    wire N__66761;
    wire N__66760;
    wire N__66757;
    wire N__66750;
    wire N__66747;
    wire N__66744;
    wire N__66741;
    wire N__66738;
    wire N__66735;
    wire N__66732;
    wire N__66729;
    wire N__66726;
    wire N__66723;
    wire N__66720;
    wire N__66717;
    wire N__66714;
    wire N__66711;
    wire N__66708;
    wire N__66705;
    wire N__66698;
    wire N__66695;
    wire N__66688;
    wire N__66685;
    wire N__66676;
    wire N__66673;
    wire N__66668;
    wire N__66663;
    wire N__66658;
    wire N__66649;
    wire N__66646;
    wire N__66643;
    wire N__66640;
    wire N__66639;
    wire N__66638;
    wire N__66635;
    wire N__66632;
    wire N__66631;
    wire N__66630;
    wire N__66629;
    wire N__66626;
    wire N__66625;
    wire N__66622;
    wire N__66619;
    wire N__66616;
    wire N__66613;
    wire N__66612;
    wire N__66609;
    wire N__66608;
    wire N__66605;
    wire N__66604;
    wire N__66601;
    wire N__66600;
    wire N__66599;
    wire N__66598;
    wire N__66595;
    wire N__66592;
    wire N__66589;
    wire N__66586;
    wire N__66583;
    wire N__66580;
    wire N__66577;
    wire N__66576;
    wire N__66575;
    wire N__66574;
    wire N__66571;
    wire N__66568;
    wire N__66565;
    wire N__66562;
    wire N__66559;
    wire N__66556;
    wire N__66549;
    wire N__66542;
    wire N__66539;
    wire N__66538;
    wire N__66535;
    wire N__66534;
    wire N__66531;
    wire N__66528;
    wire N__66525;
    wire N__66522;
    wire N__66521;
    wire N__66520;
    wire N__66519;
    wire N__66518;
    wire N__66517;
    wire N__66516;
    wire N__66515;
    wire N__66512;
    wire N__66509;
    wire N__66506;
    wire N__66503;
    wire N__66496;
    wire N__66493;
    wire N__66486;
    wire N__66483;
    wire N__66478;
    wire N__66475;
    wire N__66472;
    wire N__66469;
    wire N__66468;
    wire N__66465;
    wire N__66464;
    wire N__66461;
    wire N__66458;
    wire N__66455;
    wire N__66448;
    wire N__66445;
    wire N__66442;
    wire N__66435;
    wire N__66432;
    wire N__66429;
    wire N__66416;
    wire N__66411;
    wire N__66408;
    wire N__66393;
    wire N__66388;
    wire N__66385;
    wire N__66382;
    wire N__66379;
    wire N__66376;
    wire N__66373;
    wire N__66370;
    wire N__66367;
    wire N__66364;
    wire N__66361;
    wire N__66360;
    wire N__66359;
    wire N__66356;
    wire N__66353;
    wire N__66350;
    wire N__66349;
    wire N__66348;
    wire N__66347;
    wire N__66346;
    wire N__66345;
    wire N__66344;
    wire N__66343;
    wire N__66340;
    wire N__66337;
    wire N__66334;
    wire N__66331;
    wire N__66328;
    wire N__66327;
    wire N__66324;
    wire N__66321;
    wire N__66318;
    wire N__66315;
    wire N__66312;
    wire N__66307;
    wire N__66304;
    wire N__66301;
    wire N__66298;
    wire N__66295;
    wire N__66294;
    wire N__66293;
    wire N__66290;
    wire N__66287;
    wire N__66286;
    wire N__66283;
    wire N__66280;
    wire N__66277;
    wire N__66268;
    wire N__66265;
    wire N__66262;
    wire N__66261;
    wire N__66260;
    wire N__66259;
    wire N__66256;
    wire N__66253;
    wire N__66250;
    wire N__66247;
    wire N__66244;
    wire N__66235;
    wire N__66232;
    wire N__66229;
    wire N__66226;
    wire N__66221;
    wire N__66220;
    wire N__66219;
    wire N__66218;
    wire N__66217;
    wire N__66214;
    wire N__66211;
    wire N__66208;
    wire N__66201;
    wire N__66198;
    wire N__66193;
    wire N__66192;
    wire N__66189;
    wire N__66188;
    wire N__66185;
    wire N__66184;
    wire N__66181;
    wire N__66180;
    wire N__66177;
    wire N__66174;
    wire N__66169;
    wire N__66166;
    wire N__66163;
    wire N__66160;
    wire N__66143;
    wire N__66140;
    wire N__66137;
    wire N__66132;
    wire N__66127;
    wire N__66118;
    wire N__66115;
    wire N__66112;
    wire N__66109;
    wire N__66106;
    wire N__66103;
    wire N__66100;
    wire N__66099;
    wire N__66098;
    wire N__66095;
    wire N__66094;
    wire N__66093;
    wire N__66092;
    wire N__66091;
    wire N__66090;
    wire N__66087;
    wire N__66086;
    wire N__66083;
    wire N__66080;
    wire N__66077;
    wire N__66074;
    wire N__66071;
    wire N__66070;
    wire N__66067;
    wire N__66064;
    wire N__66063;
    wire N__66060;
    wire N__66057;
    wire N__66056;
    wire N__66053;
    wire N__66050;
    wire N__66047;
    wire N__66044;
    wire N__66041;
    wire N__66040;
    wire N__66037;
    wire N__66036;
    wire N__66033;
    wire N__66032;
    wire N__66031;
    wire N__66030;
    wire N__66029;
    wire N__66028;
    wire N__66025;
    wire N__66022;
    wire N__66019;
    wire N__66016;
    wire N__66013;
    wire N__66012;
    wire N__66005;
    wire N__66002;
    wire N__65999;
    wire N__65996;
    wire N__65993;
    wire N__65990;
    wire N__65987;
    wire N__65984;
    wire N__65983;
    wire N__65980;
    wire N__65979;
    wire N__65976;
    wire N__65975;
    wire N__65972;
    wire N__65969;
    wire N__65966;
    wire N__65963;
    wire N__65958;
    wire N__65955;
    wire N__65952;
    wire N__65941;
    wire N__65938;
    wire N__65935;
    wire N__65928;
    wire N__65917;
    wire N__65914;
    wire N__65911;
    wire N__65908;
    wire N__65905;
    wire N__65902;
    wire N__65897;
    wire N__65890;
    wire N__65887;
    wire N__65884;
    wire N__65877;
    wire N__65872;
    wire N__65863;
    wire N__65860;
    wire N__65857;
    wire N__65854;
    wire N__65851;
    wire N__65848;
    wire N__65845;
    wire N__65844;
    wire N__65843;
    wire N__65840;
    wire N__65839;
    wire N__65836;
    wire N__65833;
    wire N__65832;
    wire N__65831;
    wire N__65830;
    wire N__65829;
    wire N__65828;
    wire N__65825;
    wire N__65822;
    wire N__65819;
    wire N__65816;
    wire N__65813;
    wire N__65810;
    wire N__65809;
    wire N__65808;
    wire N__65807;
    wire N__65804;
    wire N__65801;
    wire N__65798;
    wire N__65795;
    wire N__65792;
    wire N__65791;
    wire N__65786;
    wire N__65783;
    wire N__65780;
    wire N__65777;
    wire N__65776;
    wire N__65773;
    wire N__65770;
    wire N__65767;
    wire N__65764;
    wire N__65761;
    wire N__65756;
    wire N__65753;
    wire N__65746;
    wire N__65743;
    wire N__65740;
    wire N__65739;
    wire N__65738;
    wire N__65737;
    wire N__65736;
    wire N__65735;
    wire N__65734;
    wire N__65731;
    wire N__65728;
    wire N__65725;
    wire N__65718;
    wire N__65715;
    wire N__65710;
    wire N__65707;
    wire N__65704;
    wire N__65701;
    wire N__65698;
    wire N__65697;
    wire N__65694;
    wire N__65691;
    wire N__65688;
    wire N__65683;
    wire N__65680;
    wire N__65675;
    wire N__65670;
    wire N__65667;
    wire N__65662;
    wire N__65653;
    wire N__65648;
    wire N__65645;
    wire N__65636;
    wire N__65629;
    wire N__65626;
    wire N__65623;
    wire N__65620;
    wire N__65617;
    wire N__65614;
    wire N__65611;
    wire N__65610;
    wire N__65609;
    wire N__65606;
    wire N__65603;
    wire N__65602;
    wire N__65601;
    wire N__65600;
    wire N__65597;
    wire N__65596;
    wire N__65595;
    wire N__65592;
    wire N__65589;
    wire N__65586;
    wire N__65583;
    wire N__65582;
    wire N__65581;
    wire N__65580;
    wire N__65577;
    wire N__65574;
    wire N__65571;
    wire N__65570;
    wire N__65567;
    wire N__65562;
    wire N__65559;
    wire N__65556;
    wire N__65553;
    wire N__65550;
    wire N__65547;
    wire N__65546;
    wire N__65543;
    wire N__65540;
    wire N__65537;
    wire N__65534;
    wire N__65531;
    wire N__65524;
    wire N__65521;
    wire N__65518;
    wire N__65515;
    wire N__65512;
    wire N__65511;
    wire N__65510;
    wire N__65509;
    wire N__65508;
    wire N__65507;
    wire N__65504;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65492;
    wire N__65483;
    wire N__65480;
    wire N__65477;
    wire N__65468;
    wire N__65467;
    wire N__65464;
    wire N__65459;
    wire N__65456;
    wire N__65453;
    wire N__65448;
    wire N__65445;
    wire N__65442;
    wire N__65439;
    wire N__65438;
    wire N__65437;
    wire N__65432;
    wire N__65427;
    wire N__65418;
    wire N__65413;
    wire N__65404;
    wire N__65401;
    wire N__65398;
    wire N__65395;
    wire N__65392;
    wire N__65389;
    wire N__65388;
    wire N__65387;
    wire N__65386;
    wire N__65385;
    wire N__65384;
    wire N__65381;
    wire N__65378;
    wire N__65375;
    wire N__65374;
    wire N__65371;
    wire N__65368;
    wire N__65365;
    wire N__65362;
    wire N__65361;
    wire N__65356;
    wire N__65353;
    wire N__65352;
    wire N__65349;
    wire N__65348;
    wire N__65343;
    wire N__65342;
    wire N__65341;
    wire N__65338;
    wire N__65335;
    wire N__65330;
    wire N__65327;
    wire N__65324;
    wire N__65321;
    wire N__65320;
    wire N__65317;
    wire N__65314;
    wire N__65313;
    wire N__65310;
    wire N__65301;
    wire N__65296;
    wire N__65293;
    wire N__65288;
    wire N__65285;
    wire N__65284;
    wire N__65281;
    wire N__65274;
    wire N__65271;
    wire N__65268;
    wire N__65265;
    wire N__65264;
    wire N__65261;
    wire N__65258;
    wire N__65251;
    wire N__65248;
    wire N__65245;
    wire N__65242;
    wire N__65239;
    wire N__65236;
    wire N__65227;
    wire N__65224;
    wire N__65221;
    wire N__65218;
    wire N__65215;
    wire N__65212;
    wire N__65209;
    wire N__65206;
    wire N__65203;
    wire N__65202;
    wire N__65201;
    wire N__65198;
    wire N__65195;
    wire N__65194;
    wire N__65193;
    wire N__65192;
    wire N__65189;
    wire N__65188;
    wire N__65185;
    wire N__65182;
    wire N__65179;
    wire N__65178;
    wire N__65175;
    wire N__65172;
    wire N__65171;
    wire N__65170;
    wire N__65169;
    wire N__65166;
    wire N__65163;
    wire N__65156;
    wire N__65153;
    wire N__65152;
    wire N__65149;
    wire N__65146;
    wire N__65143;
    wire N__65140;
    wire N__65139;
    wire N__65136;
    wire N__65135;
    wire N__65132;
    wire N__65129;
    wire N__65126;
    wire N__65123;
    wire N__65120;
    wire N__65119;
    wire N__65118;
    wire N__65109;
    wire N__65106;
    wire N__65103;
    wire N__65100;
    wire N__65095;
    wire N__65090;
    wire N__65087;
    wire N__65082;
    wire N__65077;
    wire N__65072;
    wire N__65065;
    wire N__65062;
    wire N__65061;
    wire N__65058;
    wire N__65055;
    wire N__65050;
    wire N__65047;
    wire N__65038;
    wire N__65035;
    wire N__65032;
    wire N__65029;
    wire N__65026;
    wire N__65023;
    wire N__65020;
    wire N__65017;
    wire N__65016;
    wire N__65015;
    wire N__65014;
    wire N__65013;
    wire N__65012;
    wire N__65011;
    wire N__65010;
    wire N__65009;
    wire N__65008;
    wire N__65007;
    wire N__65006;
    wire N__65005;
    wire N__65004;
    wire N__65001;
    wire N__64998;
    wire N__64995;
    wire N__64992;
    wire N__64989;
    wire N__64986;
    wire N__64983;
    wire N__64980;
    wire N__64977;
    wire N__64974;
    wire N__64971;
    wire N__64968;
    wire N__64965;
    wire N__64964;
    wire N__64961;
    wire N__64960;
    wire N__64957;
    wire N__64956;
    wire N__64955;
    wire N__64948;
    wire N__64947;
    wire N__64940;
    wire N__64933;
    wire N__64922;
    wire N__64921;
    wire N__64918;
    wire N__64915;
    wire N__64914;
    wire N__64911;
    wire N__64910;
    wire N__64907;
    wire N__64904;
    wire N__64901;
    wire N__64900;
    wire N__64899;
    wire N__64892;
    wire N__64889;
    wire N__64888;
    wire N__64887;
    wire N__64884;
    wire N__64881;
    wire N__64878;
    wire N__64875;
    wire N__64872;
    wire N__64869;
    wire N__64864;
    wire N__64863;
    wire N__64862;
    wire N__64859;
    wire N__64856;
    wire N__64851;
    wire N__64848;
    wire N__64845;
    wire N__64844;
    wire N__64837;
    wire N__64832;
    wire N__64829;
    wire N__64826;
    wire N__64823;
    wire N__64820;
    wire N__64817;
    wire N__64810;
    wire N__64807;
    wire N__64804;
    wire N__64801;
    wire N__64798;
    wire N__64787;
    wire N__64782;
    wire N__64779;
    wire N__64776;
    wire N__64771;
    wire N__64766;
    wire N__64759;
    wire N__64758;
    wire N__64755;
    wire N__64754;
    wire N__64753;
    wire N__64750;
    wire N__64749;
    wire N__64748;
    wire N__64747;
    wire N__64744;
    wire N__64741;
    wire N__64738;
    wire N__64735;
    wire N__64734;
    wire N__64731;
    wire N__64728;
    wire N__64727;
    wire N__64726;
    wire N__64723;
    wire N__64720;
    wire N__64717;
    wire N__64714;
    wire N__64713;
    wire N__64712;
    wire N__64709;
    wire N__64706;
    wire N__64703;
    wire N__64700;
    wire N__64697;
    wire N__64694;
    wire N__64693;
    wire N__64690;
    wire N__64683;
    wire N__64680;
    wire N__64677;
    wire N__64674;
    wire N__64671;
    wire N__64666;
    wire N__64663;
    wire N__64660;
    wire N__64657;
    wire N__64648;
    wire N__64647;
    wire N__64646;
    wire N__64645;
    wire N__64644;
    wire N__64643;
    wire N__64642;
    wire N__64641;
    wire N__64640;
    wire N__64639;
    wire N__64638;
    wire N__64633;
    wire N__64632;
    wire N__64625;
    wire N__64622;
    wire N__64619;
    wire N__64616;
    wire N__64613;
    wire N__64612;
    wire N__64609;
    wire N__64606;
    wire N__64603;
    wire N__64600;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64592;
    wire N__64589;
    wire N__64588;
    wire N__64585;
    wire N__64582;
    wire N__64579;
    wire N__64576;
    wire N__64573;
    wire N__64570;
    wire N__64565;
    wire N__64556;
    wire N__64549;
    wire N__64538;
    wire N__64533;
    wire N__64528;
    wire N__64519;
    wire N__64516;
    wire N__64507;
    wire N__64504;
    wire N__64501;
    wire N__64498;
    wire N__64497;
    wire N__64496;
    wire N__64493;
    wire N__64490;
    wire N__64489;
    wire N__64488;
    wire N__64485;
    wire N__64482;
    wire N__64479;
    wire N__64478;
    wire N__64475;
    wire N__64472;
    wire N__64471;
    wire N__64470;
    wire N__64467;
    wire N__64466;
    wire N__64461;
    wire N__64458;
    wire N__64455;
    wire N__64454;
    wire N__64453;
    wire N__64452;
    wire N__64451;
    wire N__64450;
    wire N__64447;
    wire N__64444;
    wire N__64441;
    wire N__64440;
    wire N__64439;
    wire N__64438;
    wire N__64437;
    wire N__64434;
    wire N__64431;
    wire N__64426;
    wire N__64423;
    wire N__64420;
    wire N__64417;
    wire N__64414;
    wire N__64411;
    wire N__64408;
    wire N__64403;
    wire N__64400;
    wire N__64397;
    wire N__64396;
    wire N__64393;
    wire N__64392;
    wire N__64389;
    wire N__64388;
    wire N__64385;
    wire N__64384;
    wire N__64383;
    wire N__64382;
    wire N__64381;
    wire N__64378;
    wire N__64375;
    wire N__64368;
    wire N__64365;
    wire N__64362;
    wire N__64359;
    wire N__64356;
    wire N__64349;
    wire N__64336;
    wire N__64335;
    wire N__64332;
    wire N__64331;
    wire N__64328;
    wire N__64327;
    wire N__64324;
    wire N__64323;
    wire N__64320;
    wire N__64315;
    wire N__64308;
    wire N__64303;
    wire N__64298;
    wire N__64281;
    wire N__64278;
    wire N__64275;
    wire N__64268;
    wire N__64261;
    wire N__64258;
    wire N__64255;
    wire N__64252;
    wire N__64249;
    wire N__64246;
    wire N__64243;
    wire N__64242;
    wire N__64241;
    wire N__64240;
    wire N__64239;
    wire N__64238;
    wire N__64237;
    wire N__64236;
    wire N__64235;
    wire N__64234;
    wire N__64233;
    wire N__64232;
    wire N__64231;
    wire N__64230;
    wire N__64227;
    wire N__64224;
    wire N__64221;
    wire N__64220;
    wire N__64219;
    wire N__64216;
    wire N__64215;
    wire N__64212;
    wire N__64211;
    wire N__64208;
    wire N__64207;
    wire N__64204;
    wire N__64201;
    wire N__64200;
    wire N__64197;
    wire N__64196;
    wire N__64193;
    wire N__64192;
    wire N__64189;
    wire N__64186;
    wire N__64183;
    wire N__64182;
    wire N__64179;
    wire N__64178;
    wire N__64175;
    wire N__64172;
    wire N__64169;
    wire N__64166;
    wire N__64149;
    wire N__64146;
    wire N__64133;
    wire N__64132;
    wire N__64129;
    wire N__64126;
    wire N__64123;
    wire N__64120;
    wire N__64117;
    wire N__64112;
    wire N__64111;
    wire N__64108;
    wire N__64105;
    wire N__64102;
    wire N__64101;
    wire N__64098;
    wire N__64095;
    wire N__64092;
    wire N__64091;
    wire N__64090;
    wire N__64081;
    wire N__64078;
    wire N__64075;
    wire N__64072;
    wire N__64067;
    wire N__64064;
    wire N__64061;
    wire N__64054;
    wire N__64051;
    wire N__64048;
    wire N__64043;
    wire N__64038;
    wire N__64031;
    wire N__64026;
    wire N__64023;
    wire N__64020;
    wire N__64017;
    wire N__64014;
    wire N__64009;
    wire N__64000;
    wire N__63997;
    wire N__63994;
    wire N__63991;
    wire N__63988;
    wire N__63985;
    wire N__63982;
    wire N__63981;
    wire N__63980;
    wire N__63979;
    wire N__63976;
    wire N__63975;
    wire N__63974;
    wire N__63971;
    wire N__63968;
    wire N__63967;
    wire N__63964;
    wire N__63963;
    wire N__63962;
    wire N__63959;
    wire N__63956;
    wire N__63955;
    wire N__63952;
    wire N__63951;
    wire N__63950;
    wire N__63949;
    wire N__63948;
    wire N__63947;
    wire N__63946;
    wire N__63943;
    wire N__63940;
    wire N__63937;
    wire N__63936;
    wire N__63933;
    wire N__63930;
    wire N__63929;
    wire N__63926;
    wire N__63921;
    wire N__63918;
    wire N__63915;
    wire N__63912;
    wire N__63909;
    wire N__63906;
    wire N__63903;
    wire N__63900;
    wire N__63897;
    wire N__63896;
    wire N__63895;
    wire N__63894;
    wire N__63893;
    wire N__63892;
    wire N__63891;
    wire N__63890;
    wire N__63889;
    wire N__63888;
    wire N__63885;
    wire N__63882;
    wire N__63879;
    wire N__63876;
    wire N__63875;
    wire N__63872;
    wire N__63869;
    wire N__63866;
    wire N__63863;
    wire N__63862;
    wire N__63859;
    wire N__63856;
    wire N__63853;
    wire N__63846;
    wire N__63839;
    wire N__63836;
    wire N__63833;
    wire N__63830;
    wire N__63827;
    wire N__63824;
    wire N__63821;
    wire N__63818;
    wire N__63815;
    wire N__63812;
    wire N__63805;
    wire N__63802;
    wire N__63799;
    wire N__63794;
    wire N__63791;
    wire N__63788;
    wire N__63785;
    wire N__63780;
    wire N__63777;
    wire N__63772;
    wire N__63763;
    wire N__63754;
    wire N__63751;
    wire N__63746;
    wire N__63739;
    wire N__63734;
    wire N__63731;
    wire N__63720;
    wire N__63715;
    wire N__63706;
    wire N__63703;
    wire N__63700;
    wire N__63697;
    wire N__63694;
    wire N__63691;
    wire N__63688;
    wire N__63687;
    wire N__63686;
    wire N__63683;
    wire N__63682;
    wire N__63679;
    wire N__63676;
    wire N__63673;
    wire N__63670;
    wire N__63669;
    wire N__63668;
    wire N__63665;
    wire N__63662;
    wire N__63659;
    wire N__63656;
    wire N__63655;
    wire N__63652;
    wire N__63649;
    wire N__63648;
    wire N__63647;
    wire N__63644;
    wire N__63641;
    wire N__63636;
    wire N__63635;
    wire N__63634;
    wire N__63633;
    wire N__63632;
    wire N__63631;
    wire N__63630;
    wire N__63627;
    wire N__63626;
    wire N__63625;
    wire N__63624;
    wire N__63623;
    wire N__63622;
    wire N__63619;
    wire N__63616;
    wire N__63613;
    wire N__63610;
    wire N__63609;
    wire N__63608;
    wire N__63607;
    wire N__63600;
    wire N__63599;
    wire N__63596;
    wire N__63595;
    wire N__63592;
    wire N__63591;
    wire N__63588;
    wire N__63587;
    wire N__63584;
    wire N__63581;
    wire N__63578;
    wire N__63575;
    wire N__63572;
    wire N__63569;
    wire N__63566;
    wire N__63565;
    wire N__63562;
    wire N__63561;
    wire N__63558;
    wire N__63553;
    wire N__63550;
    wire N__63547;
    wire N__63544;
    wire N__63541;
    wire N__63538;
    wire N__63535;
    wire N__63518;
    wire N__63515;
    wire N__63510;
    wire N__63507;
    wire N__63504;
    wire N__63493;
    wire N__63488;
    wire N__63485;
    wire N__63482;
    wire N__63479;
    wire N__63472;
    wire N__63469;
    wire N__63464;
    wire N__63457;
    wire N__63454;
    wire N__63451;
    wire N__63448;
    wire N__63443;
    wire N__63438;
    wire N__63433;
    wire N__63424;
    wire N__63421;
    wire N__63418;
    wire N__63415;
    wire N__63412;
    wire N__63409;
    wire N__63406;
    wire N__63405;
    wire N__63402;
    wire N__63401;
    wire N__63400;
    wire N__63399;
    wire N__63396;
    wire N__63393;
    wire N__63390;
    wire N__63389;
    wire N__63386;
    wire N__63385;
    wire N__63384;
    wire N__63383;
    wire N__63382;
    wire N__63379;
    wire N__63378;
    wire N__63377;
    wire N__63374;
    wire N__63371;
    wire N__63368;
    wire N__63365;
    wire N__63362;
    wire N__63361;
    wire N__63360;
    wire N__63359;
    wire N__63358;
    wire N__63355;
    wire N__63352;
    wire N__63349;
    wire N__63346;
    wire N__63343;
    wire N__63340;
    wire N__63337;
    wire N__63336;
    wire N__63329;
    wire N__63326;
    wire N__63323;
    wire N__63320;
    wire N__63319;
    wire N__63316;
    wire N__63315;
    wire N__63312;
    wire N__63311;
    wire N__63308;
    wire N__63305;
    wire N__63302;
    wire N__63299;
    wire N__63296;
    wire N__63293;
    wire N__63290;
    wire N__63287;
    wire N__63286;
    wire N__63285;
    wire N__63284;
    wire N__63281;
    wire N__63280;
    wire N__63279;
    wire N__63274;
    wire N__63271;
    wire N__63268;
    wire N__63255;
    wire N__63252;
    wire N__63247;
    wire N__63238;
    wire N__63237;
    wire N__63234;
    wire N__63233;
    wire N__63230;
    wire N__63229;
    wire N__63226;
    wire N__63221;
    wire N__63218;
    wire N__63215;
    wire N__63210;
    wire N__63207;
    wire N__63200;
    wire N__63187;
    wire N__63184;
    wire N__63181;
    wire N__63180;
    wire N__63177;
    wire N__63174;
    wire N__63167;
    wire N__63162;
    wire N__63159;
    wire N__63148;
    wire N__63145;
    wire N__63142;
    wire N__63139;
    wire N__63136;
    wire N__63135;
    wire N__63134;
    wire N__63133;
    wire N__63132;
    wire N__63131;
    wire N__63128;
    wire N__63127;
    wire N__63124;
    wire N__63121;
    wire N__63118;
    wire N__63115;
    wire N__63114;
    wire N__63113;
    wire N__63112;
    wire N__63111;
    wire N__63110;
    wire N__63109;
    wire N__63106;
    wire N__63103;
    wire N__63100;
    wire N__63099;
    wire N__63098;
    wire N__63097;
    wire N__63096;
    wire N__63095;
    wire N__63094;
    wire N__63093;
    wire N__63084;
    wire N__63081;
    wire N__63078;
    wire N__63075;
    wire N__63072;
    wire N__63069;
    wire N__63066;
    wire N__63065;
    wire N__63062;
    wire N__63059;
    wire N__63056;
    wire N__63053;
    wire N__63052;
    wire N__63049;
    wire N__63048;
    wire N__63045;
    wire N__63044;
    wire N__63041;
    wire N__63038;
    wire N__63035;
    wire N__63032;
    wire N__63031;
    wire N__63028;
    wire N__63019;
    wire N__63016;
    wire N__63013;
    wire N__63010;
    wire N__63003;
    wire N__63000;
    wire N__62999;
    wire N__62986;
    wire N__62983;
    wire N__62978;
    wire N__62975;
    wire N__62974;
    wire N__62971;
    wire N__62968;
    wire N__62963;
    wire N__62960;
    wire N__62959;
    wire N__62954;
    wire N__62951;
    wire N__62948;
    wire N__62945;
    wire N__62942;
    wire N__62939;
    wire N__62938;
    wire N__62935;
    wire N__62930;
    wire N__62925;
    wire N__62922;
    wire N__62919;
    wire N__62916;
    wire N__62913;
    wire N__62906;
    wire N__62903;
    wire N__62900;
    wire N__62895;
    wire N__62892;
    wire N__62887;
    wire N__62882;
    wire N__62879;
    wire N__62872;
    wire N__62869;
    wire N__62866;
    wire N__62861;
    wire N__62854;
    wire N__62851;
    wire N__62848;
    wire N__62845;
    wire N__62842;
    wire N__62839;
    wire N__62836;
    wire N__62833;
    wire N__62830;
    wire N__62827;
    wire N__62824;
    wire N__62821;
    wire N__62818;
    wire N__62815;
    wire N__62812;
    wire N__62809;
    wire N__62806;
    wire N__62803;
    wire N__62800;
    wire N__62797;
    wire N__62794;
    wire N__62791;
    wire N__62788;
    wire N__62785;
    wire N__62782;
    wire N__62779;
    wire N__62776;
    wire N__62773;
    wire N__62770;
    wire N__62767;
    wire N__62764;
    wire N__62761;
    wire N__62758;
    wire N__62755;
    wire N__62752;
    wire N__62749;
    wire N__62746;
    wire N__62743;
    wire N__62740;
    wire N__62737;
    wire N__62734;
    wire N__62731;
    wire N__62728;
    wire N__62725;
    wire N__62722;
    wire N__62721;
    wire N__62718;
    wire N__62715;
    wire N__62714;
    wire N__62711;
    wire N__62708;
    wire N__62705;
    wire N__62698;
    wire N__62697;
    wire N__62694;
    wire N__62691;
    wire N__62688;
    wire N__62687;
    wire N__62684;
    wire N__62681;
    wire N__62678;
    wire N__62671;
    wire N__62668;
    wire N__62667;
    wire N__62664;
    wire N__62661;
    wire N__62660;
    wire N__62655;
    wire N__62652;
    wire N__62647;
    wire N__62644;
    wire N__62641;
    wire N__62638;
    wire N__62635;
    wire N__62632;
    wire N__62629;
    wire N__62626;
    wire N__62623;
    wire N__62620;
    wire N__62617;
    wire N__62614;
    wire N__62611;
    wire N__62608;
    wire N__62605;
    wire N__62602;
    wire N__62599;
    wire N__62596;
    wire N__62593;
    wire N__62590;
    wire N__62587;
    wire N__62584;
    wire N__62581;
    wire N__62578;
    wire N__62575;
    wire N__62572;
    wire N__62569;
    wire N__62566;
    wire N__62565;
    wire N__62564;
    wire N__62561;
    wire N__62556;
    wire N__62551;
    wire N__62548;
    wire N__62547;
    wire N__62544;
    wire N__62541;
    wire N__62536;
    wire N__62535;
    wire N__62534;
    wire N__62531;
    wire N__62528;
    wire N__62525;
    wire N__62518;
    wire N__62517;
    wire N__62516;
    wire N__62513;
    wire N__62510;
    wire N__62507;
    wire N__62504;
    wire N__62501;
    wire N__62494;
    wire N__62491;
    wire N__62490;
    wire N__62487;
    wire N__62484;
    wire N__62483;
    wire N__62480;
    wire N__62477;
    wire N__62474;
    wire N__62467;
    wire N__62464;
    wire N__62461;
    wire N__62460;
    wire N__62459;
    wire N__62456;
    wire N__62453;
    wire N__62450;
    wire N__62443;
    wire N__62440;
    wire N__62437;
    wire N__62436;
    wire N__62435;
    wire N__62432;
    wire N__62429;
    wire N__62426;
    wire N__62419;
    wire N__62416;
    wire N__62415;
    wire N__62412;
    wire N__62411;
    wire N__62408;
    wire N__62405;
    wire N__62402;
    wire N__62395;
    wire N__62392;
    wire N__62389;
    wire N__62388;
    wire N__62387;
    wire N__62384;
    wire N__62381;
    wire N__62378;
    wire N__62371;
    wire N__62368;
    wire N__62367;
    wire N__62366;
    wire N__62363;
    wire N__62360;
    wire N__62357;
    wire N__62350;
    wire N__62347;
    wire N__62344;
    wire N__62341;
    wire N__62340;
    wire N__62339;
    wire N__62336;
    wire N__62333;
    wire N__62330;
    wire N__62323;
    wire N__62320;
    wire N__62317;
    wire N__62314;
    wire N__62311;
    wire N__62308;
    wire N__62307;
    wire N__62304;
    wire N__62301;
    wire N__62300;
    wire N__62297;
    wire N__62294;
    wire N__62291;
    wire N__62284;
    wire N__62283;
    wire N__62280;
    wire N__62279;
    wire N__62276;
    wire N__62273;
    wire N__62270;
    wire N__62267;
    wire N__62264;
    wire N__62261;
    wire N__62254;
    wire N__62251;
    wire N__62250;
    wire N__62247;
    wire N__62244;
    wire N__62243;
    wire N__62238;
    wire N__62235;
    wire N__62230;
    wire N__62227;
    wire N__62226;
    wire N__62223;
    wire N__62220;
    wire N__62215;
    wire N__62214;
    wire N__62211;
    wire N__62208;
    wire N__62203;
    wire N__62202;
    wire N__62199;
    wire N__62196;
    wire N__62191;
    wire N__62190;
    wire N__62187;
    wire N__62184;
    wire N__62179;
    wire N__62176;
    wire N__62175;
    wire N__62172;
    wire N__62169;
    wire N__62166;
    wire N__62165;
    wire N__62160;
    wire N__62157;
    wire N__62152;
    wire N__62149;
    wire N__62146;
    wire N__62143;
    wire N__62142;
    wire N__62139;
    wire N__62136;
    wire N__62131;
    wire N__62130;
    wire N__62127;
    wire N__62124;
    wire N__62119;
    wire N__62118;
    wire N__62117;
    wire N__62116;
    wire N__62115;
    wire N__62114;
    wire N__62113;
    wire N__62112;
    wire N__62111;
    wire N__62110;
    wire N__62109;
    wire N__62108;
    wire N__62107;
    wire N__62106;
    wire N__62105;
    wire N__62104;
    wire N__62071;
    wire N__62068;
    wire N__62065;
    wire N__62064;
    wire N__62061;
    wire N__62060;
    wire N__62057;
    wire N__62054;
    wire N__62051;
    wire N__62048;
    wire N__62045;
    wire N__62040;
    wire N__62035;
    wire N__62032;
    wire N__62029;
    wire N__62028;
    wire N__62027;
    wire N__62026;
    wire N__62025;
    wire N__62024;
    wire N__62023;
    wire N__62022;
    wire N__62021;
    wire N__62020;
    wire N__62019;
    wire N__62018;
    wire N__62017;
    wire N__62016;
    wire N__62015;
    wire N__61998;
    wire N__61987;
    wire N__61986;
    wire N__61985;
    wire N__61982;
    wire N__61981;
    wire N__61978;
    wire N__61977;
    wire N__61976;
    wire N__61975;
    wire N__61974;
    wire N__61973;
    wire N__61972;
    wire N__61971;
    wire N__61970;
    wire N__61969;
    wire N__61968;
    wire N__61967;
    wire N__61966;
    wire N__61961;
    wire N__61956;
    wire N__61943;
    wire N__61934;
    wire N__61923;
    wire N__61912;
    wire N__61911;
    wire N__61910;
    wire N__61909;
    wire N__61908;
    wire N__61907;
    wire N__61906;
    wire N__61905;
    wire N__61904;
    wire N__61903;
    wire N__61902;
    wire N__61901;
    wire N__61900;
    wire N__61899;
    wire N__61898;
    wire N__61897;
    wire N__61896;
    wire N__61895;
    wire N__61894;
    wire N__61893;
    wire N__61892;
    wire N__61891;
    wire N__61890;
    wire N__61889;
    wire N__61888;
    wire N__61887;
    wire N__61886;
    wire N__61885;
    wire N__61884;
    wire N__61883;
    wire N__61878;
    wire N__61869;
    wire N__61856;
    wire N__61839;
    wire N__61834;
    wire N__61827;
    wire N__61822;
    wire N__61815;
    wire N__61798;
    wire N__61795;
    wire N__61792;
    wire N__61789;
    wire N__61786;
    wire N__61783;
    wire N__61780;
    wire N__61777;
    wire N__61776;
    wire N__61775;
    wire N__61772;
    wire N__61767;
    wire N__61762;
    wire N__61759;
    wire N__61758;
    wire N__61755;
    wire N__61754;
    wire N__61751;
    wire N__61748;
    wire N__61743;
    wire N__61738;
    wire N__61735;
    wire N__61732;
    wire N__61731;
    wire N__61730;
    wire N__61727;
    wire N__61722;
    wire N__61717;
    wire N__61716;
    wire N__61713;
    wire N__61712;
    wire N__61709;
    wire N__61706;
    wire N__61703;
    wire N__61700;
    wire N__61697;
    wire N__61692;
    wire N__61687;
    wire N__61686;
    wire N__61685;
    wire N__61680;
    wire N__61677;
    wire N__61674;
    wire N__61671;
    wire N__61668;
    wire N__61665;
    wire N__61660;
    wire N__61657;
    wire N__61656;
    wire N__61655;
    wire N__61650;
    wire N__61647;
    wire N__61642;
    wire N__61639;
    wire N__61636;
    wire N__61633;
    wire N__61630;
    wire N__61629;
    wire N__61626;
    wire N__61623;
    wire N__61622;
    wire N__61619;
    wire N__61616;
    wire N__61613;
    wire N__61610;
    wire N__61605;
    wire N__61600;
    wire N__61597;
    wire N__61596;
    wire N__61593;
    wire N__61592;
    wire N__61589;
    wire N__61586;
    wire N__61583;
    wire N__61580;
    wire N__61575;
    wire N__61570;
    wire N__61567;
    wire N__61564;
    wire N__61561;
    wire N__61558;
    wire N__61555;
    wire N__61552;
    wire N__61551;
    wire N__61550;
    wire N__61547;
    wire N__61542;
    wire N__61539;
    wire N__61536;
    wire N__61531;
    wire N__61530;
    wire N__61529;
    wire N__61526;
    wire N__61521;
    wire N__61516;
    wire N__61513;
    wire N__61510;
    wire N__61507;
    wire N__61504;
    wire N__61501;
    wire N__61498;
    wire N__61495;
    wire N__61492;
    wire N__61489;
    wire N__61486;
    wire N__61483;
    wire N__61480;
    wire N__61479;
    wire N__61478;
    wire N__61477;
    wire N__61476;
    wire N__61475;
    wire N__61472;
    wire N__61471;
    wire N__61470;
    wire N__61469;
    wire N__61466;
    wire N__61463;
    wire N__61462;
    wire N__61461;
    wire N__61460;
    wire N__61459;
    wire N__61458;
    wire N__61455;
    wire N__61454;
    wire N__61451;
    wire N__61450;
    wire N__61449;
    wire N__61446;
    wire N__61437;
    wire N__61426;
    wire N__61421;
    wire N__61418;
    wire N__61415;
    wire N__61412;
    wire N__61405;
    wire N__61390;
    wire N__61389;
    wire N__61388;
    wire N__61387;
    wire N__61386;
    wire N__61383;
    wire N__61382;
    wire N__61381;
    wire N__61380;
    wire N__61379;
    wire N__61378;
    wire N__61377;
    wire N__61376;
    wire N__61375;
    wire N__61374;
    wire N__61373;
    wire N__61372;
    wire N__61371;
    wire N__61368;
    wire N__61365;
    wire N__61356;
    wire N__61347;
    wire N__61336;
    wire N__61331;
    wire N__61318;
    wire N__61315;
    wire N__61312;
    wire N__61309;
    wire N__61306;
    wire N__61303;
    wire N__61300;
    wire N__61297;
    wire N__61294;
    wire N__61291;
    wire N__61288;
    wire N__61285;
    wire N__61282;
    wire N__61279;
    wire N__61276;
    wire N__61273;
    wire N__61270;
    wire N__61267;
    wire N__61264;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61252;
    wire N__61249;
    wire N__61246;
    wire N__61243;
    wire N__61240;
    wire N__61237;
    wire N__61236;
    wire N__61233;
    wire N__61230;
    wire N__61227;
    wire N__61224;
    wire N__61221;
    wire N__61218;
    wire N__61213;
    wire N__61210;
    wire N__61207;
    wire N__61204;
    wire N__61201;
    wire N__61200;
    wire N__61197;
    wire N__61194;
    wire N__61189;
    wire N__61186;
    wire N__61183;
    wire N__61180;
    wire N__61177;
    wire N__61174;
    wire N__61171;
    wire N__61168;
    wire N__61165;
    wire N__61162;
    wire N__61159;
    wire N__61156;
    wire N__61153;
    wire N__61150;
    wire N__61147;
    wire N__61144;
    wire N__61141;
    wire N__61138;
    wire N__61135;
    wire N__61132;
    wire N__61129;
    wire N__61126;
    wire N__61123;
    wire N__61120;
    wire N__61117;
    wire N__61114;
    wire N__61111;
    wire N__61108;
    wire N__61105;
    wire N__61102;
    wire N__61099;
    wire N__61096;
    wire N__61093;
    wire N__61090;
    wire N__61087;
    wire N__61084;
    wire N__61081;
    wire N__61078;
    wire N__61075;
    wire N__61072;
    wire N__61069;
    wire N__61066;
    wire N__61063;
    wire N__61060;
    wire N__61057;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61042;
    wire N__61039;
    wire N__61036;
    wire N__61033;
    wire N__61030;
    wire N__61027;
    wire N__61024;
    wire N__61021;
    wire N__61018;
    wire N__61015;
    wire N__61012;
    wire N__61009;
    wire N__61006;
    wire N__61003;
    wire N__61000;
    wire N__60997;
    wire N__60994;
    wire N__60991;
    wire N__60988;
    wire N__60985;
    wire N__60982;
    wire N__60979;
    wire N__60976;
    wire N__60973;
    wire N__60970;
    wire N__60967;
    wire N__60966;
    wire N__60963;
    wire N__60960;
    wire N__60959;
    wire N__60958;
    wire N__60957;
    wire N__60956;
    wire N__60955;
    wire N__60954;
    wire N__60953;
    wire N__60952;
    wire N__60951;
    wire N__60946;
    wire N__60943;
    wire N__60940;
    wire N__60939;
    wire N__60938;
    wire N__60935;
    wire N__60934;
    wire N__60931;
    wire N__60930;
    wire N__60927;
    wire N__60926;
    wire N__60923;
    wire N__60922;
    wire N__60919;
    wire N__60918;
    wire N__60915;
    wire N__60914;
    wire N__60911;
    wire N__60904;
    wire N__60903;
    wire N__60902;
    wire N__60899;
    wire N__60886;
    wire N__60869;
    wire N__60866;
    wire N__60863;
    wire N__60862;
    wire N__60859;
    wire N__60858;
    wire N__60857;
    wire N__60856;
    wire N__60853;
    wire N__60848;
    wire N__60843;
    wire N__60840;
    wire N__60839;
    wire N__60836;
    wire N__60833;
    wire N__60830;
    wire N__60829;
    wire N__60828;
    wire N__60825;
    wire N__60822;
    wire N__60817;
    wire N__60814;
    wire N__60811;
    wire N__60806;
    wire N__60803;
    wire N__60800;
    wire N__60797;
    wire N__60796;
    wire N__60793;
    wire N__60786;
    wire N__60783;
    wire N__60774;
    wire N__60771;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60757;
    wire N__60748;
    wire N__60745;
    wire N__60742;
    wire N__60739;
    wire N__60736;
    wire N__60733;
    wire N__60730;
    wire N__60727;
    wire N__60724;
    wire N__60721;
    wire N__60718;
    wire N__60715;
    wire N__60712;
    wire N__60709;
    wire N__60706;
    wire N__60703;
    wire N__60700;
    wire N__60697;
    wire N__60694;
    wire N__60691;
    wire N__60688;
    wire N__60685;
    wire N__60682;
    wire N__60679;
    wire N__60676;
    wire N__60673;
    wire N__60670;
    wire N__60667;
    wire N__60664;
    wire N__60661;
    wire N__60658;
    wire N__60655;
    wire N__60652;
    wire N__60649;
    wire N__60646;
    wire N__60643;
    wire N__60640;
    wire N__60637;
    wire N__60634;
    wire N__60631;
    wire N__60628;
    wire N__60625;
    wire N__60622;
    wire N__60619;
    wire N__60616;
    wire N__60613;
    wire N__60610;
    wire N__60607;
    wire N__60604;
    wire N__60601;
    wire N__60598;
    wire N__60595;
    wire N__60592;
    wire N__60589;
    wire N__60586;
    wire N__60583;
    wire N__60580;
    wire N__60577;
    wire N__60574;
    wire N__60571;
    wire N__60568;
    wire N__60565;
    wire N__60562;
    wire N__60559;
    wire N__60556;
    wire N__60553;
    wire N__60550;
    wire N__60547;
    wire N__60544;
    wire N__60541;
    wire N__60538;
    wire N__60535;
    wire N__60532;
    wire N__60529;
    wire N__60526;
    wire N__60523;
    wire N__60520;
    wire N__60517;
    wire N__60514;
    wire N__60511;
    wire N__60508;
    wire N__60505;
    wire N__60502;
    wire N__60499;
    wire N__60496;
    wire N__60493;
    wire N__60490;
    wire N__60487;
    wire N__60484;
    wire N__60481;
    wire N__60478;
    wire N__60475;
    wire N__60472;
    wire N__60469;
    wire N__60466;
    wire N__60463;
    wire N__60460;
    wire N__60457;
    wire N__60454;
    wire N__60451;
    wire N__60448;
    wire N__60447;
    wire N__60444;
    wire N__60443;
    wire N__60442;
    wire N__60441;
    wire N__60438;
    wire N__60433;
    wire N__60426;
    wire N__60421;
    wire N__60418;
    wire N__60415;
    wire N__60412;
    wire N__60411;
    wire N__60408;
    wire N__60405;
    wire N__60402;
    wire N__60399;
    wire N__60398;
    wire N__60395;
    wire N__60392;
    wire N__60389;
    wire N__60382;
    wire N__60381;
    wire N__60376;
    wire N__60375;
    wire N__60372;
    wire N__60369;
    wire N__60366;
    wire N__60363;
    wire N__60358;
    wire N__60355;
    wire N__60354;
    wire N__60351;
    wire N__60348;
    wire N__60345;
    wire N__60342;
    wire N__60341;
    wire N__60336;
    wire N__60333;
    wire N__60328;
    wire N__60327;
    wire N__60322;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60310;
    wire N__60309;
    wire N__60304;
    wire N__60303;
    wire N__60300;
    wire N__60297;
    wire N__60292;
    wire N__60289;
    wire N__60286;
    wire N__60285;
    wire N__60282;
    wire N__60279;
    wire N__60274;
    wire N__60271;
    wire N__60270;
    wire N__60267;
    wire N__60264;
    wire N__60259;
    wire N__60258;
    wire N__60255;
    wire N__60252;
    wire N__60251;
    wire N__60248;
    wire N__60245;
    wire N__60242;
    wire N__60239;
    wire N__60234;
    wire N__60229;
    wire N__60226;
    wire N__60223;
    wire N__60222;
    wire N__60219;
    wire N__60216;
    wire N__60215;
    wire N__60212;
    wire N__60209;
    wire N__60206;
    wire N__60199;
    wire N__60196;
    wire N__60193;
    wire N__60190;
    wire N__60189;
    wire N__60186;
    wire N__60183;
    wire N__60178;
    wire N__60175;
    wire N__60174;
    wire N__60171;
    wire N__60168;
    wire N__60163;
    wire N__60160;
    wire N__60157;
    wire N__60154;
    wire N__60151;
    wire N__60148;
    wire N__60147;
    wire N__60144;
    wire N__60141;
    wire N__60140;
    wire N__60137;
    wire N__60132;
    wire N__60127;
    wire N__60124;
    wire N__60123;
    wire N__60120;
    wire N__60117;
    wire N__60112;
    wire N__60111;
    wire N__60110;
    wire N__60107;
    wire N__60102;
    wire N__60097;
    wire N__60094;
    wire N__60093;
    wire N__60092;
    wire N__60089;
    wire N__60084;
    wire N__60079;
    wire N__60076;
    wire N__60073;
    wire N__60070;
    wire N__60069;
    wire N__60068;
    wire N__60065;
    wire N__60060;
    wire N__60055;
    wire N__60052;
    wire N__60049;
    wire N__60046;
    wire N__60043;
    wire N__60040;
    wire N__60037;
    wire N__60034;
    wire N__60031;
    wire N__60028;
    wire N__60025;
    wire N__60022;
    wire N__60019;
    wire N__60016;
    wire N__60013;
    wire N__60010;
    wire N__60007;
    wire N__60006;
    wire N__60005;
    wire N__59998;
    wire N__59995;
    wire N__59992;
    wire N__59989;
    wire N__59986;
    wire N__59983;
    wire N__59980;
    wire N__59977;
    wire N__59974;
    wire N__59973;
    wire N__59972;
    wire N__59965;
    wire N__59962;
    wire N__59959;
    wire N__59956;
    wire N__59953;
    wire N__59950;
    wire N__59947;
    wire N__59944;
    wire N__59941;
    wire N__59938;
    wire N__59935;
    wire N__59932;
    wire N__59929;
    wire N__59926;
    wire N__59923;
    wire N__59920;
    wire N__59917;
    wire N__59914;
    wire N__59911;
    wire N__59908;
    wire N__59905;
    wire N__59902;
    wire N__59899;
    wire N__59896;
    wire N__59893;
    wire N__59890;
    wire N__59887;
    wire N__59884;
    wire N__59881;
    wire N__59878;
    wire N__59875;
    wire N__59872;
    wire N__59869;
    wire N__59866;
    wire N__59863;
    wire N__59860;
    wire N__59857;
    wire N__59854;
    wire N__59851;
    wire N__59848;
    wire N__59845;
    wire N__59842;
    wire N__59839;
    wire N__59836;
    wire N__59833;
    wire N__59830;
    wire N__59827;
    wire N__59824;
    wire N__59821;
    wire N__59818;
    wire N__59815;
    wire N__59812;
    wire N__59809;
    wire N__59806;
    wire N__59803;
    wire N__59800;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59787;
    wire N__59786;
    wire N__59783;
    wire N__59778;
    wire N__59773;
    wire N__59770;
    wire N__59767;
    wire N__59764;
    wire N__59761;
    wire N__59758;
    wire N__59755;
    wire N__59752;
    wire N__59749;
    wire N__59746;
    wire N__59743;
    wire N__59740;
    wire N__59737;
    wire N__59734;
    wire N__59731;
    wire N__59728;
    wire N__59725;
    wire N__59722;
    wire N__59719;
    wire N__59716;
    wire N__59713;
    wire N__59710;
    wire N__59707;
    wire N__59704;
    wire N__59701;
    wire N__59698;
    wire N__59695;
    wire N__59692;
    wire N__59689;
    wire N__59686;
    wire N__59683;
    wire N__59680;
    wire N__59677;
    wire N__59674;
    wire N__59671;
    wire N__59668;
    wire N__59665;
    wire N__59662;
    wire N__59659;
    wire N__59656;
    wire N__59653;
    wire N__59650;
    wire N__59647;
    wire N__59644;
    wire N__59641;
    wire N__59638;
    wire N__59635;
    wire N__59632;
    wire N__59629;
    wire N__59626;
    wire N__59623;
    wire N__59620;
    wire N__59617;
    wire N__59614;
    wire N__59611;
    wire N__59608;
    wire N__59605;
    wire N__59602;
    wire N__59599;
    wire N__59596;
    wire N__59593;
    wire N__59590;
    wire N__59587;
    wire N__59584;
    wire N__59581;
    wire N__59578;
    wire N__59575;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59560;
    wire N__59557;
    wire N__59554;
    wire N__59551;
    wire N__59548;
    wire N__59545;
    wire N__59542;
    wire N__59539;
    wire N__59536;
    wire N__59533;
    wire N__59530;
    wire N__59527;
    wire N__59524;
    wire N__59521;
    wire N__59518;
    wire N__59515;
    wire N__59512;
    wire N__59509;
    wire N__59506;
    wire N__59503;
    wire N__59500;
    wire N__59497;
    wire N__59494;
    wire N__59491;
    wire N__59488;
    wire N__59485;
    wire N__59482;
    wire N__59481;
    wire N__59476;
    wire N__59473;
    wire N__59470;
    wire N__59467;
    wire N__59466;
    wire N__59465;
    wire N__59462;
    wire N__59459;
    wire N__59456;
    wire N__59449;
    wire N__59446;
    wire N__59443;
    wire N__59442;
    wire N__59441;
    wire N__59440;
    wire N__59437;
    wire N__59434;
    wire N__59433;
    wire N__59430;
    wire N__59429;
    wire N__59428;
    wire N__59427;
    wire N__59426;
    wire N__59425;
    wire N__59424;
    wire N__59423;
    wire N__59420;
    wire N__59419;
    wire N__59418;
    wire N__59417;
    wire N__59416;
    wire N__59415;
    wire N__59412;
    wire N__59409;
    wire N__59402;
    wire N__59391;
    wire N__59388;
    wire N__59381;
    wire N__59374;
    wire N__59359;
    wire N__59358;
    wire N__59355;
    wire N__59352;
    wire N__59351;
    wire N__59350;
    wire N__59345;
    wire N__59342;
    wire N__59339;
    wire N__59336;
    wire N__59331;
    wire N__59326;
    wire N__59325;
    wire N__59322;
    wire N__59319;
    wire N__59316;
    wire N__59315;
    wire N__59312;
    wire N__59309;
    wire N__59308;
    wire N__59307;
    wire N__59306;
    wire N__59305;
    wire N__59304;
    wire N__59301;
    wire N__59300;
    wire N__59299;
    wire N__59298;
    wire N__59297;
    wire N__59296;
    wire N__59295;
    wire N__59294;
    wire N__59293;
    wire N__59292;
    wire N__59287;
    wire N__59280;
    wire N__59269;
    wire N__59266;
    wire N__59259;
    wire N__59252;
    wire N__59239;
    wire N__59236;
    wire N__59233;
    wire N__59230;
    wire N__59227;
    wire N__59224;
    wire N__59221;
    wire N__59218;
    wire N__59215;
    wire N__59212;
    wire N__59209;
    wire N__59206;
    wire N__59203;
    wire N__59200;
    wire N__59197;
    wire N__59196;
    wire N__59191;
    wire N__59188;
    wire N__59185;
    wire N__59182;
    wire N__59181;
    wire N__59180;
    wire N__59177;
    wire N__59174;
    wire N__59171;
    wire N__59164;
    wire N__59161;
    wire N__59158;
    wire N__59155;
    wire N__59152;
    wire N__59151;
    wire N__59150;
    wire N__59147;
    wire N__59144;
    wire N__59141;
    wire N__59134;
    wire N__59131;
    wire N__59128;
    wire N__59125;
    wire N__59122;
    wire N__59119;
    wire N__59116;
    wire N__59113;
    wire N__59110;
    wire N__59107;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59092;
    wire N__59089;
    wire N__59086;
    wire N__59083;
    wire N__59080;
    wire N__59077;
    wire N__59074;
    wire N__59071;
    wire N__59068;
    wire N__59065;
    wire N__59062;
    wire N__59059;
    wire N__59056;
    wire N__59053;
    wire N__59050;
    wire N__59047;
    wire N__59044;
    wire N__59041;
    wire N__59038;
    wire N__59035;
    wire N__59032;
    wire N__59029;
    wire N__59026;
    wire N__59023;
    wire N__59020;
    wire N__59017;
    wire N__59014;
    wire N__59011;
    wire N__59008;
    wire N__59005;
    wire N__59002;
    wire N__58999;
    wire N__58996;
    wire N__58993;
    wire N__58990;
    wire N__58987;
    wire N__58984;
    wire N__58983;
    wire N__58980;
    wire N__58977;
    wire N__58972;
    wire N__58969;
    wire N__58966;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58951;
    wire N__58948;
    wire N__58945;
    wire N__58942;
    wire N__58939;
    wire N__58936;
    wire N__58933;
    wire N__58930;
    wire N__58927;
    wire N__58924;
    wire N__58921;
    wire N__58918;
    wire N__58915;
    wire N__58912;
    wire N__58911;
    wire N__58910;
    wire N__58909;
    wire N__58908;
    wire N__58907;
    wire N__58906;
    wire N__58905;
    wire N__58904;
    wire N__58903;
    wire N__58902;
    wire N__58901;
    wire N__58900;
    wire N__58899;
    wire N__58896;
    wire N__58895;
    wire N__58892;
    wire N__58891;
    wire N__58888;
    wire N__58887;
    wire N__58884;
    wire N__58881;
    wire N__58878;
    wire N__58875;
    wire N__58874;
    wire N__58871;
    wire N__58870;
    wire N__58867;
    wire N__58866;
    wire N__58865;
    wire N__58864;
    wire N__58861;
    wire N__58860;
    wire N__58857;
    wire N__58856;
    wire N__58853;
    wire N__58852;
    wire N__58849;
    wire N__58846;
    wire N__58845;
    wire N__58842;
    wire N__58829;
    wire N__58826;
    wire N__58823;
    wire N__58820;
    wire N__58817;
    wire N__58814;
    wire N__58811;
    wire N__58810;
    wire N__58807;
    wire N__58804;
    wire N__58801;
    wire N__58784;
    wire N__58781;
    wire N__58780;
    wire N__58777;
    wire N__58772;
    wire N__58765;
    wire N__58762;
    wire N__58759;
    wire N__58756;
    wire N__58755;
    wire N__58752;
    wire N__58747;
    wire N__58740;
    wire N__58737;
    wire N__58734;
    wire N__58731;
    wire N__58722;
    wire N__58719;
    wire N__58716;
    wire N__58707;
    wire N__58698;
    wire N__58695;
    wire N__58692;
    wire N__58687;
    wire N__58684;
    wire N__58681;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58651;
    wire N__58648;
    wire N__58645;
    wire N__58642;
    wire N__58639;
    wire N__58636;
    wire N__58633;
    wire N__58630;
    wire N__58627;
    wire N__58624;
    wire N__58621;
    wire N__58618;
    wire N__58615;
    wire N__58612;
    wire N__58609;
    wire N__58606;
    wire N__58603;
    wire N__58600;
    wire N__58597;
    wire N__58594;
    wire N__58591;
    wire N__58588;
    wire N__58585;
    wire N__58582;
    wire N__58579;
    wire N__58576;
    wire N__58573;
    wire N__58570;
    wire N__58567;
    wire N__58564;
    wire N__58561;
    wire N__58558;
    wire N__58555;
    wire N__58552;
    wire N__58549;
    wire N__58546;
    wire N__58543;
    wire N__58540;
    wire N__58537;
    wire N__58534;
    wire N__58531;
    wire N__58528;
    wire N__58525;
    wire N__58522;
    wire N__58519;
    wire N__58516;
    wire N__58513;
    wire N__58512;
    wire N__58509;
    wire N__58506;
    wire N__58503;
    wire N__58500;
    wire N__58497;
    wire N__58494;
    wire N__58489;
    wire N__58488;
    wire N__58487;
    wire N__58482;
    wire N__58479;
    wire N__58476;
    wire N__58473;
    wire N__58470;
    wire N__58467;
    wire N__58464;
    wire N__58459;
    wire N__58456;
    wire N__58453;
    wire N__58452;
    wire N__58451;
    wire N__58450;
    wire N__58447;
    wire N__58446;
    wire N__58443;
    wire N__58442;
    wire N__58439;
    wire N__58438;
    wire N__58435;
    wire N__58434;
    wire N__58433;
    wire N__58430;
    wire N__58415;
    wire N__58412;
    wire N__58405;
    wire N__58404;
    wire N__58403;
    wire N__58400;
    wire N__58399;
    wire N__58396;
    wire N__58395;
    wire N__58392;
    wire N__58381;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58369;
    wire N__58368;
    wire N__58367;
    wire N__58364;
    wire N__58361;
    wire N__58358;
    wire N__58353;
    wire N__58350;
    wire N__58347;
    wire N__58344;
    wire N__58339;
    wire N__58336;
    wire N__58333;
    wire N__58330;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58309;
    wire N__58306;
    wire N__58303;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58279;
    wire N__58278;
    wire N__58275;
    wire N__58272;
    wire N__58269;
    wire N__58266;
    wire N__58263;
    wire N__58260;
    wire N__58255;
    wire N__58252;
    wire N__58249;
    wire N__58246;
    wire N__58243;
    wire N__58240;
    wire N__58239;
    wire N__58238;
    wire N__58235;
    wire N__58232;
    wire N__58229;
    wire N__58222;
    wire N__58219;
    wire N__58216;
    wire N__58213;
    wire N__58212;
    wire N__58209;
    wire N__58206;
    wire N__58203;
    wire N__58200;
    wire N__58197;
    wire N__58194;
    wire N__58191;
    wire N__58186;
    wire N__58183;
    wire N__58180;
    wire N__58177;
    wire N__58174;
    wire N__58171;
    wire N__58170;
    wire N__58169;
    wire N__58164;
    wire N__58161;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58147;
    wire N__58144;
    wire N__58141;
    wire N__58140;
    wire N__58137;
    wire N__58134;
    wire N__58129;
    wire N__58126;
    wire N__58123;
    wire N__58120;
    wire N__58117;
    wire N__58114;
    wire N__58111;
    wire N__58110;
    wire N__58109;
    wire N__58106;
    wire N__58101;
    wire N__58098;
    wire N__58095;
    wire N__58092;
    wire N__58089;
    wire N__58084;
    wire N__58081;
    wire N__58080;
    wire N__58077;
    wire N__58074;
    wire N__58071;
    wire N__58068;
    wire N__58065;
    wire N__58062;
    wire N__58057;
    wire N__58054;
    wire N__58051;
    wire N__58048;
    wire N__58045;
    wire N__58042;
    wire N__58041;
    wire N__58040;
    wire N__58035;
    wire N__58032;
    wire N__58029;
    wire N__58026;
    wire N__58021;
    wire N__58018;
    wire N__58015;
    wire N__58012;
    wire N__58011;
    wire N__58008;
    wire N__58005;
    wire N__58002;
    wire N__57999;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57987;
    wire N__57986;
    wire N__57981;
    wire N__57978;
    wire N__57973;
    wire N__57970;
    wire N__57967;
    wire N__57964;
    wire N__57963;
    wire N__57960;
    wire N__57957;
    wire N__57954;
    wire N__57951;
    wire N__57948;
    wire N__57945;
    wire N__57940;
    wire N__57939;
    wire N__57938;
    wire N__57935;
    wire N__57932;
    wire N__57929;
    wire N__57922;
    wire N__57919;
    wire N__57916;
    wire N__57913;
    wire N__57910;
    wire N__57909;
    wire N__57906;
    wire N__57903;
    wire N__57898;
    wire N__57895;
    wire N__57892;
    wire N__57889;
    wire N__57888;
    wire N__57887;
    wire N__57884;
    wire N__57879;
    wire N__57876;
    wire N__57871;
    wire N__57868;
    wire N__57865;
    wire N__57862;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57841;
    wire N__57838;
    wire N__57835;
    wire N__57832;
    wire N__57829;
    wire N__57826;
    wire N__57823;
    wire N__57820;
    wire N__57817;
    wire N__57814;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57802;
    wire N__57799;
    wire N__57796;
    wire N__57793;
    wire N__57790;
    wire N__57787;
    wire N__57786;
    wire N__57785;
    wire N__57782;
    wire N__57779;
    wire N__57776;
    wire N__57773;
    wire N__57770;
    wire N__57767;
    wire N__57762;
    wire N__57759;
    wire N__57754;
    wire N__57751;
    wire N__57748;
    wire N__57745;
    wire N__57744;
    wire N__57741;
    wire N__57738;
    wire N__57733;
    wire N__57730;
    wire N__57727;
    wire N__57724;
    wire N__57721;
    wire N__57718;
    wire N__57717;
    wire N__57716;
    wire N__57713;
    wire N__57710;
    wire N__57707;
    wire N__57704;
    wire N__57699;
    wire N__57696;
    wire N__57693;
    wire N__57688;
    wire N__57685;
    wire N__57684;
    wire N__57681;
    wire N__57678;
    wire N__57675;
    wire N__57672;
    wire N__57669;
    wire N__57666;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57646;
    wire N__57643;
    wire N__57640;
    wire N__57639;
    wire N__57636;
    wire N__57635;
    wire N__57632;
    wire N__57629;
    wire N__57626;
    wire N__57623;
    wire N__57620;
    wire N__57615;
    wire N__57612;
    wire N__57609;
    wire N__57604;
    wire N__57601;
    wire N__57600;
    wire N__57597;
    wire N__57594;
    wire N__57591;
    wire N__57588;
    wire N__57585;
    wire N__57582;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57565;
    wire N__57562;
    wire N__57561;
    wire N__57558;
    wire N__57555;
    wire N__57552;
    wire N__57551;
    wire N__57548;
    wire N__57545;
    wire N__57542;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57525;
    wire N__57522;
    wire N__57519;
    wire N__57514;
    wire N__57511;
    wire N__57508;
    wire N__57505;
    wire N__57502;
    wire N__57499;
    wire N__57496;
    wire N__57493;
    wire N__57492;
    wire N__57491;
    wire N__57488;
    wire N__57485;
    wire N__57482;
    wire N__57479;
    wire N__57474;
    wire N__57469;
    wire N__57466;
    wire N__57463;
    wire N__57460;
    wire N__57457;
    wire N__57456;
    wire N__57453;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57439;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57424;
    wire N__57421;
    wire N__57420;
    wire N__57419;
    wire N__57416;
    wire N__57411;
    wire N__57408;
    wire N__57405;
    wire N__57402;
    wire N__57399;
    wire N__57396;
    wire N__57393;
    wire N__57388;
    wire N__57385;
    wire N__57384;
    wire N__57381;
    wire N__57378;
    wire N__57375;
    wire N__57372;
    wire N__57367;
    wire N__57364;
    wire N__57361;
    wire N__57358;
    wire N__57355;
    wire N__57352;
    wire N__57349;
    wire N__57346;
    wire N__57343;
    wire N__57340;
    wire N__57337;
    wire N__57334;
    wire N__57333;
    wire N__57330;
    wire N__57327;
    wire N__57324;
    wire N__57321;
    wire N__57316;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57304;
    wire N__57301;
    wire N__57298;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57285;
    wire N__57280;
    wire N__57277;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57253;
    wire N__57250;
    wire N__57247;
    wire N__57244;
    wire N__57241;
    wire N__57238;
    wire N__57235;
    wire N__57232;
    wire N__57229;
    wire N__57226;
    wire N__57223;
    wire N__57220;
    wire N__57219;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57202;
    wire N__57199;
    wire N__57196;
    wire N__57195;
    wire N__57192;
    wire N__57189;
    wire N__57186;
    wire N__57183;
    wire N__57178;
    wire N__57175;
    wire N__57172;
    wire N__57169;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57157;
    wire N__57154;
    wire N__57153;
    wire N__57150;
    wire N__57147;
    wire N__57144;
    wire N__57141;
    wire N__57136;
    wire N__57133;
    wire N__57130;
    wire N__57127;
    wire N__57124;
    wire N__57121;
    wire N__57118;
    wire N__57115;
    wire N__57114;
    wire N__57111;
    wire N__57108;
    wire N__57103;
    wire N__57100;
    wire N__57097;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57070;
    wire N__57067;
    wire N__57064;
    wire N__57061;
    wire N__57058;
    wire N__57055;
    wire N__57052;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57040;
    wire N__57037;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57025;
    wire N__57022;
    wire N__57019;
    wire N__57016;
    wire N__57013;
    wire N__57010;
    wire N__57007;
    wire N__57004;
    wire N__57001;
    wire N__56998;
    wire N__56995;
    wire N__56992;
    wire N__56989;
    wire N__56986;
    wire N__56983;
    wire N__56980;
    wire N__56977;
    wire N__56974;
    wire N__56971;
    wire N__56968;
    wire N__56965;
    wire N__56962;
    wire N__56959;
    wire N__56956;
    wire N__56953;
    wire N__56950;
    wire N__56947;
    wire N__56944;
    wire N__56941;
    wire N__56938;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56926;
    wire N__56923;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56913;
    wire N__56910;
    wire N__56907;
    wire N__56904;
    wire N__56901;
    wire N__56896;
    wire N__56893;
    wire N__56890;
    wire N__56887;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56869;
    wire N__56866;
    wire N__56863;
    wire N__56860;
    wire N__56857;
    wire N__56854;
    wire N__56851;
    wire N__56848;
    wire N__56845;
    wire N__56842;
    wire N__56839;
    wire N__56836;
    wire N__56833;
    wire N__56830;
    wire N__56827;
    wire N__56824;
    wire N__56823;
    wire N__56822;
    wire N__56821;
    wire N__56820;
    wire N__56819;
    wire N__56818;
    wire N__56817;
    wire N__56814;
    wire N__56813;
    wire N__56812;
    wire N__56811;
    wire N__56810;
    wire N__56809;
    wire N__56808;
    wire N__56807;
    wire N__56806;
    wire N__56805;
    wire N__56804;
    wire N__56803;
    wire N__56802;
    wire N__56801;
    wire N__56794;
    wire N__56785;
    wire N__56784;
    wire N__56783;
    wire N__56782;
    wire N__56781;
    wire N__56780;
    wire N__56779;
    wire N__56778;
    wire N__56775;
    wire N__56766;
    wire N__56757;
    wire N__56752;
    wire N__56745;
    wire N__56740;
    wire N__56733;
    wire N__56724;
    wire N__56707;
    wire N__56704;
    wire N__56701;
    wire N__56698;
    wire N__56695;
    wire N__56692;
    wire N__56689;
    wire N__56686;
    wire N__56683;
    wire N__56680;
    wire N__56677;
    wire N__56676;
    wire N__56671;
    wire N__56668;
    wire N__56665;
    wire N__56662;
    wire N__56659;
    wire N__56656;
    wire N__56653;
    wire N__56650;
    wire N__56647;
    wire N__56644;
    wire N__56641;
    wire N__56638;
    wire N__56635;
    wire N__56632;
    wire N__56629;
    wire N__56626;
    wire N__56623;
    wire N__56620;
    wire N__56617;
    wire N__56614;
    wire N__56611;
    wire N__56608;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56596;
    wire N__56593;
    wire N__56590;
    wire N__56587;
    wire N__56584;
    wire N__56581;
    wire N__56578;
    wire N__56575;
    wire N__56572;
    wire N__56569;
    wire N__56566;
    wire N__56563;
    wire N__56560;
    wire N__56557;
    wire N__56554;
    wire N__56551;
    wire N__56548;
    wire N__56545;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56533;
    wire N__56530;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56512;
    wire N__56509;
    wire N__56506;
    wire N__56503;
    wire N__56500;
    wire N__56497;
    wire N__56494;
    wire N__56493;
    wire N__56492;
    wire N__56485;
    wire N__56484;
    wire N__56483;
    wire N__56482;
    wire N__56481;
    wire N__56480;
    wire N__56479;
    wire N__56478;
    wire N__56477;
    wire N__56476;
    wire N__56473;
    wire N__56464;
    wire N__56463;
    wire N__56462;
    wire N__56461;
    wire N__56460;
    wire N__56459;
    wire N__56458;
    wire N__56457;
    wire N__56456;
    wire N__56455;
    wire N__56454;
    wire N__56451;
    wire N__56450;
    wire N__56449;
    wire N__56448;
    wire N__56447;
    wire N__56444;
    wire N__56443;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56433;
    wire N__56428;
    wire N__56425;
    wire N__56412;
    wire N__56399;
    wire N__56390;
    wire N__56383;
    wire N__56368;
    wire N__56367;
    wire N__56366;
    wire N__56365;
    wire N__56364;
    wire N__56363;
    wire N__56362;
    wire N__56361;
    wire N__56360;
    wire N__56353;
    wire N__56352;
    wire N__56349;
    wire N__56346;
    wire N__56345;
    wire N__56344;
    wire N__56343;
    wire N__56342;
    wire N__56335;
    wire N__56332;
    wire N__56331;
    wire N__56330;
    wire N__56329;
    wire N__56326;
    wire N__56313;
    wire N__56310;
    wire N__56309;
    wire N__56308;
    wire N__56307;
    wire N__56306;
    wire N__56305;
    wire N__56304;
    wire N__56303;
    wire N__56302;
    wire N__56301;
    wire N__56300;
    wire N__56299;
    wire N__56298;
    wire N__56297;
    wire N__56294;
    wire N__56285;
    wire N__56278;
    wire N__56269;
    wire N__56260;
    wire N__56251;
    wire N__56248;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56224;
    wire N__56221;
    wire N__56218;
    wire N__56215;
    wire N__56214;
    wire N__56211;
    wire N__56208;
    wire N__56207;
    wire N__56206;
    wire N__56205;
    wire N__56204;
    wire N__56201;
    wire N__56198;
    wire N__56197;
    wire N__56194;
    wire N__56191;
    wire N__56190;
    wire N__56189;
    wire N__56186;
    wire N__56183;
    wire N__56182;
    wire N__56179;
    wire N__56176;
    wire N__56173;
    wire N__56170;
    wire N__56167;
    wire N__56164;
    wire N__56161;
    wire N__56160;
    wire N__56157;
    wire N__56154;
    wire N__56151;
    wire N__56150;
    wire N__56149;
    wire N__56148;
    wire N__56147;
    wire N__56146;
    wire N__56145;
    wire N__56142;
    wire N__56139;
    wire N__56136;
    wire N__56131;
    wire N__56128;
    wire N__56125;
    wire N__56122;
    wire N__56121;
    wire N__56116;
    wire N__56113;
    wire N__56110;
    wire N__56107;
    wire N__56106;
    wire N__56103;
    wire N__56102;
    wire N__56099;
    wire N__56098;
    wire N__56095;
    wire N__56094;
    wire N__56091;
    wire N__56090;
    wire N__56083;
    wire N__56076;
    wire N__56073;
    wire N__56070;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56042;
    wire N__56039;
    wire N__56038;
    wire N__56035;
    wire N__56030;
    wire N__56027;
    wire N__56020;
    wire N__56017;
    wire N__56014;
    wire N__56013;
    wire N__56010;
    wire N__56007;
    wire N__56004;
    wire N__55995;
    wire N__55990;
    wire N__55981;
    wire N__55978;
    wire N__55975;
    wire N__55972;
    wire N__55969;
    wire N__55966;
    wire N__55965;
    wire N__55964;
    wire N__55961;
    wire N__55960;
    wire N__55957;
    wire N__55956;
    wire N__55953;
    wire N__55950;
    wire N__55947;
    wire N__55946;
    wire N__55945;
    wire N__55944;
    wire N__55941;
    wire N__55940;
    wire N__55939;
    wire N__55936;
    wire N__55933;
    wire N__55928;
    wire N__55925;
    wire N__55922;
    wire N__55919;
    wire N__55918;
    wire N__55917;
    wire N__55916;
    wire N__55915;
    wire N__55912;
    wire N__55909;
    wire N__55906;
    wire N__55903;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55888;
    wire N__55885;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55875;
    wire N__55874;
    wire N__55873;
    wire N__55872;
    wire N__55869;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55849;
    wire N__55846;
    wire N__55843;
    wire N__55840;
    wire N__55839;
    wire N__55836;
    wire N__55835;
    wire N__55832;
    wire N__55831;
    wire N__55828;
    wire N__55827;
    wire N__55824;
    wire N__55823;
    wire N__55820;
    wire N__55813;
    wire N__55806;
    wire N__55803;
    wire N__55800;
    wire N__55797;
    wire N__55794;
    wire N__55777;
    wire N__55774;
    wire N__55769;
    wire N__55760;
    wire N__55753;
    wire N__55750;
    wire N__55747;
    wire N__55744;
    wire N__55741;
    wire N__55738;
    wire N__55737;
    wire N__55736;
    wire N__55733;
    wire N__55730;
    wire N__55729;
    wire N__55726;
    wire N__55725;
    wire N__55724;
    wire N__55723;
    wire N__55722;
    wire N__55719;
    wire N__55718;
    wire N__55717;
    wire N__55714;
    wire N__55711;
    wire N__55708;
    wire N__55705;
    wire N__55702;
    wire N__55699;
    wire N__55698;
    wire N__55697;
    wire N__55694;
    wire N__55691;
    wire N__55688;
    wire N__55685;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55673;
    wire N__55670;
    wire N__55667;
    wire N__55664;
    wire N__55663;
    wire N__55660;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55642;
    wire N__55633;
    wire N__55630;
    wire N__55627;
    wire N__55624;
    wire N__55621;
    wire N__55620;
    wire N__55619;
    wire N__55618;
    wire N__55617;
    wire N__55616;
    wire N__55615;
    wire N__55612;
    wire N__55605;
    wire N__55598;
    wire N__55595;
    wire N__55592;
    wire N__55589;
    wire N__55586;
    wire N__55583;
    wire N__55582;
    wire N__55579;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55567;
    wire N__55564;
    wire N__55557;
    wire N__55554;
    wire N__55549;
    wire N__55540;
    wire N__55537;
    wire N__55522;
    wire N__55519;
    wire N__55516;
    wire N__55513;
    wire N__55512;
    wire N__55511;
    wire N__55510;
    wire N__55509;
    wire N__55506;
    wire N__55497;
    wire N__55496;
    wire N__55495;
    wire N__55494;
    wire N__55493;
    wire N__55492;
    wire N__55491;
    wire N__55490;
    wire N__55489;
    wire N__55488;
    wire N__55487;
    wire N__55486;
    wire N__55481;
    wire N__55472;
    wire N__55465;
    wire N__55456;
    wire N__55455;
    wire N__55454;
    wire N__55453;
    wire N__55452;
    wire N__55451;
    wire N__55450;
    wire N__55449;
    wire N__55448;
    wire N__55447;
    wire N__55446;
    wire N__55445;
    wire N__55444;
    wire N__55435;
    wire N__55430;
    wire N__55423;
    wire N__55416;
    wire N__55407;
    wire N__55404;
    wire N__55395;
    wire N__55390;
    wire N__55387;
    wire N__55384;
    wire N__55381;
    wire N__55378;
    wire N__55377;
    wire N__55374;
    wire N__55371;
    wire N__55370;
    wire N__55367;
    wire N__55366;
    wire N__55365;
    wire N__55364;
    wire N__55363;
    wire N__55360;
    wire N__55357;
    wire N__55356;
    wire N__55353;
    wire N__55350;
    wire N__55349;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55341;
    wire N__55338;
    wire N__55337;
    wire N__55334;
    wire N__55331;
    wire N__55328;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55316;
    wire N__55313;
    wire N__55310;
    wire N__55307;
    wire N__55306;
    wire N__55303;
    wire N__55300;
    wire N__55297;
    wire N__55294;
    wire N__55291;
    wire N__55286;
    wire N__55283;
    wire N__55280;
    wire N__55275;
    wire N__55272;
    wire N__55269;
    wire N__55268;
    wire N__55267;
    wire N__55266;
    wire N__55263;
    wire N__55260;
    wire N__55253;
    wire N__55242;
    wire N__55239;
    wire N__55234;
    wire N__55233;
    wire N__55230;
    wire N__55229;
    wire N__55224;
    wire N__55221;
    wire N__55216;
    wire N__55213;
    wire N__55210;
    wire N__55207;
    wire N__55204;
    wire N__55189;
    wire N__55186;
    wire N__55183;
    wire N__55182;
    wire N__55181;
    wire N__55180;
    wire N__55179;
    wire N__55176;
    wire N__55173;
    wire N__55170;
    wire N__55167;
    wire N__55166;
    wire N__55163;
    wire N__55156;
    wire N__55155;
    wire N__55152;
    wire N__55151;
    wire N__55150;
    wire N__55147;
    wire N__55144;
    wire N__55141;
    wire N__55138;
    wire N__55135;
    wire N__55132;
    wire N__55129;
    wire N__55126;
    wire N__55125;
    wire N__55124;
    wire N__55123;
    wire N__55122;
    wire N__55115;
    wire N__55106;
    wire N__55103;
    wire N__55100;
    wire N__55097;
    wire N__55094;
    wire N__55093;
    wire N__55090;
    wire N__55089;
    wire N__55084;
    wire N__55077;
    wire N__55074;
    wire N__55073;
    wire N__55070;
    wire N__55067;
    wire N__55060;
    wire N__55057;
    wire N__55048;
    wire N__55045;
    wire N__55042;
    wire N__55039;
    wire N__55036;
    wire N__55033;
    wire N__55032;
    wire N__55027;
    wire N__55024;
    wire N__55021;
    wire N__55018;
    wire N__55015;
    wire N__55012;
    wire N__55009;
    wire N__55006;
    wire N__55005;
    wire N__55002;
    wire N__55001;
    wire N__54998;
    wire N__54997;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54989;
    wire N__54988;
    wire N__54987;
    wire N__54984;
    wire N__54981;
    wire N__54978;
    wire N__54973;
    wire N__54970;
    wire N__54969;
    wire N__54966;
    wire N__54963;
    wire N__54960;
    wire N__54959;
    wire N__54958;
    wire N__54955;
    wire N__54952;
    wire N__54947;
    wire N__54946;
    wire N__54945;
    wire N__54942;
    wire N__54941;
    wire N__54940;
    wire N__54935;
    wire N__54932;
    wire N__54929;
    wire N__54926;
    wire N__54923;
    wire N__54918;
    wire N__54915;
    wire N__54914;
    wire N__54911;
    wire N__54908;
    wire N__54905;
    wire N__54902;
    wire N__54895;
    wire N__54886;
    wire N__54883;
    wire N__54880;
    wire N__54873;
    wire N__54862;
    wire N__54859;
    wire N__54856;
    wire N__54853;
    wire N__54850;
    wire N__54847;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54832;
    wire N__54829;
    wire N__54826;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54814;
    wire N__54813;
    wire N__54810;
    wire N__54807;
    wire N__54806;
    wire N__54805;
    wire N__54804;
    wire N__54803;
    wire N__54802;
    wire N__54801;
    wire N__54800;
    wire N__54799;
    wire N__54798;
    wire N__54797;
    wire N__54796;
    wire N__54793;
    wire N__54790;
    wire N__54787;
    wire N__54784;
    wire N__54781;
    wire N__54778;
    wire N__54775;
    wire N__54774;
    wire N__54773;
    wire N__54772;
    wire N__54771;
    wire N__54770;
    wire N__54769;
    wire N__54768;
    wire N__54765;
    wire N__54762;
    wire N__54761;
    wire N__54758;
    wire N__54757;
    wire N__54754;
    wire N__54751;
    wire N__54750;
    wire N__54747;
    wire N__54742;
    wire N__54739;
    wire N__54736;
    wire N__54733;
    wire N__54730;
    wire N__54727;
    wire N__54724;
    wire N__54721;
    wire N__54718;
    wire N__54715;
    wire N__54714;
    wire N__54713;
    wire N__54710;
    wire N__54709;
    wire N__54706;
    wire N__54705;
    wire N__54702;
    wire N__54699;
    wire N__54696;
    wire N__54681;
    wire N__54680;
    wire N__54675;
    wire N__54672;
    wire N__54665;
    wire N__54662;
    wire N__54659;
    wire N__54656;
    wire N__54653;
    wire N__54650;
    wire N__54637;
    wire N__54632;
    wire N__54629;
    wire N__54626;
    wire N__54625;
    wire N__54620;
    wire N__54609;
    wire N__54606;
    wire N__54599;
    wire N__54596;
    wire N__54593;
    wire N__54590;
    wire N__54585;
    wire N__54580;
    wire N__54577;
    wire N__54568;
    wire N__54565;
    wire N__54562;
    wire N__54559;
    wire N__54556;
    wire N__54553;
    wire N__54550;
    wire N__54547;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54534;
    wire N__54531;
    wire N__54530;
    wire N__54527;
    wire N__54526;
    wire N__54525;
    wire N__54522;
    wire N__54521;
    wire N__54518;
    wire N__54517;
    wire N__54516;
    wire N__54513;
    wire N__54512;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54505;
    wire N__54502;
    wire N__54501;
    wire N__54500;
    wire N__54499;
    wire N__54498;
    wire N__54497;
    wire N__54494;
    wire N__54491;
    wire N__54488;
    wire N__54485;
    wire N__54482;
    wire N__54481;
    wire N__54480;
    wire N__54477;
    wire N__54474;
    wire N__54473;
    wire N__54470;
    wire N__54469;
    wire N__54466;
    wire N__54463;
    wire N__54460;
    wire N__54457;
    wire N__54454;
    wire N__54451;
    wire N__54450;
    wire N__54449;
    wire N__54446;
    wire N__54445;
    wire N__54442;
    wire N__54441;
    wire N__54438;
    wire N__54437;
    wire N__54434;
    wire N__54433;
    wire N__54426;
    wire N__54423;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54400;
    wire N__54397;
    wire N__54390;
    wire N__54387;
    wire N__54386;
    wire N__54383;
    wire N__54374;
    wire N__54365;
    wire N__54362;
    wire N__54355;
    wire N__54352;
    wire N__54349;
    wire N__54344;
    wire N__54341;
    wire N__54336;
    wire N__54333;
    wire N__54324;
    wire N__54317;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54303;
    wire N__54300;
    wire N__54293;
    wire N__54286;
    wire N__54283;
    wire N__54280;
    wire N__54277;
    wire N__54274;
    wire N__54271;
    wire N__54268;
    wire N__54265;
    wire N__54264;
    wire N__54261;
    wire N__54258;
    wire N__54257;
    wire N__54256;
    wire N__54255;
    wire N__54254;
    wire N__54253;
    wire N__54252;
    wire N__54251;
    wire N__54250;
    wire N__54249;
    wire N__54248;
    wire N__54245;
    wire N__54242;
    wire N__54239;
    wire N__54236;
    wire N__54233;
    wire N__54232;
    wire N__54229;
    wire N__54228;
    wire N__54225;
    wire N__54224;
    wire N__54221;
    wire N__54220;
    wire N__54217;
    wire N__54214;
    wire N__54211;
    wire N__54208;
    wire N__54207;
    wire N__54202;
    wire N__54199;
    wire N__54196;
    wire N__54195;
    wire N__54194;
    wire N__54193;
    wire N__54190;
    wire N__54177;
    wire N__54176;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54166;
    wire N__54163;
    wire N__54160;
    wire N__54157;
    wire N__54156;
    wire N__54153;
    wire N__54148;
    wire N__54145;
    wire N__54142;
    wire N__54139;
    wire N__54138;
    wire N__54137;
    wire N__54136;
    wire N__54135;
    wire N__54132;
    wire N__54129;
    wire N__54126;
    wire N__54123;
    wire N__54120;
    wire N__54111;
    wire N__54108;
    wire N__54105;
    wire N__54100;
    wire N__54091;
    wire N__54088;
    wire N__54085;
    wire N__54084;
    wire N__54081;
    wire N__54080;
    wire N__54077;
    wire N__54070;
    wire N__54063;
    wire N__54060;
    wire N__54055;
    wire N__54046;
    wire N__54043;
    wire N__54038;
    wire N__54033;
    wire N__54028;
    wire N__54025;
    wire N__54016;
    wire N__54013;
    wire N__54010;
    wire N__54007;
    wire N__54004;
    wire N__54001;
    wire N__54000;
    wire N__53999;
    wire N__53996;
    wire N__53993;
    wire N__53992;
    wire N__53991;
    wire N__53990;
    wire N__53987;
    wire N__53986;
    wire N__53983;
    wire N__53980;
    wire N__53977;
    wire N__53974;
    wire N__53971;
    wire N__53970;
    wire N__53969;
    wire N__53966;
    wire N__53963;
    wire N__53958;
    wire N__53955;
    wire N__53952;
    wire N__53949;
    wire N__53946;
    wire N__53943;
    wire N__53942;
    wire N__53941;
    wire N__53940;
    wire N__53939;
    wire N__53938;
    wire N__53937;
    wire N__53934;
    wire N__53931;
    wire N__53922;
    wire N__53919;
    wire N__53916;
    wire N__53915;
    wire N__53912;
    wire N__53911;
    wire N__53908;
    wire N__53907;
    wire N__53904;
    wire N__53903;
    wire N__53900;
    wire N__53897;
    wire N__53894;
    wire N__53889;
    wire N__53888;
    wire N__53887;
    wire N__53886;
    wire N__53885;
    wire N__53884;
    wire N__53883;
    wire N__53882;
    wire N__53881;
    wire N__53876;
    wire N__53873;
    wire N__53870;
    wire N__53867;
    wire N__53854;
    wire N__53851;
    wire N__53848;
    wire N__53845;
    wire N__53842;
    wire N__53839;
    wire N__53836;
    wire N__53833;
    wire N__53832;
    wire N__53829;
    wire N__53826;
    wire N__53823;
    wire N__53820;
    wire N__53819;
    wire N__53816;
    wire N__53805;
    wire N__53802;
    wire N__53799;
    wire N__53796;
    wire N__53785;
    wire N__53778;
    wire N__53775;
    wire N__53772;
    wire N__53769;
    wire N__53766;
    wire N__53757;
    wire N__53754;
    wire N__53743;
    wire N__53740;
    wire N__53737;
    wire N__53734;
    wire N__53731;
    wire N__53728;
    wire N__53725;
    wire N__53724;
    wire N__53723;
    wire N__53722;
    wire N__53719;
    wire N__53716;
    wire N__53715;
    wire N__53712;
    wire N__53711;
    wire N__53708;
    wire N__53707;
    wire N__53706;
    wire N__53705;
    wire N__53702;
    wire N__53699;
    wire N__53696;
    wire N__53695;
    wire N__53694;
    wire N__53693;
    wire N__53690;
    wire N__53687;
    wire N__53684;
    wire N__53681;
    wire N__53680;
    wire N__53677;
    wire N__53674;
    wire N__53669;
    wire N__53666;
    wire N__53665;
    wire N__53662;
    wire N__53661;
    wire N__53658;
    wire N__53657;
    wire N__53654;
    wire N__53651;
    wire N__53650;
    wire N__53647;
    wire N__53644;
    wire N__53641;
    wire N__53638;
    wire N__53637;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53625;
    wire N__53612;
    wire N__53611;
    wire N__53610;
    wire N__53609;
    wire N__53608;
    wire N__53607;
    wire N__53604;
    wire N__53601;
    wire N__53592;
    wire N__53589;
    wire N__53586;
    wire N__53585;
    wire N__53582;
    wire N__53575;
    wire N__53572;
    wire N__53569;
    wire N__53568;
    wire N__53567;
    wire N__53564;
    wire N__53563;
    wire N__53560;
    wire N__53559;
    wire N__53556;
    wire N__53547;
    wire N__53544;
    wire N__53541;
    wire N__53534;
    wire N__53529;
    wire N__53516;
    wire N__53511;
    wire N__53508;
    wire N__53501;
    wire N__53494;
    wire N__53491;
    wire N__53488;
    wire N__53485;
    wire N__53482;
    wire N__53479;
    wire N__53478;
    wire N__53475;
    wire N__53474;
    wire N__53471;
    wire N__53470;
    wire N__53469;
    wire N__53468;
    wire N__53467;
    wire N__53466;
    wire N__53465;
    wire N__53464;
    wire N__53461;
    wire N__53458;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53446;
    wire N__53445;
    wire N__53442;
    wire N__53439;
    wire N__53438;
    wire N__53435;
    wire N__53434;
    wire N__53431;
    wire N__53430;
    wire N__53429;
    wire N__53428;
    wire N__53427;
    wire N__53426;
    wire N__53423;
    wire N__53420;
    wire N__53417;
    wire N__53414;
    wire N__53411;
    wire N__53410;
    wire N__53409;
    wire N__53408;
    wire N__53405;
    wire N__53390;
    wire N__53387;
    wire N__53386;
    wire N__53383;
    wire N__53382;
    wire N__53379;
    wire N__53378;
    wire N__53377;
    wire N__53374;
    wire N__53373;
    wire N__53370;
    wire N__53369;
    wire N__53364;
    wire N__53359;
    wire N__53356;
    wire N__53353;
    wire N__53350;
    wire N__53347;
    wire N__53342;
    wire N__53329;
    wire N__53326;
    wire N__53323;
    wire N__53320;
    wire N__53317;
    wire N__53316;
    wire N__53313;
    wire N__53306;
    wire N__53303;
    wire N__53300;
    wire N__53297;
    wire N__53288;
    wire N__53285;
    wire N__53284;
    wire N__53281;
    wire N__53278;
    wire N__53275;
    wire N__53262;
    wire N__53259;
    wire N__53254;
    wire N__53251;
    wire N__53248;
    wire N__53245;
    wire N__53242;
    wire N__53239;
    wire N__53234;
    wire N__53227;
    wire N__53224;
    wire N__53221;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53211;
    wire N__53210;
    wire N__53207;
    wire N__53206;
    wire N__53203;
    wire N__53202;
    wire N__53201;
    wire N__53200;
    wire N__53199;
    wire N__53198;
    wire N__53197;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53191;
    wire N__53190;
    wire N__53189;
    wire N__53186;
    wire N__53183;
    wire N__53180;
    wire N__53177;
    wire N__53174;
    wire N__53171;
    wire N__53170;
    wire N__53169;
    wire N__53166;
    wire N__53165;
    wire N__53162;
    wire N__53161;
    wire N__53158;
    wire N__53155;
    wire N__53154;
    wire N__53151;
    wire N__53148;
    wire N__53147;
    wire N__53144;
    wire N__53141;
    wire N__53140;
    wire N__53137;
    wire N__53136;
    wire N__53131;
    wire N__53130;
    wire N__53127;
    wire N__53124;
    wire N__53121;
    wire N__53116;
    wire N__53103;
    wire N__53100;
    wire N__53093;
    wire N__53090;
    wire N__53089;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53075;
    wire N__53072;
    wire N__53069;
    wire N__53066;
    wire N__53059;
    wire N__53048;
    wire N__53045;
    wire N__53042;
    wire N__53037;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53020;
    wire N__53013;
    wire N__53010;
    wire N__53005;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52989;
    wire N__52986;
    wire N__52981;
    wire N__52978;
    wire N__52975;
    wire N__52970;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52936;
    wire N__52933;
    wire N__52930;
    wire N__52929;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52919;
    wire N__52912;
    wire N__52909;
    wire N__52906;
    wire N__52903;
    wire N__52900;
    wire N__52897;
    wire N__52894;
    wire N__52891;
    wire N__52888;
    wire N__52885;
    wire N__52882;
    wire N__52879;
    wire N__52876;
    wire N__52875;
    wire N__52874;
    wire N__52867;
    wire N__52864;
    wire N__52861;
    wire N__52858;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52846;
    wire N__52843;
    wire N__52842;
    wire N__52839;
    wire N__52836;
    wire N__52831;
    wire N__52828;
    wire N__52825;
    wire N__52824;
    wire N__52819;
    wire N__52816;
    wire N__52813;
    wire N__52810;
    wire N__52807;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52794;
    wire N__52789;
    wire N__52786;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52772;
    wire N__52767;
    wire N__52764;
    wire N__52759;
    wire N__52756;
    wire N__52755;
    wire N__52750;
    wire N__52747;
    wire N__52746;
    wire N__52745;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52722;
    wire N__52719;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52705;
    wire N__52704;
    wire N__52703;
    wire N__52700;
    wire N__52697;
    wire N__52694;
    wire N__52687;
    wire N__52684;
    wire N__52681;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52657;
    wire N__52654;
    wire N__52651;
    wire N__52650;
    wire N__52645;
    wire N__52642;
    wire N__52641;
    wire N__52640;
    wire N__52637;
    wire N__52634;
    wire N__52631;
    wire N__52624;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52579;
    wire N__52576;
    wire N__52573;
    wire N__52572;
    wire N__52569;
    wire N__52566;
    wire N__52561;
    wire N__52558;
    wire N__52555;
    wire N__52552;
    wire N__52549;
    wire N__52546;
    wire N__52543;
    wire N__52540;
    wire N__52537;
    wire N__52534;
    wire N__52531;
    wire N__52528;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52492;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52453;
    wire N__52450;
    wire N__52447;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52435;
    wire N__52432;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52417;
    wire N__52414;
    wire N__52411;
    wire N__52408;
    wire N__52405;
    wire N__52402;
    wire N__52399;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52344;
    wire N__52341;
    wire N__52338;
    wire N__52333;
    wire N__52330;
    wire N__52327;
    wire N__52324;
    wire N__52321;
    wire N__52318;
    wire N__52315;
    wire N__52312;
    wire N__52309;
    wire N__52306;
    wire N__52303;
    wire N__52300;
    wire N__52297;
    wire N__52294;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52210;
    wire N__52207;
    wire N__52204;
    wire N__52201;
    wire N__52198;
    wire N__52195;
    wire N__52192;
    wire N__52189;
    wire N__52186;
    wire N__52183;
    wire N__52180;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52141;
    wire N__52138;
    wire N__52135;
    wire N__52132;
    wire N__52129;
    wire N__52126;
    wire N__52123;
    wire N__52120;
    wire N__52117;
    wire N__52114;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52062;
    wire N__52059;
    wire N__52056;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52018;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51997;
    wire N__51994;
    wire N__51991;
    wire N__51988;
    wire N__51985;
    wire N__51982;
    wire N__51979;
    wire N__51976;
    wire N__51973;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51946;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51934;
    wire N__51931;
    wire N__51928;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51913;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51901;
    wire N__51898;
    wire N__51895;
    wire N__51892;
    wire N__51889;
    wire N__51886;
    wire N__51883;
    wire N__51880;
    wire N__51877;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51844;
    wire N__51841;
    wire N__51838;
    wire N__51835;
    wire N__51832;
    wire N__51829;
    wire N__51826;
    wire N__51823;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51808;
    wire N__51805;
    wire N__51802;
    wire N__51799;
    wire N__51796;
    wire N__51793;
    wire N__51790;
    wire N__51787;
    wire N__51784;
    wire N__51781;
    wire N__51778;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51748;
    wire N__51745;
    wire N__51742;
    wire N__51739;
    wire N__51736;
    wire N__51733;
    wire N__51730;
    wire N__51727;
    wire N__51724;
    wire N__51721;
    wire N__51718;
    wire N__51715;
    wire N__51712;
    wire N__51709;
    wire N__51706;
    wire N__51703;
    wire N__51700;
    wire N__51697;
    wire N__51694;
    wire N__51691;
    wire N__51688;
    wire N__51685;
    wire N__51682;
    wire N__51679;
    wire N__51676;
    wire N__51673;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51628;
    wire N__51625;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51580;
    wire N__51577;
    wire N__51574;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51541;
    wire N__51538;
    wire N__51535;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51523;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51463;
    wire N__51460;
    wire N__51457;
    wire N__51454;
    wire N__51451;
    wire N__51448;
    wire N__51445;
    wire N__51442;
    wire N__51439;
    wire N__51436;
    wire N__51433;
    wire N__51430;
    wire N__51427;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51388;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51376;
    wire N__51373;
    wire N__51370;
    wire N__51367;
    wire N__51364;
    wire N__51361;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51343;
    wire N__51340;
    wire N__51337;
    wire N__51334;
    wire N__51331;
    wire N__51328;
    wire N__51325;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51313;
    wire N__51310;
    wire N__51307;
    wire N__51304;
    wire N__51301;
    wire N__51298;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51286;
    wire N__51283;
    wire N__51280;
    wire N__51277;
    wire N__51274;
    wire N__51271;
    wire N__51268;
    wire N__51265;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51253;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51214;
    wire N__51211;
    wire N__51208;
    wire N__51205;
    wire N__51204;
    wire N__51201;
    wire N__51198;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51190;
    wire N__51187;
    wire N__51182;
    wire N__51179;
    wire N__51176;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51160;
    wire N__51159;
    wire N__51158;
    wire N__51153;
    wire N__51150;
    wire N__51149;
    wire N__51146;
    wire N__51143;
    wire N__51140;
    wire N__51139;
    wire N__51132;
    wire N__51129;
    wire N__51128;
    wire N__51127;
    wire N__51122;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51108;
    wire N__51105;
    wire N__51102;
    wire N__51097;
    wire N__51094;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51082;
    wire N__51079;
    wire N__51078;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51061;
    wire N__51058;
    wire N__51055;
    wire N__51054;
    wire N__51049;
    wire N__51046;
    wire N__51043;
    wire N__51042;
    wire N__51041;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51025;
    wire N__51022;
    wire N__51021;
    wire N__51018;
    wire N__51015;
    wire N__51010;
    wire N__51009;
    wire N__51008;
    wire N__51005;
    wire N__51002;
    wire N__50999;
    wire N__50996;
    wire N__50993;
    wire N__50990;
    wire N__50983;
    wire N__50980;
    wire N__50977;
    wire N__50976;
    wire N__50975;
    wire N__50972;
    wire N__50967;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50953;
    wire N__50950;
    wire N__50949;
    wire N__50948;
    wire N__50945;
    wire N__50940;
    wire N__50935;
    wire N__50932;
    wire N__50931;
    wire N__50926;
    wire N__50923;
    wire N__50922;
    wire N__50919;
    wire N__50916;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50906;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50890;
    wire N__50887;
    wire N__50884;
    wire N__50881;
    wire N__50878;
    wire N__50877;
    wire N__50874;
    wire N__50873;
    wire N__50870;
    wire N__50867;
    wire N__50862;
    wire N__50859;
    wire N__50856;
    wire N__50851;
    wire N__50848;
    wire N__50845;
    wire N__50842;
    wire N__50839;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50827;
    wire N__50824;
    wire N__50821;
    wire N__50818;
    wire N__50815;
    wire N__50812;
    wire N__50809;
    wire N__50806;
    wire N__50803;
    wire N__50800;
    wire N__50797;
    wire N__50794;
    wire N__50791;
    wire N__50788;
    wire N__50785;
    wire N__50782;
    wire N__50779;
    wire N__50776;
    wire N__50773;
    wire N__50770;
    wire N__50767;
    wire N__50764;
    wire N__50761;
    wire N__50758;
    wire N__50755;
    wire N__50752;
    wire N__50749;
    wire N__50746;
    wire N__50743;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50731;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50719;
    wire N__50716;
    wire N__50713;
    wire N__50712;
    wire N__50709;
    wire N__50708;
    wire N__50703;
    wire N__50700;
    wire N__50697;
    wire N__50694;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50681;
    wire N__50676;
    wire N__50671;
    wire N__50668;
    wire N__50665;
    wire N__50664;
    wire N__50659;
    wire N__50656;
    wire N__50655;
    wire N__50654;
    wire N__50651;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50636;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50620;
    wire N__50617;
    wire N__50614;
    wire N__50611;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50572;
    wire N__50569;
    wire N__50566;
    wire N__50563;
    wire N__50560;
    wire N__50557;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50545;
    wire N__50542;
    wire N__50539;
    wire N__50536;
    wire N__50533;
    wire N__50530;
    wire N__50527;
    wire N__50524;
    wire N__50521;
    wire N__50518;
    wire N__50515;
    wire N__50512;
    wire N__50509;
    wire N__50506;
    wire N__50503;
    wire N__50500;
    wire N__50497;
    wire N__50494;
    wire N__50491;
    wire N__50488;
    wire N__50485;
    wire N__50482;
    wire N__50479;
    wire N__50476;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50455;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50434;
    wire N__50431;
    wire N__50428;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50404;
    wire N__50401;
    wire N__50398;
    wire N__50395;
    wire N__50392;
    wire N__50389;
    wire N__50386;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50364;
    wire N__50363;
    wire N__50362;
    wire N__50359;
    wire N__50354;
    wire N__50351;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50339;
    wire N__50336;
    wire N__50333;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50308;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50155;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50101;
    wire N__50098;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50086;
    wire N__50083;
    wire N__50080;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50011;
    wire N__50008;
    wire N__50005;
    wire N__50002;
    wire N__49999;
    wire N__49996;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49972;
    wire N__49969;
    wire N__49966;
    wire N__49963;
    wire N__49960;
    wire N__49957;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49945;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49927;
    wire N__49924;
    wire N__49921;
    wire N__49918;
    wire N__49915;
    wire N__49912;
    wire N__49909;
    wire N__49906;
    wire N__49903;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49885;
    wire N__49882;
    wire N__49879;
    wire N__49876;
    wire N__49873;
    wire N__49870;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49858;
    wire N__49855;
    wire N__49852;
    wire N__49849;
    wire N__49846;
    wire N__49843;
    wire N__49840;
    wire N__49837;
    wire N__49834;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49811;
    wire N__49808;
    wire N__49803;
    wire N__49798;
    wire N__49795;
    wire N__49794;
    wire N__49791;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49771;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49763;
    wire N__49760;
    wire N__49755;
    wire N__49750;
    wire N__49747;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49702;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49681;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49597;
    wire N__49594;
    wire N__49591;
    wire N__49588;
    wire N__49585;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49543;
    wire N__49540;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49528;
    wire N__49525;
    wire N__49522;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49510;
    wire N__49507;
    wire N__49504;
    wire N__49501;
    wire N__49498;
    wire N__49495;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49462;
    wire N__49459;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49411;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49396;
    wire N__49393;
    wire N__49390;
    wire N__49387;
    wire N__49384;
    wire N__49381;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49357;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49333;
    wire N__49330;
    wire N__49327;
    wire N__49324;
    wire N__49321;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49309;
    wire N__49306;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49273;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49261;
    wire N__49258;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49228;
    wire N__49225;
    wire N__49222;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49165;
    wire N__49162;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49045;
    wire N__49042;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49011;
    wire N__49008;
    wire N__49005;
    wire N__49002;
    wire N__48999;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48962;
    wire N__48959;
    wire N__48956;
    wire N__48953;
    wire N__48952;
    wire N__48947;
    wire N__48944;
    wire N__48941;
    wire N__48940;
    wire N__48939;
    wire N__48936;
    wire N__48931;
    wire N__48926;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48867;
    wire N__48864;
    wire N__48861;
    wire N__48856;
    wire N__48853;
    wire N__48850;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48823;
    wire N__48820;
    wire N__48819;
    wire N__48816;
    wire N__48813;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48793;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48724;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48502;
    wire N__48499;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48379;
    wire N__48376;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48274;
    wire N__48271;
    wire N__48268;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48211;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48187;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48130;
    wire N__48127;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48094;
    wire N__48091;
    wire N__48088;
    wire N__48085;
    wire N__48082;
    wire N__48079;
    wire N__48076;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48064;
    wire N__48061;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48031;
    wire N__48028;
    wire N__48025;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47971;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47944;
    wire N__47941;
    wire N__47938;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47917;
    wire N__47914;
    wire N__47911;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47878;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47845;
    wire N__47842;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47734;
    wire N__47731;
    wire N__47728;
    wire N__47725;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47689;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47679;
    wire N__47676;
    wire N__47673;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47623;
    wire N__47620;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47578;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47503;
    wire N__47500;
    wire N__47497;
    wire N__47494;
    wire N__47491;
    wire N__47488;
    wire N__47485;
    wire N__47482;
    wire N__47479;
    wire N__47476;
    wire N__47473;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47455;
    wire N__47452;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47359;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47338;
    wire N__47335;
    wire N__47332;
    wire N__47329;
    wire N__47326;
    wire N__47323;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47254;
    wire N__47251;
    wire N__47248;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47161;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47065;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46945;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46933;
    wire N__46930;
    wire N__46927;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46897;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46801;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46789;
    wire N__46786;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46774;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46762;
    wire N__46759;
    wire N__46756;
    wire N__46753;
    wire N__46750;
    wire N__46747;
    wire N__46746;
    wire N__46743;
    wire N__46740;
    wire N__46735;
    wire N__46732;
    wire N__46729;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46702;
    wire N__46699;
    wire N__46696;
    wire N__46693;
    wire N__46690;
    wire N__46687;
    wire N__46684;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46639;
    wire N__46636;
    wire N__46633;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46572;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46555;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46542;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46522;
    wire N__46519;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46144;
    wire N__46141;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45997;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45970;
    wire N__45967;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45925;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45901;
    wire N__45898;
    wire N__45895;
    wire N__45892;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45835;
    wire N__45832;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45760;
    wire N__45757;
    wire N__45756;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45738;
    wire N__45735;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45703;
    wire N__45700;
    wire N__45697;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45661;
    wire N__45658;
    wire N__45655;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45643;
    wire N__45640;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45632;
    wire N__45629;
    wire N__45624;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45598;
    wire N__45595;
    wire N__45594;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45582;
    wire N__45579;
    wire N__45576;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45468;
    wire N__45465;
    wire N__45460;
    wire N__45457;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45441;
    wire N__45438;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45382;
    wire N__45379;
    wire N__45376;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45325;
    wire N__45322;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45259;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45151;
    wire N__45148;
    wire N__45147;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45130;
    wire N__45129;
    wire N__45128;
    wire N__45127;
    wire N__45126;
    wire N__45125;
    wire N__45124;
    wire N__45123;
    wire N__45122;
    wire N__45121;
    wire N__45120;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45108;
    wire N__45101;
    wire N__45094;
    wire N__45089;
    wire N__45076;
    wire N__45073;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45055;
    wire N__45052;
    wire N__45051;
    wire N__45050;
    wire N__45049;
    wire N__45048;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45036;
    wire N__45031;
    wire N__45022;
    wire N__45019;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44952;
    wire N__44951;
    wire N__44950;
    wire N__44949;
    wire N__44948;
    wire N__44947;
    wire N__44946;
    wire N__44943;
    wire N__44942;
    wire N__44937;
    wire N__44934;
    wire N__44925;
    wire N__44918;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44908;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44894;
    wire N__44893;
    wire N__44890;
    wire N__44885;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44864;
    wire N__44861;
    wire N__44860;
    wire N__44857;
    wire N__44852;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44840;
    wire N__44833;
    wire N__44832;
    wire N__44829;
    wire N__44828;
    wire N__44827;
    wire N__44824;
    wire N__44823;
    wire N__44822;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44808;
    wire N__44807;
    wire N__44802;
    wire N__44795;
    wire N__44792;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44766;
    wire N__44765;
    wire N__44764;
    wire N__44759;
    wire N__44754;
    wire N__44749;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44737;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44688;
    wire N__44687;
    wire N__44684;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44668;
    wire N__44667;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44440;
    wire N__44437;
    wire N__44436;
    wire N__44435;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44423;
    wire N__44422;
    wire N__44419;
    wire N__44414;
    wire N__44411;
    wire N__44410;
    wire N__44409;
    wire N__44406;
    wire N__44401;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44392;
    wire N__44387;
    wire N__44384;
    wire N__44375;
    wire N__44368;
    wire N__44365;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44353;
    wire N__44350;
    wire N__44349;
    wire N__44346;
    wire N__44341;
    wire N__44340;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44323;
    wire N__44320;
    wire N__44319;
    wire N__44318;
    wire N__44317;
    wire N__44316;
    wire N__44315;
    wire N__44314;
    wire N__44313;
    wire N__44310;
    wire N__44305;
    wire N__44298;
    wire N__44293;
    wire N__44292;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44261;
    wire N__44254;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44242;
    wire N__44241;
    wire N__44240;
    wire N__44239;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44226;
    wire N__44225;
    wire N__44224;
    wire N__44217;
    wire N__44214;
    wire N__44209;
    wire N__44206;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44187;
    wire N__44186;
    wire N__44183;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44167;
    wire N__44166;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44151;
    wire N__44146;
    wire N__44143;
    wire N__44142;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44138;
    wire N__44133;
    wire N__44130;
    wire N__44123;
    wire N__44116;
    wire N__44115;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44091;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44083;
    wire N__44078;
    wire N__44073;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44061;
    wire N__44060;
    wire N__44059;
    wire N__44058;
    wire N__44057;
    wire N__44056;
    wire N__44047;
    wire N__44042;
    wire N__44039;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44007;
    wire N__44004;
    wire N__44003;
    wire N__44000;
    wire N__43995;
    wire N__43992;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43952;
    wire N__43949;
    wire N__43944;
    wire N__43939;
    wire N__43938;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43923;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43833;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43498;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43152;
    wire N__43147;
    wire N__43144;
    wire N__43143;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43131;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43034;
    wire N__43031;
    wire N__43026;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42703;
    wire N__42702;
    wire N__42701;
    wire N__42700;
    wire N__42699;
    wire N__42698;
    wire N__42697;
    wire N__42696;
    wire N__42693;
    wire N__42692;
    wire N__42689;
    wire N__42688;
    wire N__42685;
    wire N__42684;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42666;
    wire N__42653;
    wire N__42648;
    wire N__42645;
    wire N__42634;
    wire N__42633;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42629;
    wire N__42628;
    wire N__42623;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42611;
    wire N__42608;
    wire N__42607;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42596;
    wire N__42595;
    wire N__42594;
    wire N__42593;
    wire N__42590;
    wire N__42585;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42563;
    wire N__42560;
    wire N__42559;
    wire N__42556;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42542;
    wire N__42529;
    wire N__42526;
    wire N__42517;
    wire N__42516;
    wire N__42511;
    wire N__42508;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42463;
    wire N__42460;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42292;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42216;
    wire N__42215;
    wire N__42212;
    wire N__42211;
    wire N__42208;
    wire N__42207;
    wire N__42204;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42190;
    wire N__42187;
    wire N__42186;
    wire N__42185;
    wire N__42184;
    wire N__42183;
    wire N__42182;
    wire N__42179;
    wire N__42164;
    wire N__42161;
    wire N__42150;
    wire N__42147;
    wire N__42146;
    wire N__42143;
    wire N__42142;
    wire N__42139;
    wire N__42138;
    wire N__42137;
    wire N__42136;
    wire N__42135;
    wire N__42134;
    wire N__42131;
    wire N__42130;
    wire N__42127;
    wire N__42120;
    wire N__42107;
    wire N__42104;
    wire N__42103;
    wire N__42100;
    wire N__42099;
    wire N__42096;
    wire N__42095;
    wire N__42092;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42082;
    wire N__42077;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42047;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41977;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41947;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41719;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41709;
    wire N__41708;
    wire N__41707;
    wire N__41704;
    wire N__41701;
    wire N__41700;
    wire N__41697;
    wire N__41696;
    wire N__41693;
    wire N__41692;
    wire N__41691;
    wire N__41690;
    wire N__41689;
    wire N__41688;
    wire N__41687;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41669;
    wire N__41668;
    wire N__41667;
    wire N__41666;
    wire N__41663;
    wire N__41662;
    wire N__41661;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41653;
    wire N__41652;
    wire N__41651;
    wire N__41648;
    wire N__41647;
    wire N__41644;
    wire N__41643;
    wire N__41640;
    wire N__41639;
    wire N__41638;
    wire N__41635;
    wire N__41630;
    wire N__41621;
    wire N__41612;
    wire N__41609;
    wire N__41608;
    wire N__41605;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41597;
    wire N__41584;
    wire N__41579;
    wire N__41572;
    wire N__41569;
    wire N__41556;
    wire N__41551;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41392;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41380;
    wire N__41379;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41356;
    wire N__41355;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41250;
    wire N__41245;
    wire N__41242;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40803;
    wire N__40802;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40674;
    wire N__40671;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40659;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40501;
    wire N__40498;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40486;
    wire N__40485;
    wire N__40484;
    wire N__40481;
    wire N__40476;
    wire N__40475;
    wire N__40470;
    wire N__40467;
    wire N__40462;
    wire N__40459;
    wire N__40458;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40447;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40426;
    wire N__40421;
    wire N__40418;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40404;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40389;
    wire N__40388;
    wire N__40387;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40376;
    wire N__40373;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40360;
    wire N__40357;
    wire N__40356;
    wire N__40353;
    wire N__40352;
    wire N__40351;
    wire N__40350;
    wire N__40349;
    wire N__40348;
    wire N__40345;
    wire N__40332;
    wire N__40327;
    wire N__40314;
    wire N__40313;
    wire N__40312;
    wire N__40311;
    wire N__40308;
    wire N__40307;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40301;
    wire N__40296;
    wire N__40287;
    wire N__40284;
    wire N__40271;
    wire N__40270;
    wire N__40269;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40261;
    wire N__40258;
    wire N__40251;
    wire N__40248;
    wire N__40237;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40120;
    wire N__40117;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39487;
    wire N__39484;
    wire N__39481;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39390;
    wire N__39389;
    wire N__39388;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39384;
    wire N__39381;
    wire N__39380;
    wire N__39377;
    wire N__39376;
    wire N__39373;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39365;
    wire N__39362;
    wire N__39361;
    wire N__39358;
    wire N__39357;
    wire N__39354;
    wire N__39353;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39349;
    wire N__39348;
    wire N__39345;
    wire N__39330;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39287;
    wire N__39286;
    wire N__39283;
    wire N__39282;
    wire N__39279;
    wire N__39278;
    wire N__39275;
    wire N__39274;
    wire N__39271;
    wire N__39264;
    wire N__39257;
    wire N__39252;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39224;
    wire N__39219;
    wire N__39216;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38495;
    wire N__38492;
    wire N__38487;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37758;
    wire N__37757;
    wire N__37756;
    wire N__37755;
    wire N__37754;
    wire N__37753;
    wire N__37752;
    wire N__37751;
    wire N__37750;
    wire N__37749;
    wire N__37746;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37729;
    wire N__37726;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37720;
    wire N__37717;
    wire N__37716;
    wire N__37715;
    wire N__37714;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37700;
    wire N__37697;
    wire N__37696;
    wire N__37693;
    wire N__37680;
    wire N__37675;
    wire N__37662;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37647;
    wire N__37644;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37626;
    wire N__37623;
    wire N__37618;
    wire N__37613;
    wire N__37610;
    wire N__37599;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37429;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36720;
    wire N__36717;
    wire N__36716;
    wire N__36713;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36697;
    wire N__36694;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36681;
    wire N__36680;
    wire N__36679;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36665;
    wire N__36662;
    wire N__36661;
    wire N__36660;
    wire N__36655;
    wire N__36644;
    wire N__36641;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36567;
    wire N__36562;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36468;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36451;
    wire N__36448;
    wire N__36447;
    wire N__36444;
    wire N__36439;
    wire N__36428;
    wire N__36425;
    wire N__36420;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36132;
    wire N__36131;
    wire N__36130;
    wire N__36129;
    wire N__36128;
    wire N__36127;
    wire N__36126;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36111;
    wire N__36108;
    wire N__36107;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36095;
    wire N__36092;
    wire N__36091;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36081;
    wire N__36080;
    wire N__36079;
    wire N__36078;
    wire N__36075;
    wire N__36064;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36034;
    wire N__36033;
    wire N__36030;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36022;
    wire N__36019;
    wire N__36018;
    wire N__36015;
    wire N__36004;
    wire N__35991;
    wire N__35988;
    wire N__35977;
    wire N__35976;
    wire N__35973;
    wire N__35966;
    wire N__35963;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35894;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35884;
    wire N__35883;
    wire N__35880;
    wire N__35879;
    wire N__35876;
    wire N__35875;
    wire N__35872;
    wire N__35871;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35854;
    wire N__35851;
    wire N__35850;
    wire N__35847;
    wire N__35846;
    wire N__35843;
    wire N__35842;
    wire N__35839;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35819;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35793;
    wire N__35778;
    wire N__35775;
    wire N__35770;
    wire N__35767;
    wire N__35766;
    wire N__35763;
    wire N__35762;
    wire N__35759;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35743;
    wire N__35738;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35714;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35003;
    wire N__35000;
    wire N__34995;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34791;
    wire N__34788;
    wire N__34787;
    wire N__34784;
    wire N__34783;
    wire N__34780;
    wire N__34779;
    wire N__34776;
    wire N__34761;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34362;
    wire N__34361;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34349;
    wire N__34346;
    wire N__34339;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34321;
    wire N__34318;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34284;
    wire N__34281;
    wire N__34280;
    wire N__34279;
    wire N__34278;
    wire N__34277;
    wire N__34276;
    wire N__34275;
    wire N__34274;
    wire N__34273;
    wire N__34272;
    wire N__34267;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34246;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34236;
    wire N__34233;
    wire N__34232;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34224;
    wire N__34223;
    wire N__34222;
    wire N__34221;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34201;
    wire N__34192;
    wire N__34179;
    wire N__34174;
    wire N__34173;
    wire N__34170;
    wire N__34169;
    wire N__34166;
    wire N__34165;
    wire N__34162;
    wire N__34151;
    wire N__34146;
    wire N__34133;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34083;
    wire N__34078;
    wire N__34075;
    wire N__34074;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33500;
    wire N__33497;
    wire N__33496;
    wire N__33495;
    wire N__33490;
    wire N__33479;
    wire N__33476;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33348;
    wire N__33347;
    wire N__33346;
    wire N__33345;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33331;
    wire N__33328;
    wire N__33327;
    wire N__33324;
    wire N__33319;
    wire N__33308;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32852;
    wire N__32849;
    wire N__32848;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32805;
    wire N__32804;
    wire N__32801;
    wire N__32800;
    wire N__32799;
    wire N__32798;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32770;
    wire N__32767;
    wire N__32766;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32728;
    wire N__32725;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32697;
    wire N__32694;
    wire N__32693;
    wire N__32688;
    wire N__32683;
    wire N__32680;
    wire N__32673;
    wire N__32670;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32608;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32600;
    wire N__32597;
    wire N__32592;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32445;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32377;
    wire N__32376;
    wire N__32373;
    wire N__32372;
    wire N__32371;
    wire N__32370;
    wire N__32369;
    wire N__32368;
    wire N__32367;
    wire N__32366;
    wire N__32365;
    wire N__32364;
    wire N__32363;
    wire N__32360;
    wire N__32353;
    wire N__32352;
    wire N__32343;
    wire N__32340;
    wire N__32339;
    wire N__32336;
    wire N__32335;
    wire N__32332;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32323;
    wire N__32320;
    wire N__32319;
    wire N__32318;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32285;
    wire N__32280;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32260;
    wire N__32249;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32205;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32193;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32181;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32169;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32157;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32136;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32126;
    wire N__32125;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32110;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32093;
    wire N__32090;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32078;
    wire N__32073;
    wire N__32066;
    wire N__32059;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32041;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31926;
    wire N__31923;
    wire N__31922;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31824;
    wire N__31821;
    wire N__31820;
    wire N__31817;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31781;
    wire N__31778;
    wire N__31777;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31753;
    wire N__31748;
    wire N__31747;
    wire N__31740;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31734;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31716;
    wire N__31715;
    wire N__31714;
    wire N__31711;
    wire N__31706;
    wire N__31693;
    wire N__31688;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31572;
    wire N__31571;
    wire N__31570;
    wire N__31569;
    wire N__31568;
    wire N__31567;
    wire N__31564;
    wire N__31563;
    wire N__31562;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31547;
    wire N__31536;
    wire N__31529;
    wire N__31520;
    wire N__31519;
    wire N__31518;
    wire N__31511;
    wire N__31510;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31501;
    wire N__31500;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31496;
    wire N__31495;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31488;
    wire N__31473;
    wire N__31472;
    wire N__31469;
    wire N__31468;
    wire N__31465;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31440;
    wire N__31439;
    wire N__31434;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31406;
    wire N__31397;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31315;
    wire N__31314;
    wire N__31311;
    wire N__31310;
    wire N__31307;
    wire N__31306;
    wire N__31291;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31194;
    wire N__31193;
    wire N__31192;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31178;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31154;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30849;
    wire N__30848;
    wire N__30847;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30840;
    wire N__30839;
    wire N__30838;
    wire N__30837;
    wire N__30834;
    wire N__30833;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30825;
    wire N__30822;
    wire N__30821;
    wire N__30820;
    wire N__30817;
    wire N__30812;
    wire N__30809;
    wire N__30808;
    wire N__30805;
    wire N__30804;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30796;
    wire N__30791;
    wire N__30778;
    wire N__30773;
    wire N__30770;
    wire N__30765;
    wire N__30764;
    wire N__30751;
    wire N__30748;
    wire N__30743;
    wire N__30738;
    wire N__30735;
    wire N__30734;
    wire N__30731;
    wire N__30722;
    wire N__30719;
    wire N__30712;
    wire N__30711;
    wire N__30708;
    wire N__30707;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30676;
    wire N__30673;
    wire N__30672;
    wire N__30669;
    wire N__30668;
    wire N__30665;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30627;
    wire N__30624;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30612;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30278;
    wire N__30273;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29673;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29662;
    wire N__29659;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29633;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29610;
    wire N__29609;
    wire N__29606;
    wire N__29605;
    wire N__29602;
    wire N__29601;
    wire N__29598;
    wire N__29597;
    wire N__29596;
    wire N__29595;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29553;
    wire N__29552;
    wire N__29551;
    wire N__29548;
    wire N__29547;
    wire N__29544;
    wire N__29543;
    wire N__29540;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29534;
    wire N__29533;
    wire N__29532;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29510;
    wire N__29507;
    wire N__29506;
    wire N__29503;
    wire N__29502;
    wire N__29499;
    wire N__29498;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29473;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29442;
    wire N__29441;
    wire N__29440;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29426;
    wire N__29423;
    wire N__29422;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29402;
    wire N__29399;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29277;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28755;
    wire N__28752;
    wire N__28751;
    wire N__28750;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire pin3_clk_16mhz_pad_gb_input;
    wire VCCG0;
    wire bfn_6_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336 ;
    wire bfn_6_21_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177 ;
    wire bfn_7_19_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448 ;
    wire bfn_7_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338 ;
    wire bfn_7_21_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138 ;
    wire bfn_7_22_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252 ;
    wire bfn_7_23_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478 ;
    wire bfn_7_24_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341 ;
    wire bfn_7_25_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141 ;
    wire bfn_7_26_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256 ;
    wire bfn_9_9_0_;
    wire \foc.u_Park_Transform.n17107 ;
    wire \foc.u_Park_Transform.n17108 ;
    wire \foc.u_Park_Transform.n17109 ;
    wire \foc.u_Park_Transform.n17110 ;
    wire \foc.u_Park_Transform.n17111 ;
    wire \foc.u_Park_Transform.n17112 ;
    wire \foc.u_Park_Transform.n17113 ;
    wire \foc.u_Park_Transform.n17114 ;
    wire bfn_9_10_0_;
    wire \foc.u_Park_Transform.n17115 ;
    wire \foc.u_Park_Transform.n17116 ;
    wire \foc.u_Park_Transform.n779_adj_2070 ;
    wire bfn_9_11_0_;
    wire \foc.u_Park_Transform.n81 ;
    wire \foc.u_Park_Transform.n17118 ;
    wire \foc.u_Park_Transform.n130 ;
    wire \foc.u_Park_Transform.n17119 ;
    wire \foc.u_Park_Transform.n179 ;
    wire \foc.u_Park_Transform.n17120 ;
    wire \foc.u_Park_Transform.n228_adj_2063 ;
    wire \foc.u_Park_Transform.n17121 ;
    wire \foc.u_Park_Transform.n277_adj_2060 ;
    wire \foc.u_Park_Transform.n17122 ;
    wire \foc.u_Park_Transform.n326_adj_2056 ;
    wire \foc.u_Park_Transform.n17123 ;
    wire \foc.u_Park_Transform.n375_adj_2055 ;
    wire \foc.u_Park_Transform.n17124 ;
    wire \foc.u_Park_Transform.n17125 ;
    wire \foc.u_Park_Transform.n424_adj_2052 ;
    wire bfn_9_12_0_;
    wire \foc.u_Park_Transform.n473_adj_2050 ;
    wire \foc.u_Park_Transform.n17126 ;
    wire \foc.u_Park_Transform.n17127 ;
    wire \foc.u_Park_Transform.n17128 ;
    wire \foc.u_Park_Transform.n522_adj_2046 ;
    wire \foc.u_Park_Transform.n17129 ;
    wire \foc.u_Park_Transform.n775_adj_2047 ;
    wire bfn_9_15_0_;
    wire \foc.u_Park_Transform.n16935 ;
    wire \foc.u_Park_Transform.n16936 ;
    wire \foc.u_Park_Transform.n16937 ;
    wire \foc.u_Park_Transform.n16938 ;
    wire \foc.u_Park_Transform.n16939 ;
    wire \foc.u_Park_Transform.n16940 ;
    wire \foc.u_Park_Transform.n16941 ;
    wire \foc.u_Park_Transform.n16942 ;
    wire bfn_9_16_0_;
    wire \foc.u_Park_Transform.n16943 ;
    wire \foc.u_Park_Transform.n16944 ;
    wire \foc.u_Park_Transform.n16945 ;
    wire \foc.u_Park_Transform.n16946 ;
    wire \foc.u_Park_Transform.n775 ;
    wire bfn_9_19_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467 ;
    wire bfn_9_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471 ;
    wire bfn_9_21_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831 ;
    wire bfn_9_22_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244 ;
    wire bfn_9_23_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347 ;
    wire bfn_9_24_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147 ;
    wire bfn_9_25_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489 ;
    wire bfn_10_9_0_;
    wire \foc.u_Park_Transform.n17146 ;
    wire \foc.u_Park_Transform.n17147 ;
    wire \foc.u_Park_Transform.n17148 ;
    wire \foc.u_Park_Transform.n17149 ;
    wire \foc.u_Park_Transform.n17150 ;
    wire \foc.u_Park_Transform.n17151 ;
    wire \foc.u_Park_Transform.n17152 ;
    wire \foc.u_Park_Transform.n17153 ;
    wire bfn_10_10_0_;
    wire \foc.u_Park_Transform.n17154 ;
    wire \foc.u_Park_Transform.n17155 ;
    wire \foc.u_Park_Transform.n17156 ;
    wire \foc.u_Park_Transform.n17157 ;
    wire \foc.u_Park_Transform.n17158 ;
    wire \foc.u_Park_Transform.n17159 ;
    wire \foc.u_Park_Transform.n767 ;
    wire \foc.u_Park_Transform.n75 ;
    wire bfn_10_11_0_;
    wire \foc.u_Park_Transform.n78 ;
    wire \foc.u_Park_Transform.n124 ;
    wire \foc.u_Park_Transform.n17131 ;
    wire \foc.u_Park_Transform.n127 ;
    wire \foc.u_Park_Transform.n173 ;
    wire \foc.u_Park_Transform.n17132 ;
    wire \foc.u_Park_Transform.n176 ;
    wire \foc.u_Park_Transform.n222 ;
    wire \foc.u_Park_Transform.n17133 ;
    wire \foc.u_Park_Transform.n225 ;
    wire \foc.u_Park_Transform.n271 ;
    wire \foc.u_Park_Transform.n17134 ;
    wire \foc.u_Park_Transform.n274 ;
    wire \foc.u_Park_Transform.n320 ;
    wire \foc.u_Park_Transform.n17135 ;
    wire \foc.u_Park_Transform.n323 ;
    wire \foc.u_Park_Transform.n369 ;
    wire \foc.u_Park_Transform.n17136 ;
    wire \foc.u_Park_Transform.n372 ;
    wire \foc.u_Park_Transform.n418_adj_2024 ;
    wire \foc.u_Park_Transform.n17137 ;
    wire \foc.u_Park_Transform.n17138 ;
    wire \foc.u_Park_Transform.n421_adj_2039 ;
    wire \foc.u_Park_Transform.n467_adj_2019 ;
    wire bfn_10_12_0_;
    wire \foc.u_Park_Transform.n470_adj_2038 ;
    wire \foc.u_Park_Transform.n516_adj_2018 ;
    wire \foc.u_Park_Transform.n17139 ;
    wire \foc.u_Park_Transform.n519_adj_2035 ;
    wire \foc.u_Park_Transform.n565 ;
    wire \foc.u_Park_Transform.n17140 ;
    wire \foc.u_Park_Transform.n568_adj_2034 ;
    wire \foc.u_Park_Transform.n614_adj_2017 ;
    wire \foc.u_Park_Transform.n17141 ;
    wire \foc.u_Park_Transform.n663_adj_2016 ;
    wire \foc.u_Park_Transform.n17142 ;
    wire \foc.u_Park_Transform.n712_adj_2015 ;
    wire \foc.u_Park_Transform.n17143 ;
    wire \foc.u_Park_Transform.n617_adj_2031 ;
    wire \foc.u_Park_Transform.n17144 ;
    wire \foc.u_Park_Transform.n771_adj_2032 ;
    wire \foc.u_Park_Transform.n773 ;
    wire bfn_10_14_0_;
    wire \foc.u_Park_Transform.n18160 ;
    wire \foc.u_Park_Transform.n18161 ;
    wire \foc.u_Park_Transform.n18162 ;
    wire \foc.u_Park_Transform.n18163 ;
    wire \foc.u_Park_Transform.n18164 ;
    wire \foc.u_Park_Transform.n18165 ;
    wire \foc.u_Park_Transform.n787 ;
    wire bfn_10_15_0_;
    wire \foc.u_Park_Transform.n87 ;
    wire \foc.u_Park_Transform.n16915 ;
    wire \foc.u_Park_Transform.n136 ;
    wire \foc.u_Park_Transform.n16916 ;
    wire \foc.u_Park_Transform.n185 ;
    wire \foc.u_Park_Transform.n16917 ;
    wire \foc.u_Park_Transform.n234 ;
    wire \foc.u_Park_Transform.n16918 ;
    wire \foc.u_Park_Transform.n283 ;
    wire \foc.u_Park_Transform.n16919 ;
    wire \foc.u_Park_Transform.n16920 ;
    wire \foc.u_Park_Transform.n16921 ;
    wire \foc.u_Park_Transform.n16922 ;
    wire \foc.u_Park_Transform.n332 ;
    wire bfn_10_16_0_;
    wire \foc.u_Park_Transform.n783_adj_2167 ;
    wire \foc.u_Park_Transform.n81_adj_2120 ;
    wire bfn_10_17_0_;
    wire \foc.u_Park_Transform.n84_adj_2118 ;
    wire \foc.u_Park_Transform.n130_adj_2105 ;
    wire \foc.u_Park_Transform.n16924 ;
    wire \foc.u_Park_Transform.n133 ;
    wire \foc.u_Park_Transform.n179_adj_2076 ;
    wire \foc.u_Park_Transform.n16925 ;
    wire \foc.u_Park_Transform.n182 ;
    wire \foc.u_Park_Transform.n228 ;
    wire \foc.u_Park_Transform.n16926 ;
    wire \foc.u_Park_Transform.n231 ;
    wire \foc.u_Park_Transform.n277 ;
    wire \foc.u_Park_Transform.n16927 ;
    wire \foc.u_Park_Transform.n280 ;
    wire \foc.u_Park_Transform.n326 ;
    wire \foc.u_Park_Transform.n16928 ;
    wire \foc.u_Park_Transform.n329 ;
    wire \foc.u_Park_Transform.n375 ;
    wire \foc.u_Park_Transform.n16929 ;
    wire \foc.u_Park_Transform.n378 ;
    wire \foc.u_Park_Transform.n424 ;
    wire \foc.u_Park_Transform.n16930 ;
    wire \foc.u_Park_Transform.n16931 ;
    wire \foc.u_Park_Transform.n473 ;
    wire bfn_10_18_0_;
    wire \foc.u_Park_Transform.n619 ;
    wire \foc.u_Park_Transform.n522 ;
    wire \foc.u_Park_Transform.n16932 ;
    wire \foc.u_Park_Transform.n777 ;
    wire \foc.u_Park_Transform.n427 ;
    wire \foc.u_Park_Transform.n16933 ;
    wire \foc.u_Park_Transform.n779 ;
    wire bfn_10_19_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392 ;
    wire bfn_10_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224 ;
    wire bfn_10_21_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828 ;
    wire bfn_10_22_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420 ;
    wire bfn_10_23_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401 ;
    wire bfn_10_24_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228 ;
    wire bfn_10_25_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ;
    wire bfn_10_26_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465 ;
    wire \foc.u_Park_Transform.n84 ;
    wire bfn_11_9_0_;
    wire \foc.u_Park_Transform.n133_adj_2101 ;
    wire \foc.u_Park_Transform.n17098 ;
    wire \foc.u_Park_Transform.n182_adj_2094 ;
    wire \foc.u_Park_Transform.n17099 ;
    wire \foc.u_Park_Transform.n231_adj_2089 ;
    wire \foc.u_Park_Transform.n17100 ;
    wire \foc.u_Park_Transform.n280_adj_2087 ;
    wire \foc.u_Park_Transform.n17101 ;
    wire \foc.u_Park_Transform.n329_adj_2080 ;
    wire \foc.u_Park_Transform.n17102 ;
    wire \foc.u_Park_Transform.n378_adj_2078 ;
    wire \foc.u_Park_Transform.n17103 ;
    wire \foc.u_Park_Transform.n427_adj_2069 ;
    wire \foc.u_Park_Transform.n17104 ;
    wire \foc.u_Park_Transform.n17105 ;
    wire bfn_11_10_0_;
    wire \foc.u_Park_Transform.n783 ;
    wire \foc.u_Park_Transform.n622 ;
    wire \foc.u_Park_Transform.n781 ;
    wire \foc.u_Park_Transform.n87_adj_2138 ;
    wire bfn_11_11_0_;
    wire \foc.u_Park_Transform.n136_adj_2127 ;
    wire \foc.u_Park_Transform.n17980 ;
    wire \foc.u_Park_Transform.n185_adj_2126 ;
    wire \foc.u_Park_Transform.n17981 ;
    wire \foc.u_Park_Transform.n234_adj_2125 ;
    wire \foc.u_Park_Transform.n17982 ;
    wire \foc.u_Park_Transform.n283_adj_2122 ;
    wire \foc.u_Park_Transform.n17983 ;
    wire \foc.u_Park_Transform.n332_adj_2110 ;
    wire \foc.u_Park_Transform.n17984 ;
    wire \foc.u_Park_Transform.n17985 ;
    wire \foc.u_Park_Transform.n787_adj_2149 ;
    wire \foc.u_Park_Transform.n625 ;
    wire n21486_cascade_;
    wire n139;
    wire \foc.u_Park_Transform.n90 ;
    wire bfn_11_13_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946 ;
    wire \foc.Look_Up_Table_out1_1_6 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947 ;
    wire \foc.Look_Up_Table_out1_1_7 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948 ;
    wire \foc.Look_Up_Table_out1_1_8 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949 ;
    wire \foc.Look_Up_Table_out1_1_9 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951 ;
    wire \foc.Look_Up_Table_out1_1_10 ;
    wire bfn_11_14_0_;
    wire \foc.Look_Up_Table_out1_1_11 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956 ;
    wire \foc.Look_Up_Table_out1_1_12 ;
    wire \foc.u_Park_Transform.n785 ;
    wire \foc.u_Park_Transform.n616 ;
    wire bfn_11_15_0_;
    wire \foc.u_Park_Transform.n78_adj_2145 ;
    wire \foc.u_Park_Transform.n16948 ;
    wire \foc.u_Park_Transform.n127_adj_2119 ;
    wire \foc.u_Park_Transform.n16949 ;
    wire \foc.u_Park_Transform.n176_adj_2104 ;
    wire \foc.u_Park_Transform.n16950 ;
    wire \foc.u_Park_Transform.n225_adj_2075 ;
    wire \foc.u_Park_Transform.n16951 ;
    wire \foc.u_Park_Transform.n274_adj_2058 ;
    wire \foc.u_Park_Transform.n16952 ;
    wire \foc.u_Park_Transform.n323_adj_2057 ;
    wire \foc.u_Park_Transform.n16953 ;
    wire \foc.u_Park_Transform.n372_adj_2042 ;
    wire \foc.u_Park_Transform.n16954 ;
    wire \foc.u_Park_Transform.n16955 ;
    wire \foc.u_Park_Transform.n421 ;
    wire bfn_11_16_0_;
    wire \foc.u_Park_Transform.n470 ;
    wire \foc.u_Park_Transform.n16956 ;
    wire \foc.u_Park_Transform.n519 ;
    wire \foc.u_Park_Transform.n16957 ;
    wire \foc.u_Park_Transform.n568 ;
    wire \foc.u_Park_Transform.n16958 ;
    wire \foc.u_Park_Transform.n16959 ;
    wire \foc.u_Park_Transform.n16960 ;
    wire \foc.u_Park_Transform.n769 ;
    wire \foc.u_Park_Transform.n617 ;
    wire \foc.u_Park_Transform.n16961 ;
    wire \foc.u_Park_Transform.n771 ;
    wire bfn_11_17_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365 ;
    wire bfn_11_18_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ;
    wire bfn_11_19_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40 ;
    wire bfn_11_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329 ;
    wire bfn_11_21_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235 ;
    wire bfn_11_22_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423 ;
    wire bfn_11_23_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231 ;
    wire bfn_11_24_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO ;
    wire bfn_12_9_0_;
    wire \foc.u_Park_Transform.n72 ;
    wire \foc.u_Park_Transform.n17161 ;
    wire \foc.u_Park_Transform.n121 ;
    wire \foc.u_Park_Transform.n17162 ;
    wire \foc.u_Park_Transform.n170 ;
    wire \foc.u_Park_Transform.n17163 ;
    wire \foc.u_Park_Transform.n219 ;
    wire \foc.u_Park_Transform.n17164 ;
    wire \foc.u_Park_Transform.n268 ;
    wire \foc.u_Park_Transform.n17165 ;
    wire \foc.u_Park_Transform.n317 ;
    wire \foc.u_Park_Transform.n17166 ;
    wire \foc.u_Park_Transform.n366 ;
    wire \foc.u_Park_Transform.n17167 ;
    wire \foc.u_Park_Transform.n17168 ;
    wire \foc.u_Park_Transform.n415_adj_2008 ;
    wire bfn_12_10_0_;
    wire \foc.u_Park_Transform.n464_adj_2005 ;
    wire \foc.u_Park_Transform.n17169 ;
    wire \foc.u_Park_Transform.n513_adj_2002 ;
    wire \foc.u_Park_Transform.n17170 ;
    wire \foc.u_Park_Transform.n562_adj_2000 ;
    wire \foc.u_Park_Transform.n17171 ;
    wire \foc.u_Park_Transform.n611 ;
    wire \foc.u_Park_Transform.n17172 ;
    wire \foc.u_Park_Transform.n660 ;
    wire \foc.u_Park_Transform.n17173 ;
    wire \foc.u_Park_Transform.n709 ;
    wire \foc.u_Park_Transform.n17174 ;
    wire \foc.u_Park_Transform.n763 ;
    wire bfn_12_11_0_;
    wire \foc.u_Park_Transform.n69 ;
    wire \foc.u_Park_Transform.n17176 ;
    wire \foc.u_Park_Transform.n118 ;
    wire \foc.u_Park_Transform.n17177 ;
    wire \foc.u_Park_Transform.n167 ;
    wire \foc.u_Park_Transform.n17178 ;
    wire \foc.u_Park_Transform.n216 ;
    wire \foc.u_Park_Transform.n17179 ;
    wire \foc.u_Park_Transform.n265 ;
    wire \foc.u_Park_Transform.n17180 ;
    wire \foc.u_Park_Transform.n314 ;
    wire \foc.u_Park_Transform.n17181 ;
    wire \foc.u_Park_Transform.n363 ;
    wire \foc.u_Park_Transform.n17182 ;
    wire \foc.u_Park_Transform.n17183 ;
    wire \foc.u_Park_Transform.n412 ;
    wire bfn_12_12_0_;
    wire \foc.u_Park_Transform.n461 ;
    wire \foc.u_Park_Transform.n17184 ;
    wire \foc.u_Park_Transform.n510_adj_2004 ;
    wire \foc.u_Park_Transform.n17185 ;
    wire \foc.u_Park_Transform.n559_adj_2001 ;
    wire \foc.u_Park_Transform.n17186 ;
    wire \foc.u_Park_Transform.n608 ;
    wire \foc.u_Park_Transform.n17187 ;
    wire \foc.u_Park_Transform.n657 ;
    wire \foc.u_Park_Transform.n17188 ;
    wire \foc.u_Park_Transform.n706 ;
    wire \foc.u_Park_Transform.n17189 ;
    wire \foc.u_Park_Transform.n759_adj_2166 ;
    wire \foc.Look_Up_Table_out1_1_3 ;
    wire \foc.Look_Up_Table_out1_1_5 ;
    wire \foc.Look_Up_Table_out1_1_4 ;
    wire n4_cascade_;
    wire \foc.u_Park_Transform.n237 ;
    wire \foc.u_Park_Transform.n188 ;
    wire \foc.u_Park_Transform.n613 ;
    wire bfn_12_15_0_;
    wire \foc.u_Park_Transform.n75_adj_2123 ;
    wire \foc.u_Park_Transform.n16963 ;
    wire \foc.u_Park_Transform.n124_adj_2090 ;
    wire \foc.u_Park_Transform.n16964 ;
    wire \foc.u_Park_Transform.n173_adj_2061 ;
    wire \foc.u_Park_Transform.n16965 ;
    wire \foc.u_Park_Transform.n222_adj_2049 ;
    wire \foc.u_Park_Transform.n16966 ;
    wire \foc.u_Park_Transform.n271_adj_2043 ;
    wire \foc.u_Park_Transform.n16967 ;
    wire \foc.u_Park_Transform.n320_adj_2036 ;
    wire \foc.u_Park_Transform.n16968 ;
    wire \foc.u_Park_Transform.n369_adj_2026 ;
    wire \foc.u_Park_Transform.n16969 ;
    wire \foc.u_Park_Transform.n16970 ;
    wire \foc.u_Park_Transform.n418 ;
    wire bfn_12_16_0_;
    wire \foc.u_Park_Transform.n467 ;
    wire \foc.u_Park_Transform.n16971 ;
    wire \foc.u_Park_Transform.n516 ;
    wire \foc.u_Park_Transform.n16972 ;
    wire \foc.u_Park_Transform.n565_adj_2020 ;
    wire \foc.u_Park_Transform.n16973 ;
    wire \foc.u_Park_Transform.n614 ;
    wire \foc.u_Park_Transform.n16974 ;
    wire \foc.u_Park_Transform.n663 ;
    wire \foc.u_Park_Transform.n16975 ;
    wire \foc.u_Park_Transform.n765 ;
    wire \foc.u_Park_Transform.n712 ;
    wire \foc.u_Park_Transform.n16976 ;
    wire \foc.u_Park_Transform.n767_adj_2041 ;
    wire bfn_12_17_0_;
    wire \foc.u_Park_Transform.n16900 ;
    wire \foc.u_Park_Transform.n16901 ;
    wire \foc.u_Park_Transform.n16902 ;
    wire \foc.u_Park_Transform.n16903 ;
    wire \foc.u_Park_Transform.n16904 ;
    wire \foc.u_Park_Transform.n16905 ;
    wire \foc.u_Park_Transform.n16906 ;
    wire \foc.u_Park_Transform.n16907 ;
    wire \foc.u_Park_Transform.n766_adj_2053 ;
    wire bfn_12_18_0_;
    wire \foc.u_Park_Transform.n770 ;
    wire \foc.u_Park_Transform.n767_adj_2041_THRU_CO ;
    wire \foc.u_Park_Transform.n16908 ;
    wire \foc.u_Park_Transform.n774 ;
    wire \foc.u_Park_Transform.n771_THRU_CO ;
    wire \foc.u_Park_Transform.n16909 ;
    wire \foc.u_Park_Transform.n778 ;
    wire \foc.u_Park_Transform.n775_THRU_CO ;
    wire \foc.u_Park_Transform.n16910 ;
    wire \foc.u_Park_Transform.n782 ;
    wire \foc.u_Park_Transform.n779_THRU_CO ;
    wire \foc.u_Park_Transform.n16911 ;
    wire \foc.u_Park_Transform.n786 ;
    wire \foc.u_Park_Transform.n783_adj_2167_THRU_CO ;
    wire \foc.u_Park_Transform.n16912 ;
    wire \foc.u_Park_Transform.n787_THRU_CO ;
    wire \foc.u_Park_Transform.n16913 ;
    wire \foc.u_Park_Transform.n16914 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816 ;
    wire bfn_12_19_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219 ;
    wire bfn_12_20_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO ;
    wire bfn_12_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17656 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17657 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17658 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17659 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17660 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17661 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17662 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17663 ;
    wire bfn_12_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17664 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17665 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17666 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17667 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n775 ;
    wire bfn_12_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18107 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18108 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18109 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18110 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18111 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18112 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n372 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18113 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18114 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n421 ;
    wire bfn_12_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n470 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18115 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n519 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18116 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n568 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18117 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18118 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18119 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n617 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18120 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598 ;
    wire bfn_13_9_0_;
    wire \foc.u_Park_Transform.n17083 ;
    wire \foc.u_Park_Transform.n17084 ;
    wire \foc.u_Park_Transform.n17085 ;
    wire \foc.u_Park_Transform.n17086 ;
    wire \foc.u_Park_Transform.n17087 ;
    wire \foc.u_Park_Transform.n758_adj_2168 ;
    wire \foc.u_Park_Transform.n17088 ;
    wire \foc.u_Park_Transform.n759_adj_2166_THRU_CO ;
    wire \foc.u_Park_Transform.n762 ;
    wire \foc.u_Park_Transform.n17089 ;
    wire \foc.u_Park_Transform.n17090 ;
    wire \foc.u_Park_Transform.n766 ;
    wire \foc.u_Park_Transform.n763_THRU_CO ;
    wire bfn_13_10_0_;
    wire \foc.u_Park_Transform.n770_adj_2030 ;
    wire \foc.u_Park_Transform.n767_THRU_CO ;
    wire \foc.u_Park_Transform.n17091 ;
    wire \foc.u_Park_Transform.n774_adj_2045 ;
    wire \foc.u_Park_Transform.n771_adj_2032_THRU_CO ;
    wire \foc.u_Park_Transform.n17092 ;
    wire \foc.u_Park_Transform.n778_adj_2068 ;
    wire \foc.u_Park_Transform.n775_adj_2047_THRU_CO ;
    wire \foc.u_Park_Transform.n17093 ;
    wire \foc.u_Park_Transform.n782_adj_2109 ;
    wire \foc.u_Park_Transform.n779_adj_2070_THRU_CO ;
    wire \foc.u_Park_Transform.n17094 ;
    wire \foc.u_Park_Transform.n786_adj_2152 ;
    wire \foc.u_Park_Transform.n783_THRU_CO ;
    wire \foc.u_Park_Transform.n17095 ;
    wire \foc.u_Park_Transform.n790 ;
    wire \foc.u_Park_Transform.n787_adj_2149_THRU_CO ;
    wire \foc.u_Park_Transform.n17096 ;
    wire \foc.u_Park_Transform.n17097 ;
    wire bfn_13_11_0_;
    wire \foc.u_Park_Transform.n66 ;
    wire \foc.u_Park_Transform.n17191 ;
    wire \foc.u_Park_Transform.n115 ;
    wire \foc.u_Park_Transform.n17192 ;
    wire \foc.u_Park_Transform.n164 ;
    wire \foc.u_Park_Transform.n17193 ;
    wire \foc.u_Park_Transform.n213 ;
    wire \foc.u_Park_Transform.n17194 ;
    wire \foc.u_Park_Transform.n262_adj_1996 ;
    wire \foc.u_Park_Transform.n17195 ;
    wire \foc.u_Park_Transform.n311 ;
    wire \foc.u_Park_Transform.n17196 ;
    wire \foc.u_Park_Transform.n360 ;
    wire \foc.u_Park_Transform.n17197 ;
    wire \foc.u_Park_Transform.n17198 ;
    wire \foc.u_Park_Transform.n409 ;
    wire bfn_13_12_0_;
    wire \foc.u_Park_Transform.n458 ;
    wire \foc.u_Park_Transform.n17199 ;
    wire \foc.u_Park_Transform.n507_adj_2165 ;
    wire \foc.u_Park_Transform.n17200 ;
    wire \foc.u_Park_Transform.n556_adj_2164 ;
    wire \foc.u_Park_Transform.n17201 ;
    wire \foc.u_Park_Transform.n605_adj_2163 ;
    wire \foc.u_Park_Transform.n17202 ;
    wire \foc.u_Park_Transform.n654_adj_2162 ;
    wire \foc.u_Park_Transform.n17203 ;
    wire \foc.u_Park_Transform.n703_adj_2160 ;
    wire \foc.u_Park_Transform.n754_adj_2159 ;
    wire \foc.u_Park_Transform.n17204 ;
    wire \foc.u_Park_Transform.n755_adj_2161 ;
    wire \foc.u_Park_Transform.n755_adj_2161_THRU_CO ;
    wire bfn_13_13_0_;
    wire \foc.u_Park_Transform.n16993 ;
    wire \foc.u_Park_Transform.n16994 ;
    wire \foc.u_Park_Transform.n16995 ;
    wire \foc.u_Park_Transform.n16996 ;
    wire \foc.u_Park_Transform.n16997 ;
    wire \foc.u_Park_Transform.n16998 ;
    wire \foc.u_Park_Transform.n16999 ;
    wire \foc.u_Park_Transform.n17000 ;
    wire bfn_13_14_0_;
    wire \foc.u_Park_Transform.n17001 ;
    wire \foc.u_Park_Transform.n17002 ;
    wire \foc.u_Park_Transform.n17003 ;
    wire \foc.u_Park_Transform.n17004 ;
    wire \foc.u_Park_Transform.n17005 ;
    wire \foc.u_Park_Transform.n757 ;
    wire \foc.u_Park_Transform.n758 ;
    wire \foc.u_Park_Transform.n17006 ;
    wire \foc.u_Park_Transform.n759 ;
    wire \foc.u_Park_Transform.n759_THRU_CO ;
    wire \foc.u_Park_Transform.n610 ;
    wire \foc.u_Park_Transform.n69_adj_2059 ;
    wire bfn_13_15_0_;
    wire \foc.u_Park_Transform.n72_adj_2062 ;
    wire \foc.u_Park_Transform.n118_adj_2037 ;
    wire \foc.u_Park_Transform.n16978 ;
    wire \foc.u_Park_Transform.n121_adj_2051 ;
    wire \foc.u_Park_Transform.n167_adj_2029 ;
    wire \foc.u_Park_Transform.n16979 ;
    wire \foc.u_Park_Transform.n170_adj_2048 ;
    wire \foc.u_Park_Transform.n216_adj_2025 ;
    wire \foc.u_Park_Transform.n16980 ;
    wire \foc.u_Park_Transform.n219_adj_2040 ;
    wire \foc.u_Park_Transform.n265_adj_2023 ;
    wire \foc.u_Park_Transform.n16981 ;
    wire \foc.u_Park_Transform.n268_adj_2027 ;
    wire \foc.u_Park_Transform.n314_adj_2010 ;
    wire \foc.u_Park_Transform.n16982 ;
    wire \foc.u_Park_Transform.n317_adj_2021 ;
    wire \foc.u_Park_Transform.n363_adj_1998 ;
    wire \foc.u_Park_Transform.n16983 ;
    wire \foc.u_Park_Transform.n366_adj_2013 ;
    wire \foc.u_Park_Transform.n412_adj_1995 ;
    wire \foc.u_Park_Transform.n16984 ;
    wire \foc.u_Park_Transform.n16985 ;
    wire \foc.u_Park_Transform.n415 ;
    wire \foc.u_Park_Transform.n461_adj_2007 ;
    wire bfn_13_16_0_;
    wire \foc.u_Park_Transform.n464 ;
    wire \foc.u_Park_Transform.n510 ;
    wire \foc.u_Park_Transform.n16986 ;
    wire \foc.u_Park_Transform.n513 ;
    wire \foc.u_Park_Transform.n559 ;
    wire \foc.u_Park_Transform.n16987 ;
    wire \foc.u_Park_Transform.n562 ;
    wire \foc.u_Park_Transform.n608_adj_2067 ;
    wire \foc.u_Park_Transform.n16988 ;
    wire \foc.u_Park_Transform.n611_adj_2107 ;
    wire \foc.u_Park_Transform.n657_adj_2064 ;
    wire \foc.u_Park_Transform.n16989 ;
    wire \foc.u_Park_Transform.n660_adj_2091 ;
    wire \foc.u_Park_Transform.n607 ;
    wire \foc.u_Park_Transform.n706_adj_2044 ;
    wire \foc.u_Park_Transform.n16990 ;
    wire \foc.u_Park_Transform.n761 ;
    wire \foc.u_Park_Transform.n709_adj_2066 ;
    wire \foc.u_Park_Transform.n762_adj_2065 ;
    wire \foc.u_Park_Transform.n16991 ;
    wire \foc.u_Park_Transform.n763_adj_2054 ;
    wire \foc.u_Park_Transform.n763_adj_2054_THRU_CO ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411 ;
    wire bfn_13_17_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215 ;
    wire bfn_13_18_0_;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216 ;
    wire \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO ;
    wire \foc.Look_Up_Table_out1_1_0 ;
    wire n794;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750 ;
    wire bfn_13_20_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17856 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17857 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17858 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17859 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n326 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17860 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n375 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17861 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n424 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17862 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17863 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n473 ;
    wire bfn_13_21_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n522 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17864 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17865 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736 ;
    wire bfn_13_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17957 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17958 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17959 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17960 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17961 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17962 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17963 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17964 ;
    wire bfn_13_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17965 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n774 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17966 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17967 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17968 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17969 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17970 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17971 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17972 ;
    wire bfn_13_24_0_;
    wire bfn_13_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18092 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18093 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18094 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18095 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18096 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18097 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18098 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18099 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605 ;
    wire bfn_13_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18100 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18101 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18102 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18103 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18104 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18105 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO ;
    wire \foc.dCurrent_4 ;
    wire bfn_14_7_0_;
    wire \foc.dCurrent_5 ;
    wire \foc.u_Park_Transform.n17277 ;
    wire \foc.dCurrent_6 ;
    wire \foc.u_Park_Transform.n17278 ;
    wire \foc.dCurrent_7 ;
    wire \foc.u_Park_Transform.n17279 ;
    wire \foc.dCurrent_8 ;
    wire \foc.u_Park_Transform.n17280 ;
    wire \foc.dCurrent_9 ;
    wire \foc.u_Park_Transform.n17281 ;
    wire \foc.dCurrent_10 ;
    wire \foc.u_Park_Transform.n17282 ;
    wire \foc.dCurrent_11 ;
    wire \foc.u_Park_Transform.n17283 ;
    wire \foc.u_Park_Transform.n17284 ;
    wire \foc.dCurrent_12 ;
    wire bfn_14_8_0_;
    wire \foc.dCurrent_13 ;
    wire \foc.u_Park_Transform.n17285 ;
    wire \foc.dCurrent_14 ;
    wire \foc.u_Park_Transform.n17286 ;
    wire \foc.dCurrent_15 ;
    wire \foc.u_Park_Transform.n17287 ;
    wire \foc.dCurrent_16 ;
    wire \foc.u_Park_Transform.n17288 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_15 ;
    wire \foc.dCurrent_17 ;
    wire \foc.u_Park_Transform.n17289 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_16 ;
    wire \foc.dCurrent_18 ;
    wire \foc.u_Park_Transform.n17290 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_17 ;
    wire \foc.dCurrent_19 ;
    wire \foc.u_Park_Transform.n17291 ;
    wire \foc.u_Park_Transform.n17292 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_18 ;
    wire \foc.dCurrent_20 ;
    wire bfn_14_9_0_;
    wire \foc.u_Park_Transform.Product1_mul_temp_19 ;
    wire \foc.dCurrent_21 ;
    wire \foc.u_Park_Transform.n17293 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_20 ;
    wire \foc.dCurrent_22 ;
    wire \foc.u_Park_Transform.n17294 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_21 ;
    wire \foc.dCurrent_23 ;
    wire \foc.u_Park_Transform.n17295 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_22 ;
    wire \foc.dCurrent_24 ;
    wire \foc.u_Park_Transform.n17296 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_23 ;
    wire \foc.dCurrent_25 ;
    wire \foc.u_Park_Transform.n17297 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_24 ;
    wire \foc.u_Park_Transform.n17298 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_25 ;
    wire \foc.u_Park_Transform.n17299 ;
    wire \foc.u_Park_Transform.n17300 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_26 ;
    wire bfn_14_10_0_;
    wire \foc.u_Park_Transform.Product1_mul_temp_27 ;
    wire \foc.u_Park_Transform.n17301 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_28 ;
    wire \foc.u_Park_Transform.n17302 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_29 ;
    wire \foc.u_Park_Transform.n17303 ;
    wire \foc.dCurrent_31_cascade_ ;
    wire \foc.dCurrent_29 ;
    wire \foc.dCurrent_28 ;
    wire \foc.dCurrent_30 ;
    wire bfn_14_11_0_;
    wire \foc.u_Park_Transform.n17221 ;
    wire \foc.u_Park_Transform.n17222 ;
    wire \foc.u_Park_Transform.n17223 ;
    wire \foc.u_Park_Transform.n17224 ;
    wire \foc.u_Park_Transform.n17225 ;
    wire \foc.u_Park_Transform.n17226 ;
    wire \foc.u_Park_Transform.n17227 ;
    wire \foc.u_Park_Transform.n17228 ;
    wire bfn_14_12_0_;
    wire \foc.u_Park_Transform.n17229 ;
    wire \foc.u_Park_Transform.n17230 ;
    wire \foc.u_Park_Transform.n17231 ;
    wire \foc.u_Park_Transform.n17232 ;
    wire \foc.u_Park_Transform.n17233 ;
    wire \foc.u_Park_Transform.n746 ;
    wire \foc.u_Park_Transform.n17234 ;
    wire \foc.u_Park_Transform.n747 ;
    wire \foc.u_Park_Transform.n747_THRU_CO ;
    wire \foc.u_Park_Transform.n604 ;
    wire bfn_14_13_0_;
    wire \foc.u_Park_Transform.n66_adj_2033 ;
    wire \foc.u_Park_Transform.n17008 ;
    wire \foc.u_Park_Transform.n115_adj_2028 ;
    wire \foc.u_Park_Transform.n17009 ;
    wire \foc.u_Park_Transform.n164_adj_2014 ;
    wire \foc.u_Park_Transform.n17010 ;
    wire \foc.u_Park_Transform.n213_adj_1999 ;
    wire \foc.u_Park_Transform.n17011 ;
    wire \foc.u_Park_Transform.n262 ;
    wire \foc.u_Park_Transform.n17012 ;
    wire \foc.u_Park_Transform.n311_adj_2022 ;
    wire \foc.u_Park_Transform.n17013 ;
    wire \foc.u_Park_Transform.n360_adj_2009 ;
    wire \foc.u_Park_Transform.n17014 ;
    wire \foc.u_Park_Transform.n17015 ;
    wire \foc.u_Park_Transform.n409_adj_1997 ;
    wire bfn_14_14_0_;
    wire \foc.u_Park_Transform.n458_adj_2093 ;
    wire \foc.u_Park_Transform.n17016 ;
    wire \foc.u_Park_Transform.n507 ;
    wire \foc.u_Park_Transform.n17017 ;
    wire \foc.u_Park_Transform.n556 ;
    wire \foc.u_Park_Transform.n17018 ;
    wire \foc.u_Park_Transform.n605 ;
    wire \foc.u_Park_Transform.n17019 ;
    wire \foc.u_Park_Transform.n654 ;
    wire \foc.u_Park_Transform.n17020 ;
    wire \foc.u_Park_Transform.n753 ;
    wire \foc.u_Park_Transform.n703 ;
    wire \foc.u_Park_Transform.n754 ;
    wire \foc.u_Park_Transform.n17021 ;
    wire \foc.u_Park_Transform.n755 ;
    wire \foc.u_Park_Transform.n755_THRU_CO ;
    wire bfn_14_15_0_;
    wire \foc.u_Park_Transform.n17068 ;
    wire \foc.u_Park_Transform.n17069 ;
    wire \foc.u_Park_Transform.n17070 ;
    wire \foc.u_Park_Transform.n17071 ;
    wire \foc.u_Park_Transform.n17072 ;
    wire \foc.u_Park_Transform.n17073 ;
    wire \foc.u_Park_Transform.n17074 ;
    wire \foc.u_Park_Transform.n17075 ;
    wire bfn_14_16_0_;
    wire \foc.u_Park_Transform.n17076 ;
    wire \foc.u_Park_Transform.n17077 ;
    wire \foc.u_Park_Transform.n17078 ;
    wire \foc.u_Park_Transform.n17079 ;
    wire \foc.u_Park_Transform.n17080 ;
    wire \foc.u_Park_Transform.n738_adj_2003 ;
    wire \foc.u_Park_Transform.n17081 ;
    wire \foc.u_Park_Transform.n739_adj_2006 ;
    wire \foc.u_Park_Transform.n739_adj_2006_THRU_CO ;
    wire \foc.u_Park_Transform.Product4_mul_temp_2 ;
    wire bfn_14_17_0_;
    wire \foc.u_Park_Transform.Product4_mul_temp_3 ;
    wire \foc.u_Park_Transform.n15748 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_4 ;
    wire \foc.u_Park_Transform.n15749 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_5 ;
    wire \foc.u_Park_Transform.n15750 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_6 ;
    wire \foc.u_Park_Transform.n15751 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_7 ;
    wire \foc.u_Park_Transform.n15752 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_8 ;
    wire \foc.u_Park_Transform.n15753 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_9 ;
    wire \foc.u_Park_Transform.n15754 ;
    wire \foc.u_Park_Transform.n15755 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_10 ;
    wire bfn_14_18_0_;
    wire \foc.u_Park_Transform.Product4_mul_temp_11 ;
    wire \foc.u_Park_Transform.n15756 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_12 ;
    wire \foc.u_Park_Transform.n15757 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_13 ;
    wire \foc.u_Park_Transform.n15758 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_14 ;
    wire \foc.u_Park_Transform.n15759 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_15 ;
    wire \foc.u_Park_Transform.n15760 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_16 ;
    wire \foc.u_Park_Transform.n15761 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_17 ;
    wire \foc.u_Park_Transform.n15762 ;
    wire \foc.u_Park_Transform.n15763 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_18 ;
    wire bfn_14_19_0_;
    wire \foc.u_Park_Transform.Product4_mul_temp_19 ;
    wire \foc.u_Park_Transform.n15764 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_20 ;
    wire \foc.u_Park_Transform.n15765 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_21 ;
    wire \foc.u_Park_Transform.n15766 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_22 ;
    wire \foc.u_Park_Transform.n15767 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_23 ;
    wire \foc.u_Park_Transform.n15768 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_24 ;
    wire \foc.u_Park_Transform.n15769 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_25 ;
    wire \foc.u_Park_Transform.n15770 ;
    wire \foc.u_Park_Transform.n15771 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_26 ;
    wire bfn_14_20_0_;
    wire \foc.u_Park_Transform.Product4_mul_temp_27 ;
    wire \foc.u_Park_Transform.n15772 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_28 ;
    wire \foc.u_Park_Transform.n15773 ;
    wire \foc.u_Park_Transform.Product4_mul_temp_29 ;
    wire \foc.u_Park_Transform.n15774 ;
    wire \foc.qCurrent_21 ;
    wire \foc.qCurrent_29 ;
    wire \foc.qCurrent_23 ;
    wire \foc.qCurrent_30 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749 ;
    wire bfn_14_21_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17727 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17728 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17729 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17730 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17731 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17732 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17733 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17734 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735 ;
    wire bfn_14_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO ;
    wire bfn_14_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18047 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18048 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18049 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18050 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18051 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18052 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18053 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18054 ;
    wire bfn_14_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18055 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18056 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18057 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18058 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18059 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18060 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO ;
    wire bfn_14_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18032 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18033 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18034 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18035 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18036 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18037 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18038 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18039 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675 ;
    wire bfn_14_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18040 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18041 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18042 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18043 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18044 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18045 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO ;
    wire bfn_15_5_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15775 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n30 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15776 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n29 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15777 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n28 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15778 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15779 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15780 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15781 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15782 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n24 ;
    wire bfn_15_6_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n23 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15783 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n22 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15784 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15785 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15786 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15787 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15788 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15789 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15790 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n16 ;
    wire bfn_15_7_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15791 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15792 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n13 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15793 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15794 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n11 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15795 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n10 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15796 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15797 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15798 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n8 ;
    wire bfn_15_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15799 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15800 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n5 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15801 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15802 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n3 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15803 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n2 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15804 ;
    wire \foc.dCurrent_26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n7 ;
    wire \foc.dCurrent_3 ;
    wire bfn_15_9_0_;
    wire \foc.u_Park_Transform.Product1_mul_temp_2 ;
    wire \foc.u_Park_Transform.n17251 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_3 ;
    wire \foc.u_Park_Transform.n17252 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_4 ;
    wire \foc.u_Park_Transform.n17253 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_5 ;
    wire \foc.u_Park_Transform.n17254 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_6 ;
    wire \foc.u_Park_Transform.n17255 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_7 ;
    wire \foc.u_Park_Transform.n17256 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_8 ;
    wire \foc.u_Park_Transform.n17257 ;
    wire \foc.u_Park_Transform.n17258 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_9 ;
    wire bfn_15_10_0_;
    wire \foc.u_Park_Transform.Product1_mul_temp_10 ;
    wire \foc.u_Park_Transform.n17259 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_11 ;
    wire \foc.u_Park_Transform.n17260 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_12 ;
    wire \foc.u_Park_Transform.n17261 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_13 ;
    wire \foc.u_Park_Transform.n17262 ;
    wire \foc.u_Park_Transform.dCurrent_2 ;
    wire \foc.u_Park_Transform.Product1_mul_temp_14 ;
    wire \foc.u_Park_Transform.n17263 ;
    wire \foc.u_Park_Transform.n737 ;
    wire \foc.u_Park_Transform.n738 ;
    wire \foc.u_Park_Transform.n17264 ;
    wire \foc.u_Park_Transform.n739 ;
    wire \foc.u_Park_Transform.n739_THRU_CO ;
    wire \foc.u_Park_Transform.n54_adj_2095 ;
    wire bfn_15_11_0_;
    wire \foc.u_Park_Transform.n57_adj_2116 ;
    wire \foc.u_Park_Transform.n103_adj_2092 ;
    wire \foc.u_Park_Transform.n17236 ;
    wire \foc.u_Park_Transform.n106_adj_2115 ;
    wire \foc.u_Park_Transform.n152_adj_2088 ;
    wire \foc.u_Park_Transform.n17237 ;
    wire \foc.u_Park_Transform.n155_adj_2114 ;
    wire \foc.u_Park_Transform.n201_adj_2085 ;
    wire \foc.u_Park_Transform.n17238 ;
    wire \foc.u_Park_Transform.n204_adj_2113 ;
    wire \foc.u_Park_Transform.n250_adj_2084 ;
    wire \foc.u_Park_Transform.n17239 ;
    wire \foc.u_Park_Transform.n253_adj_2112 ;
    wire \foc.u_Park_Transform.n299_adj_2083 ;
    wire \foc.u_Park_Transform.n17240 ;
    wire \foc.u_Park_Transform.n302_adj_2111 ;
    wire \foc.u_Park_Transform.n348_adj_2082 ;
    wire \foc.u_Park_Transform.n17241 ;
    wire \foc.u_Park_Transform.n351_adj_2108 ;
    wire \foc.u_Park_Transform.n397_adj_2081 ;
    wire \foc.u_Park_Transform.n17242 ;
    wire \foc.u_Park_Transform.n17243 ;
    wire \foc.u_Park_Transform.n400_adj_2106 ;
    wire \foc.u_Park_Transform.n446_adj_2079 ;
    wire bfn_15_12_0_;
    wire \foc.u_Park_Transform.n449_adj_2103 ;
    wire \foc.u_Park_Transform.n495_adj_2077 ;
    wire \foc.u_Park_Transform.n17244 ;
    wire \foc.u_Park_Transform.n498_adj_2102 ;
    wire \foc.u_Park_Transform.n544_adj_2074 ;
    wire \foc.u_Park_Transform.n17245 ;
    wire \foc.u_Park_Transform.n547_adj_2100 ;
    wire \foc.u_Park_Transform.n593_adj_2073 ;
    wire \foc.u_Park_Transform.n17246 ;
    wire \foc.u_Park_Transform.n596_adj_2099 ;
    wire \foc.u_Park_Transform.n642_adj_2072 ;
    wire \foc.u_Park_Transform.n17247 ;
    wire \foc.u_Park_Transform.n645_adj_2098 ;
    wire \foc.u_Park_Transform.n691_adj_2071 ;
    wire \foc.u_Park_Transform.n17248 ;
    wire \foc.u_Park_Transform.n694_adj_2097 ;
    wire \foc.u_Park_Transform.n742 ;
    wire \foc.u_Park_Transform.n17249 ;
    wire \foc.u_Park_Transform.n743 ;
    wire \foc.u_Park_Transform.n743_THRU_CO ;
    wire bfn_15_13_0_;
    wire \foc.u_Park_Transform.n63 ;
    wire \foc.u_Park_Transform.n17023 ;
    wire \foc.u_Park_Transform.n112 ;
    wire \foc.u_Park_Transform.n17024 ;
    wire \foc.u_Park_Transform.n161 ;
    wire \foc.u_Park_Transform.n17025 ;
    wire \foc.u_Park_Transform.n210 ;
    wire \foc.u_Park_Transform.n17026 ;
    wire \foc.u_Park_Transform.n259 ;
    wire \foc.u_Park_Transform.n17027 ;
    wire \foc.u_Park_Transform.n308 ;
    wire \foc.u_Park_Transform.n17028 ;
    wire \foc.u_Park_Transform.n357 ;
    wire \foc.u_Park_Transform.n17029 ;
    wire \foc.u_Park_Transform.n17030 ;
    wire \foc.u_Park_Transform.n406 ;
    wire bfn_15_14_0_;
    wire \foc.u_Park_Transform.n455 ;
    wire \foc.u_Park_Transform.n17031 ;
    wire \foc.u_Park_Transform.n504 ;
    wire \foc.u_Park_Transform.n17032 ;
    wire \foc.u_Park_Transform.n553 ;
    wire \foc.u_Park_Transform.n17033 ;
    wire \foc.u_Park_Transform.n602 ;
    wire \foc.u_Park_Transform.n17034 ;
    wire \foc.u_Park_Transform.n651 ;
    wire \foc.u_Park_Transform.n17035 ;
    wire \foc.u_Park_Transform.n700 ;
    wire \foc.u_Park_Transform.n750_adj_2117 ;
    wire \foc.u_Park_Transform.n17036 ;
    wire \foc.u_Park_Transform.n751 ;
    wire \foc.u_Park_Transform.n751_THRU_CO ;
    wire \foc.u_Park_Transform.n54 ;
    wire bfn_15_15_0_;
    wire \foc.u_Park_Transform.n103 ;
    wire \foc.u_Park_Transform.n17053 ;
    wire \foc.u_Park_Transform.n152 ;
    wire \foc.u_Park_Transform.n17054 ;
    wire \foc.u_Park_Transform.n201 ;
    wire \foc.u_Park_Transform.n17055 ;
    wire \foc.u_Park_Transform.n250 ;
    wire \foc.u_Park_Transform.n17056 ;
    wire \foc.u_Park_Transform.n299 ;
    wire \foc.u_Park_Transform.n17057 ;
    wire \foc.u_Park_Transform.n348 ;
    wire \foc.u_Park_Transform.n17058 ;
    wire \foc.u_Park_Transform.n397 ;
    wire \foc.u_Park_Transform.n17059 ;
    wire \foc.u_Park_Transform.n17060 ;
    wire \foc.u_Park_Transform.n446 ;
    wire bfn_15_16_0_;
    wire \foc.u_Park_Transform.n495 ;
    wire \foc.u_Park_Transform.n17061 ;
    wire \foc.u_Park_Transform.n544 ;
    wire \foc.u_Park_Transform.n17062 ;
    wire \foc.u_Park_Transform.n593 ;
    wire \foc.u_Park_Transform.n17063 ;
    wire \foc.u_Park_Transform.n642 ;
    wire \foc.u_Park_Transform.n17064 ;
    wire \foc.u_Park_Transform.n691 ;
    wire \foc.u_Park_Transform.n17065 ;
    wire \foc.u_Park_Transform.n742_adj_2086 ;
    wire \foc.u_Park_Transform.n17066 ;
    wire \foc.u_Park_Transform.n743_adj_2096 ;
    wire \foc.u_Park_Transform.n743_adj_2096_THRU_CO ;
    wire \foc.qCurrent_6 ;
    wire \foc.u_Park_Transform.n741 ;
    wire Look_Up_Table_out1_1_14;
    wire Look_Up_Table_out1_1_15;
    wire \foc.qCurrent_8 ;
    wire \foc.Look_Up_Table_out1_1_1 ;
    wire \foc.u_Park_Transform.n592 ;
    wire \foc.qCurrent_3 ;
    wire \foc.qCurrent_18 ;
    wire \foc.qCurrent_19 ;
    wire \foc.qCurrent_13 ;
    wire \foc.qCurrent_16 ;
    wire \foc.qCurrent_14 ;
    wire \foc.qCurrent_4 ;
    wire \foc.qCurrent_11 ;
    wire \foc.qCurrent_15 ;
    wire \foc.qCurrent_22 ;
    wire \foc.qCurrent_17 ;
    wire \foc.qCurrent_24 ;
    wire \foc.qCurrent_27 ;
    wire \foc.qCurrent_26 ;
    wire \foc.qCurrent_12 ;
    wire \foc.qCurrent_28 ;
    wire \foc.qCurrent_20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_ ;
    wire \foc.qCurrent_31 ;
    wire \foc.qCurrent_25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730 ;
    wire bfn_15_21_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17973 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17974 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17975 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17976 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17977 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17978 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733 ;
    wire n794_adj_2425;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666 ;
    wire bfn_15_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18062 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18063 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18064 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18065 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18066 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18067 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18068 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18069 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658 ;
    wire bfn_15_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18070 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18071 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18072 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18073 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18074 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18075 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650 ;
    wire bfn_15_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18077 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18078 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18079 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18080 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18081 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18082 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18083 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18084 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642 ;
    wire bfn_15_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18085 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18086 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18087 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18088 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18089 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18090 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24 ;
    wire \foc.dCurrent_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n6 ;
    wire \foc.u_Park_Transform.n601 ;
    wire \foc.u_Park_Transform.n60_adj_2140 ;
    wire bfn_16_11_0_;
    wire \foc.u_Park_Transform.n63_adj_2158 ;
    wire \foc.u_Park_Transform.n109_adj_2139 ;
    wire \foc.u_Park_Transform.n17206 ;
    wire \foc.u_Park_Transform.n112_adj_2157 ;
    wire \foc.u_Park_Transform.n158_adj_2137 ;
    wire \foc.u_Park_Transform.n17207 ;
    wire \foc.u_Park_Transform.n161_adj_2156 ;
    wire \foc.u_Park_Transform.n207_adj_2136 ;
    wire \foc.u_Park_Transform.n17208 ;
    wire \foc.u_Park_Transform.n210_adj_2155 ;
    wire \foc.u_Park_Transform.n256_adj_2135 ;
    wire \foc.u_Park_Transform.n17209 ;
    wire \foc.u_Park_Transform.n259_adj_2154 ;
    wire \foc.u_Park_Transform.n305_adj_2134 ;
    wire \foc.u_Park_Transform.n17210 ;
    wire \foc.u_Park_Transform.n308_adj_2153 ;
    wire \foc.u_Park_Transform.n354_adj_2133 ;
    wire \foc.u_Park_Transform.n17211 ;
    wire \foc.u_Park_Transform.n357_adj_2151 ;
    wire \foc.u_Park_Transform.n403_adj_2132 ;
    wire \foc.u_Park_Transform.n17212 ;
    wire \foc.u_Park_Transform.n17213 ;
    wire \foc.u_Park_Transform.n406_adj_2150 ;
    wire \foc.u_Park_Transform.n452_adj_2131 ;
    wire bfn_16_12_0_;
    wire \foc.u_Park_Transform.n455_adj_2148 ;
    wire \foc.u_Park_Transform.n501_adj_2130 ;
    wire \foc.u_Park_Transform.n17214 ;
    wire \foc.u_Park_Transform.n504_adj_2147 ;
    wire \foc.u_Park_Transform.n550_adj_2129 ;
    wire \foc.u_Park_Transform.n17215 ;
    wire \foc.u_Park_Transform.n553_adj_2146 ;
    wire \foc.u_Park_Transform.n599_adj_2128 ;
    wire \foc.u_Park_Transform.n17216 ;
    wire \foc.u_Park_Transform.n602_adj_2144 ;
    wire \foc.u_Park_Transform.n648_adj_2124 ;
    wire \foc.u_Park_Transform.n17217 ;
    wire \foc.u_Park_Transform.n651_adj_2143 ;
    wire \foc.u_Park_Transform.n697_adj_2121 ;
    wire \foc.u_Park_Transform.n17218 ;
    wire \foc.u_Park_Transform.n749 ;
    wire \foc.u_Park_Transform.n700_adj_2141 ;
    wire \foc.u_Park_Transform.n750 ;
    wire \foc.u_Park_Transform.n17219 ;
    wire \foc.u_Park_Transform.n751_adj_2142 ;
    wire \foc.u_Park_Transform.n751_adj_2142_THRU_CO ;
    wire \foc.u_Park_Transform.n598 ;
    wire \foc.u_Park_Transform.n57 ;
    wire bfn_16_13_0_;
    wire \foc.u_Park_Transform.n60 ;
    wire \foc.u_Park_Transform.n106 ;
    wire \foc.u_Park_Transform.n17038 ;
    wire \foc.u_Park_Transform.n109 ;
    wire \foc.u_Park_Transform.n155 ;
    wire \foc.u_Park_Transform.n17039 ;
    wire \foc.u_Park_Transform.n158 ;
    wire \foc.u_Park_Transform.n204 ;
    wire \foc.u_Park_Transform.n17040 ;
    wire \foc.u_Park_Transform.n207 ;
    wire \foc.u_Park_Transform.n253 ;
    wire \foc.u_Park_Transform.n17041 ;
    wire \foc.u_Park_Transform.n256 ;
    wire \foc.u_Park_Transform.n302 ;
    wire \foc.u_Park_Transform.n17042 ;
    wire \foc.u_Park_Transform.n305 ;
    wire \foc.u_Park_Transform.n351 ;
    wire \foc.u_Park_Transform.n17043 ;
    wire \foc.u_Park_Transform.n354 ;
    wire \foc.u_Park_Transform.n400 ;
    wire \foc.u_Park_Transform.n17044 ;
    wire \foc.u_Park_Transform.n17045 ;
    wire \foc.u_Park_Transform.n403 ;
    wire \foc.u_Park_Transform.n449 ;
    wire bfn_16_14_0_;
    wire \foc.u_Park_Transform.n452 ;
    wire \foc.u_Park_Transform.n498 ;
    wire \foc.u_Park_Transform.n17046 ;
    wire \foc.u_Park_Transform.n501 ;
    wire \foc.u_Park_Transform.n547 ;
    wire \foc.u_Park_Transform.n17047 ;
    wire \foc.u_Park_Transform.n550 ;
    wire \foc.u_Park_Transform.n596 ;
    wire \foc.u_Park_Transform.n17048 ;
    wire \foc.u_Park_Transform.n599 ;
    wire \foc.u_Park_Transform.n645 ;
    wire \foc.u_Park_Transform.n17049 ;
    wire \foc.u_Park_Transform.n648 ;
    wire \foc.u_Park_Transform.n694 ;
    wire \foc.u_Park_Transform.n17050 ;
    wire \foc.u_Park_Transform.n745 ;
    wire \foc.u_Park_Transform.n697 ;
    wire \foc.u_Park_Transform.n746_adj_2011 ;
    wire \foc.u_Park_Transform.n17051 ;
    wire \foc.u_Park_Transform.n747_adj_2012 ;
    wire \foc.u_Park_Transform.n747_adj_2012_THRU_CO ;
    wire \foc.u_Park_Transform.n6_cascade_ ;
    wire \foc.Look_Up_Table_out1_1_2 ;
    wire \foc.u_Park_Transform.n595 ;
    wire n4;
    wire \foc.qCurrent_10 ;
    wire \foc.qCurrent_7 ;
    wire \foc.qCurrent_5 ;
    wire \foc.qCurrent_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n30 ;
    wire \foc.u_DQ_Current_Control.n31 ;
    wire bfn_16_18_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n29 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15720 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n28 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15721 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15722 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n26 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15723 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15724 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n24 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15725 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n23 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15726 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15727 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n22 ;
    wire bfn_16_19_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15728 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15729 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15730 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15731 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15732 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n16 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15733 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15734 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15735 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n14 ;
    wire bfn_16_20_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n13 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15736 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n12 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15737 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n11 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15738 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n10 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15739 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15740 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n8 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15741 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n7 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15742 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15743 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n6 ;
    wire bfn_16_21_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n5 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15744 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n4 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15745 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n3 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15746 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n2 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15747 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22 ;
    wire bfn_16_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17987 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17988 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17989 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17990 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17991 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17992 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17993 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17994 ;
    wire bfn_16_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17995 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17996 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17997 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17998 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n17999 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18000 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n739 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO ;
    wire bfn_16_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18017 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18018 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18019 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18020 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18021 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18022 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18023 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18024 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691 ;
    wire bfn_16_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18025 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18026 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18027 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18028 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18029 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18030 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n54 ;
    wire bfn_16_27_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n103 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18002 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n152 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18003 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n201 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18004 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n250 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18005 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n299 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18006 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n348 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18007 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n397 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18008 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18009 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n446 ;
    wire bfn_16_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n495 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18010 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n544 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18011 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n593 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18012 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n642 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18013 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18014 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18015 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO ;
    wire bfn_17_5_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18135 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18136 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18137 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18138 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18139 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18140 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18141 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18142 ;
    wire bfn_17_6_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400 ;
    wire bfn_17_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n90 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18167 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18168 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18169 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n283 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18170 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n332 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18171 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18172 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n787 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n188 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n139 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n237 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n4 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n12 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19273 ;
    wire n142_adj_2419;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19269 ;
    wire \foc.u_Park_Transform.n7_cascade_ ;
    wire \foc.u_Park_Transform.n791 ;
    wire \foc.u_Park_Transform.n4_cascade_ ;
    wire Look_Up_Table_out1_1_13;
    wire \foc.u_Park_Transform.n14 ;
    wire n628_cascade_;
    wire \foc.u_Park_Transform.n12 ;
    wire n142;
    wire n628;
    wire \foc.u_Park_Transform.n18_cascade_ ;
    wire \foc.u_Park_Transform.n19845 ;
    wire \foc.u_Park_Transform.n26 ;
    wire bfn_17_15_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17781 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17782 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17783 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17784 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17785 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17786 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17787 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17788 ;
    wire bfn_17_16_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17789 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17790 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17791 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17792 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17793 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17794 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n755 ;
    wire bfn_17_18_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17766 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n112 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17767 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n161 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17768 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n210 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17769 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n259 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17770 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17771 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17772 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17773 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363 ;
    wire bfn_17_19_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17774 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n504 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17775 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n553 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17776 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n602 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17777 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17778 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17779 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n751 ;
    wire n142_adj_2422_cascade_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756 ;
    wire Amp25_out1_14;
    wire n142_adj_2422;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727 ;
    wire n141_adj_2421_cascade_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18 ;
    wire Error_sub_temp_30_adj_2385;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n737 ;
    wire bfn_17_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n741 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18369 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n745 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18370 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n749 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18371 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n753 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18372 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n757 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18373 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n761 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18374 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n765 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18375 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18376 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n769 ;
    wire bfn_17_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n773 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18377 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n777 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18378 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n781 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18379 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n785 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18380 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n789 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18381 ;
    wire n793_adj_2424;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18382 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n795 ;
    wire bfn_18_5_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n84 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17266 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n133 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17267 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n182 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17268 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n231 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17269 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n280 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17270 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n329 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17271 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n378 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17272 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17273 ;
    wire bfn_18_6_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17274 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n427 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17275 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22 ;
    wire bfn_18_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17942 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17943 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17944 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17945 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17946 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17947 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17948 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17949 ;
    wire bfn_18_9_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17950 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n777 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17951 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n781 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17952 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n785 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17953 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n789 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17954 ;
    wire n793;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17955 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n795 ;
    wire bfn_18_10_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17882 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17883 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17884 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17885 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17886 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17887 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17888 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17889 ;
    wire bfn_18_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17890 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17891 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17892 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17893 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17894 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17895 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n779 ;
    wire bfn_18_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17867 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17868 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17869 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17870 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17871 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17872 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17873 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17874 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435 ;
    wire bfn_18_13_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17875 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17876 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n571 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17877 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n620 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17878 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n669 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17879 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n718 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17880 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n775 ;
    wire bfn_18_14_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17841 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17842 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17843 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17844 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17845 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17846 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17847 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17848 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465 ;
    wire bfn_18_15_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17849 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17850 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17851 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17852 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n666 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17853 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n715 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17854 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353 ;
    wire bfn_18_16_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n75 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17826 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17827 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17828 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17829 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17830 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17831 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17832 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17833 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500 ;
    wire bfn_18_17_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17834 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17835 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17836 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17837 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17838 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17839 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n767 ;
    wire bfn_18_18_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n60 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17751 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17752 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17753 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n207 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17754 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n256 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17755 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n305 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17756 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17757 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17758 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365 ;
    wire bfn_18_19_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17759 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n501 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17760 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n550 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17761 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n599 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17762 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17763 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n697 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17764 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n747 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20174 ;
    wire bfn_18_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15883 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15884 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15885 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15886 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15887 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15888 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15889 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15890 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8 ;
    wire bfn_18_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15891 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15892 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15893 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15894 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15895 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15896 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15897 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15898 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16 ;
    wire bfn_18_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15899 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15900 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15901 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15902 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15903 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15904 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15905 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15906 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24 ;
    wire bfn_18_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15907 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15908 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15909 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15910 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15911 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15912 ;
    wire bfn_18_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n93 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18354 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n142 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18355 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n191 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18356 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n240 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18357 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n289 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18358 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n338 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18359 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n387 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18360 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18361 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n436 ;
    wire bfn_18_27_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n485 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18362 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n534 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18363 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n583 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18364 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n632 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18365 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n681 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18366 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n730 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18367 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n791 ;
    wire bfn_19_5_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17641 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17642 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17643 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17644 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17645 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17646 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17647 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17648 ;
    wire bfn_19_6_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17649 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17650 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17651 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17652 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17653 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n769 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17654 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n771 ;
    wire bfn_19_7_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17626 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n124 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17627 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n173 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17628 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n222 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17629 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n271 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17630 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n320 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17631 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n369 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17632 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17633 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n418 ;
    wire bfn_19_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n467 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17634 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n516 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17635 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n565 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17636 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n614 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17637 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n663 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17638 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n765 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n712 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17639 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382 ;
    wire bfn_19_9_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n93 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17927 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17928 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n191 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17929 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n240 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17930 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n289 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17931 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n338 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17932 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n387 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17933 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17934 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n436 ;
    wire bfn_19_10_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n485 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17935 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n534 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17936 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n583 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17937 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n632 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17938 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n681 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17939 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n730 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17940 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416 ;
    wire bfn_19_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17912 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17913 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17914 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17915 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n286 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17916 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n335 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17917 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n384 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17918 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17919 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n433 ;
    wire bfn_19_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n482 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17920 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n531 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17921 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n580 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17922 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n629 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17923 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n678 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17924 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n727 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17925 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421 ;
    wire bfn_19_13_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n72 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17811 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n121 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17812 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n170 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17813 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n219 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17814 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17815 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17816 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17817 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17818 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n415 ;
    wire bfn_19_14_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17819 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17820 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17821 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17822 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17823 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n709 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17824 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n763 ;
    wire bfn_19_15_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n69 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n115 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17796 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n118 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n164 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17797 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n167 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n213 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17798 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n216 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17799 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n265 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17800 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n360 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17801 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n409 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17802 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17803 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n412 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n458 ;
    wire bfn_19_16_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n461 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n507 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17804 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n510 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17805 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17806 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17807 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17808 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17809 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354 ;
    wire bfn_19_17_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17711 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17712 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n746 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17713 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n750 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17714 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n754 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17715 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n758 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17716 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n762 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17717 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17718 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n766 ;
    wire bfn_19_18_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n770 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17719 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n774 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17720 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n778 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17721 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17722 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n786 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17723 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17724 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17725 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17726 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO ;
    wire bfn_19_19_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20870 ;
    wire \foc.preSatVoltage_10 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n738 ;
    wire bfn_19_21_0_;
    wire Error_sub_temp_31_adj_2384;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18144 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n8356 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18145 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18146 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18147 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18148 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18149 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18150 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18151 ;
    wire bfn_19_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18152 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18153 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18154 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18155 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18156 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n790 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18157 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n794 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18158 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18159 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n796 ;
    wire bfn_19_23_0_;
    wire bfn_19_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n60 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18189 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18190 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18191 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18192 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18193 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18194 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18195 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18196 ;
    wire bfn_19_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18197 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18198 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18199 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18200 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18201 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n746 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18202 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n747 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO ;
    wire bfn_19_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n90 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18339 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n139 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18340 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n188 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18341 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n237 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18342 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n286 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18343 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n335 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18344 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n384 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18345 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18346 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n433 ;
    wire bfn_19_27_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n482 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18347 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n531 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18348 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n580 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18349 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n629 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18350 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n678 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18351 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n727 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n786 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18352 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n787 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO ;
    wire bfn_19_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n87 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18324 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n136 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18325 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n185 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18326 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n234 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18327 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n283 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18328 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n332 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18329 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n381 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18330 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18331 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n430 ;
    wire bfn_19_29_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n479 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18332 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n528 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18333 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n577 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18334 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n626 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18335 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n675 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18336 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n724 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n782 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18337 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n783 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n78 ;
    wire bfn_20_5_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n81 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n127 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18122 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n130 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n176 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18123 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n179 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n225 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18124 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n228 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n274 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18125 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n277 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n323 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18126 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n326 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n372 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18127 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n375 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n421 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18128 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18129 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n424 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n470 ;
    wire bfn_20_6_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n473 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n519 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18130 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n568 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18131 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n617 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18132 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n773 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n522 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n18133 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357 ;
    wire bfn_20_7_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17611 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17612 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17613 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17614 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n268 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17615 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n317 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17616 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n366 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17617 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17618 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449 ;
    wire bfn_20_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n464 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17619 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n513 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17620 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n562 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17621 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n611 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17622 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n660 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17623 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n761 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17624 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386 ;
    wire bfn_20_9_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17581 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17582 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17583 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17584 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17585 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17586 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17587 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17588 ;
    wire bfn_20_10_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17589 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17590 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17591 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17592 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17593 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n753 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17594 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404 ;
    wire bfn_20_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n87 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17897 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n136 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17898 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n185 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17899 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n234 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17900 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17901 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17902 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n381 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17903 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17904 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n430 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n476 ;
    wire bfn_20_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n479 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n525 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17905 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n528 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n574 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17906 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n577 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n623 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17907 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n626 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n672 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17908 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n675 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n721 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17909 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n724 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n782 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17910 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n783 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO ;
    wire Error_sub_temp_30;
    wire bfn_20_14_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17505 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17506 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17507 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17508 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17509 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17510 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17511 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17512 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO ;
    wire bfn_20_15_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17513 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17514 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17515 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17516 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17517 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n790 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17518 ;
    wire n794_adj_2420;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n791 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17519 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17520 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n796 ;
    wire bfn_20_16_0_;
    wire \foc.preSatVoltage_19 ;
    wire \foc.qVoltage_10 ;
    wire \foc.preSatVoltage_22 ;
    wire \foc.qVoltage_13 ;
    wire \foc.qVoltage_3 ;
    wire \foc.preSatVoltage_13 ;
    wire \foc.qVoltage_4_cascade_ ;
    wire \foc.preSatVoltage_12 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17 ;
    wire \foc.qVoltage_8_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n8265 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19884 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n27 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20590 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20614 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_ ;
    wire \foc.qVoltage_7 ;
    wire Error_sub_temp_31;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_ ;
    wire Saturate_out1_31__N_266_adj_2417_cascade_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20620 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20608 ;
    wire Saturate_out1_31__N_267_adj_2418_cascade_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20676 ;
    wire bfn_20_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n63 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n109 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18204 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n158 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18205 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n207 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18206 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n256 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18207 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n305 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18208 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n354 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18209 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n403 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18210 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18211 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n452 ;
    wire bfn_20_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n501 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18212 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n550 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18213 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n599 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18214 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n648 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18215 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n697 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18216 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n750 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18217 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n751 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO ;
    wire bfn_20_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n66 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n112 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18219 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n161 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18220 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n210 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18221 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n259 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18222 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n308 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18223 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n357 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18224 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n406 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18225 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18226 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n455 ;
    wire bfn_20_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n504 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18227 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n553 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18228 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n602 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18229 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n651 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18230 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n700 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18231 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n754 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18232 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n755 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO ;
    wire bfn_20_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n84 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18309 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n133 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18310 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n182 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18311 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n231 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18312 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n280 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18313 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n329 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18314 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n378 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18315 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18316 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n427 ;
    wire bfn_20_29_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n476 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18317 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n525 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18318 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n574 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18319 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n623 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18320 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n672 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18321 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n721 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n778 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18322 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n779 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n66 ;
    wire bfn_21_7_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17596 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17597 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17598 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n262 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17599 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n311 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17600 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n314 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17601 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n363 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17602 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17603 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468 ;
    wire bfn_21_8_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17604 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n556 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17605 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n559 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n605 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17606 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n608 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n654 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17607 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n657 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n703 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17608 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n757 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n706 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17609 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n759 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO ;
    wire bfn_21_9_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n63 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17566 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17567 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17568 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17569 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17570 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n308 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17571 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n357 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17572 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17573 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n406 ;
    wire bfn_21_10_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n455 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17574 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17575 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17576 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17577 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n651 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17578 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n749 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n700 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17579 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO ;
    wire bfn_21_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17551 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n109 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17552 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n158 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17553 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17554 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17555 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17556 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n354 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17557 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17558 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n403 ;
    wire bfn_21_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n452 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17559 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17560 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17561 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17562 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n648 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17563 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n745 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17564 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO ;
    wire \foc.dVoltage_2_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_ ;
    wire \foc.dVoltage_15 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_ ;
    wire \foc.dVoltage_10 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_ ;
    wire \foc.qVoltage_5_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20604 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20588 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896 ;
    wire \foc.Out_31__N_333_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31 ;
    wire \foc.Out_31__N_332_cascade_ ;
    wire \foc.qVoltage_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18 ;
    wire \foc.qVoltage_14_cascade_ ;
    wire \foc.preSatVoltage_23 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24 ;
    wire \foc.qVoltage_15 ;
    wire bfn_21_17_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n57 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17736 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n108 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n106 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17737 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n111 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17738 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n114 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17739 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n253 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n117 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17740 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n120 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17741 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n351 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n123 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17742 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17743 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n126 ;
    wire bfn_21_18_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n129 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17744 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n132 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17745 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n135 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17746 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n138 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17747 ;
    wire n141;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n691 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17748 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427 ;
    wire n146;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n742 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17749 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n743 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO ;
    wire Saturate_out1_31__N_266_adj_2417;
    wire Saturate_out1_31__N_267_adj_2418;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19308 ;
    wire bfn_21_21_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n57 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18174 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n106 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18175 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n155 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18176 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n204 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18177 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n253 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18178 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n302 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18179 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n351 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18180 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18181 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n400 ;
    wire bfn_21_22_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n449 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18182 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n498 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18183 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n547 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18184 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n596 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18185 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n645 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n691 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18186 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n694 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n742 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18187 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n743 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4 ;
    wire bfn_21_23_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15913 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15914 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15915 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15916 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15917 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15918 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15919 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15920 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12 ;
    wire bfn_21_24_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15921 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15922 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15923 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15924 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15925 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15926 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15927 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15928 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20 ;
    wire bfn_21_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21 ;
    wire Add_add_temp_21_adj_2399;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15929 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22 ;
    wire Add_add_temp_22_adj_2398;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15930 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23 ;
    wire Add_add_temp_23_adj_2397;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15931 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24 ;
    wire Add_add_temp_24_adj_2396;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15932 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25 ;
    wire Add_add_temp_25_adj_2395;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15933 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26 ;
    wire Add_add_temp_26_adj_2394;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15934 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27 ;
    wire Add_add_temp_27_adj_2393;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15935 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15936 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28 ;
    wire Add_add_temp_28_adj_2392;
    wire bfn_21_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29 ;
    wire Add_add_temp_29_adj_2391;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15937 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30 ;
    wire Add_add_temp_30_adj_2390;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15938 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27 ;
    wire Add_add_temp_31_adj_2389;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15939 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28 ;
    wire Add_add_temp_32_adj_2388;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15940 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29 ;
    wire Add_add_temp_33_adj_2387;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15941 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30 ;
    wire Add_add_temp_34_adj_2386;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15942 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15943 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31 ;
    wire bfn_21_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n81 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18294 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n130 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18295 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n179 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18296 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n228 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18297 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n277 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18298 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18299 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18300 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18301 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586 ;
    wire bfn_21_29_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18302 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18303 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n571 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18304 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n620 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18305 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n669 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18306 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n718 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18307 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n105 ;
    wire bfn_22_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17536 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17537 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n155 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17538 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n204 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17539 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17540 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n302 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17541 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17542 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17543 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n400 ;
    wire bfn_22_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n449 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17544 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n498 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17545 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n547 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17546 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n596 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17547 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n645 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17548 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n694 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n741 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17549 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20556 ;
    wire \foc.dVoltage_5_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20554 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_ ;
    wire \foc.dVoltage_12 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20560 ;
    wire \foc.Out_31__N_332_adj_2312_cascade_ ;
    wire \foc.dVoltage_8 ;
    wire \foc.Out_31__N_333_adj_2310_cascade_ ;
    wire \foc.dVoltage_14 ;
    wire \foc.dVoltage_3_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20572 ;
    wire \foc.dVoltage_11_cascade_ ;
    wire \foc.dVoltage_9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20566 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11 ;
    wire \foc.qVoltage_2_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20594 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20612 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20618 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15 ;
    wire \foc.qVoltage_6 ;
    wire \foc.Out_31__N_332 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21 ;
    wire \foc.Out_31__N_333 ;
    wire \foc.qVoltage_12 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_ ;
    wire Saturate_out1_31__N_267_cascade_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20634 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4 ;
    wire bfn_22_19_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15973 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15974 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15975 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15976 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15977 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15978 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15979 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15980 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12 ;
    wire bfn_22_20_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15981 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15982 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15983 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15984 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15985 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15986 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15987 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15988 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20 ;
    wire bfn_22_21_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15989 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15990 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15991 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24 ;
    wire Add_add_temp_24;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15992 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15993 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15994 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15995 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15996 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28 ;
    wire Add_add_temp_28;
    wire bfn_22_22_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29 ;
    wire Add_add_temp_29;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15997 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15998 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15999 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n16000 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n16001 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n16002 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n16003 ;
    wire Add_add_temp_14_adj_2406;
    wire Add_add_temp_12_adj_2408;
    wire Add_add_temp_13_adj_2407;
    wire Add_add_temp_16_adj_2404;
    wire Add_add_temp_17_adj_2403;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_ ;
    wire Add_add_temp_15_adj_2405;
    wire Add_add_temp_20_adj_2400;
    wire Add_add_temp_19_adj_2401;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_ ;
    wire Add_add_temp_18_adj_2402;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19733 ;
    wire Add_add_temp_5_adj_2415;
    wire Add_add_temp_4_adj_2416;
    wire Add_add_temp_8_adj_2412;
    wire Add_add_temp_7_adj_2413;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_ ;
    wire Add_add_temp_6_adj_2414;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20704 ;
    wire bfn_22_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n69 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n115 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18234 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n164 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18235 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n213 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18236 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n262 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18237 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n311 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18238 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n360 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18239 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n409 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18240 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18241 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n458 ;
    wire bfn_22_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n507 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18242 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n556 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18243 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n605 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18244 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n654 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18245 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n703 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18246 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n758 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18247 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n759 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO ;
    wire bfn_22_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n78 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18279 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n127 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18280 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n176 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18281 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n225 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18282 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n274 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18283 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n323 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18284 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18285 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18286 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595 ;
    wire bfn_22_29_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18287 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18288 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18289 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18290 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n666 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18291 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n715 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n770 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18292 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n771 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n102 ;
    wire bfn_23_11_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n54 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17521 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n103 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17522 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n152 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17523 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n201 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17524 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n250 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17525 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n299 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17526 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n348 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17527 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17528 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n397 ;
    wire bfn_23_12_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n446 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17529 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n495 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17530 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n544 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17531 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n593 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17532 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n642 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17533 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n737 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n738 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n17534 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n739 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20546 ;
    wire \foc.dVoltage_13_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20576 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n14 ;
    wire \foc.dVoltage_6 ;
    wire \foc.Out_31__N_332_adj_2312 ;
    wire \foc.Out_31__N_333_adj_2310 ;
    wire \foc.dVoltage_7 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19858 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_ ;
    wire Add_add_temp_31;
    wire Add_add_temp_32;
    wire Add_add_temp_30;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20644 ;
    wire Add_add_temp_34;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_ ;
    wire Add_add_temp_33;
    wire Saturate_out1_31__N_266_cascade_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4 ;
    wire Add_add_temp_26;
    wire Add_add_temp_27;
    wire Add_add_temp_25;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5 ;
    wire Saturate_out1_31__N_267;
    wire Saturate_out1_31__N_266;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20688 ;
    wire Add_add_temp_17;
    wire Add_add_temp_16;
    wire Add_add_temp_15;
    wire Add_add_temp_5;
    wire Add_add_temp_4;
    wire Add_add_temp_8;
    wire Add_add_temp_7;
    wire Add_add_temp_6;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20712 ;
    wire Add_add_temp_9;
    wire Add_add_temp_11;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_ ;
    wire Add_add_temp_10;
    wire Add_add_temp_14;
    wire Add_add_temp_13;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_ ;
    wire Add_add_temp_12;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15205 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20670 ;
    wire Add_add_temp_20;
    wire Add_add_temp_18;
    wire Add_add_temp_19;
    wire Add_add_temp_21;
    wire Add_add_temp_23;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_ ;
    wire Add_add_temp_22;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20656 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31 ;
    wire pin3_clk_16mhz_N;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n19755 ;
    wire Add_add_temp_11_adj_2409;
    wire Add_add_temp_9_adj_2411;
    wire Add_add_temp_10_adj_2410;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n20718 ;
    wire bfn_23_25_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n72 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n118 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18249 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n167 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18250 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n216 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18251 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n265 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18252 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n314 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18253 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n363 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18254 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n412 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18255 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18256 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n461 ;
    wire bfn_23_26_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n510 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18257 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n559 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18258 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n608 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18259 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n657 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18260 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n706 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18261 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n762 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18262 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n763 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n102 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ;
    wire bfn_23_27_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n75 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n105 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n121 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18264 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n124 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n170 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18265 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n173 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n219 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18266 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n222 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n268 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18267 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n271 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n317 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18268 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n120 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n320 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n366 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18269 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n369 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n415 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18270 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18271 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n126 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n418 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n464 ;
    wire bfn_23_28_0_;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n467 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n513 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18272 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n516 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n562 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18273 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n565 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n135 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n611 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18274 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n614 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n660 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18275 ;
    wire n141_adj_2421;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n663 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n709 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18276 ;
    wire n146_adj_2423;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n712 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n766 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n18277 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n767 ;
    wire \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_ ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0 ;
    wire bfn_24_16_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20184 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15568 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20186 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15569 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20188 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15570 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20190 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15571 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20192 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15572 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15573 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20194 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14 ;
    wire bfn_24_17_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20196 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n20198 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15574 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15575 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17 ;
    wire \foc.preSatVoltage_10_adj_2311 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15576 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15577 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11 ;
    wire \foc.preSatVoltage_12_adj_2330 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15578 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15579 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15580 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14 ;
    wire bfn_24_18_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15581 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15582 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15583 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15584 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26 ;
    wire \foc.preSatVoltage_19_adj_2329 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15585 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15586 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15587 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15588 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22 ;
    wire bfn_24_19_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22 ;
    wire \foc.preSatVoltage_23_adj_2328 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15589 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15590 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15591 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15592 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15593 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15594 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15595 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15596 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30 ;
    wire bfn_24_20_0_;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.n15597 ;
    wire \foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31 ;
    wire _gnd_net_;

    defparam pin10_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin10_pad_iopad.PULLUP=1'b0;
    IO_PAD pin10_pad_iopad (
            .OE(N__69497),
            .DIN(N__69496),
            .DOUT(N__69495),
            .PACKAGEPIN(pin10));
    defparam pin10_pad_preio.PIN_TYPE=6'b101001;
    defparam pin10_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin10_pad_preio (
            .PADOEN(N__69497),
            .PADOUT(N__69496),
            .PADIN(N__69495),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin11_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin11_pad_iopad.PULLUP=1'b0;
    IO_PAD pin11_pad_iopad (
            .OE(N__69488),
            .DIN(N__69487),
            .DOUT(N__69486),
            .PACKAGEPIN(pin11));
    defparam pin11_pad_preio.PIN_TYPE=6'b101001;
    defparam pin11_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin11_pad_preio (
            .PADOEN(N__69488),
            .PADOUT(N__69487),
            .PADIN(N__69486),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin12_pad_iopad.PULLUP=1'b0;
    IO_PAD pin12_pad_iopad (
            .OE(N__69479),
            .DIN(N__69478),
            .DOUT(N__69477),
            .PACKAGEPIN(pin12));
    defparam pin12_pad_preio.PIN_TYPE=6'b101001;
    defparam pin12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin12_pad_preio (
            .PADOEN(N__69479),
            .PADOUT(N__69478),
            .PADIN(N__69477),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin13_pad_iopad.PULLUP=1'b0;
    IO_PAD pin13_pad_iopad (
            .OE(N__69470),
            .DIN(N__69469),
            .DOUT(N__69468),
            .PACKAGEPIN(pin13));
    defparam pin13_pad_preio.PIN_TYPE=6'b101001;
    defparam pin13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin13_pad_preio (
            .PADOEN(N__69470),
            .PADOUT(N__69469),
            .PADIN(N__69468),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin14_sdo_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin14_sdo_pad_iopad.PULLUP=1'b0;
    IO_PAD pin14_sdo_pad_iopad (
            .OE(N__69461),
            .DIN(N__69460),
            .DOUT(N__69459),
            .PACKAGEPIN(pin14_sdo));
    defparam pin14_sdo_pad_preio.PIN_TYPE=6'b101001;
    defparam pin14_sdo_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin14_sdo_pad_preio (
            .PADOEN(N__69461),
            .PADOUT(N__69460),
            .PADIN(N__69459),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin15_sdi_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin15_sdi_pad_iopad.PULLUP=1'b0;
    IO_PAD pin15_sdi_pad_iopad (
            .OE(N__69452),
            .DIN(N__69451),
            .DOUT(N__69450),
            .PACKAGEPIN(pin15_sdi));
    defparam pin15_sdi_pad_preio.PIN_TYPE=6'b101001;
    defparam pin15_sdi_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin15_sdi_pad_preio (
            .PADOEN(N__69452),
            .PADOUT(N__69451),
            .PADIN(N__69450),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin16_sck_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin16_sck_pad_iopad.PULLUP=1'b0;
    IO_PAD pin16_sck_pad_iopad (
            .OE(N__69443),
            .DIN(N__69442),
            .DOUT(N__69441),
            .PACKAGEPIN(pin16_sck));
    defparam pin16_sck_pad_preio.PIN_TYPE=6'b101001;
    defparam pin16_sck_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin16_sck_pad_preio (
            .PADOEN(N__69443),
            .PADOUT(N__69442),
            .PADIN(N__69441),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin17_ss_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin17_ss_pad_iopad.PULLUP=1'b0;
    IO_PAD pin17_ss_pad_iopad (
            .OE(N__69434),
            .DIN(N__69433),
            .DOUT(N__69432),
            .PACKAGEPIN(pin17_ss));
    defparam pin17_ss_pad_preio.PIN_TYPE=6'b101001;
    defparam pin17_ss_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin17_ss_pad_preio (
            .PADOEN(N__69434),
            .PADOUT(N__69433),
            .PADIN(N__69432),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin18_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin18_pad_iopad.PULLUP=1'b0;
    IO_PAD pin18_pad_iopad (
            .OE(N__69425),
            .DIN(N__69424),
            .DOUT(N__69423),
            .PACKAGEPIN(pin18));
    defparam pin18_pad_preio.PIN_TYPE=6'b101001;
    defparam pin18_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin18_pad_preio (
            .PADOEN(N__69425),
            .PADOUT(N__69424),
            .PADIN(N__69423),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin19_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin19_pad_iopad.PULLUP=1'b0;
    IO_PAD pin19_pad_iopad (
            .OE(N__69416),
            .DIN(N__69415),
            .DOUT(N__69414),
            .PACKAGEPIN(pin19));
    defparam pin19_pad_preio.PIN_TYPE=6'b101001;
    defparam pin19_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin19_pad_preio (
            .PADOEN(N__69416),
            .PADOUT(N__69415),
            .PADIN(N__69414),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin1_usb_dp_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin1_usb_dp_pad_iopad.PULLUP=1'b0;
    IO_PAD pin1_usb_dp_pad_iopad (
            .OE(N__69407),
            .DIN(N__69406),
            .DOUT(N__69405),
            .PACKAGEPIN(pin1_usb_dp));
    defparam pin1_usb_dp_pad_preio.PIN_TYPE=6'b101001;
    defparam pin1_usb_dp_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin1_usb_dp_pad_preio (
            .PADOEN(N__69407),
            .PADOUT(N__69406),
            .PADIN(N__69405),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin20_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin20_pad_iopad.PULLUP=1'b0;
    IO_PAD pin20_pad_iopad (
            .OE(N__69398),
            .DIN(N__69397),
            .DOUT(N__69396),
            .PACKAGEPIN(pin20));
    defparam pin20_pad_preio.PIN_TYPE=6'b101001;
    defparam pin20_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin20_pad_preio (
            .PADOEN(N__69398),
            .PADOUT(N__69397),
            .PADIN(N__69396),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin21_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin21_pad_iopad.PULLUP=1'b0;
    IO_PAD pin21_pad_iopad (
            .OE(N__69389),
            .DIN(N__69388),
            .DOUT(N__69387),
            .PACKAGEPIN(pin21));
    defparam pin21_pad_preio.PIN_TYPE=6'b101001;
    defparam pin21_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin21_pad_preio (
            .PADOEN(N__69389),
            .PADOUT(N__69388),
            .PADIN(N__69387),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin22_pad_iopad.PULLUP=1'b0;
    IO_PAD pin22_pad_iopad (
            .OE(N__69380),
            .DIN(N__69379),
            .DOUT(N__69378),
            .PACKAGEPIN(pin22));
    defparam pin22_pad_preio.PIN_TYPE=6'b101001;
    defparam pin22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin22_pad_preio (
            .PADOEN(N__69380),
            .PADOUT(N__69379),
            .PADIN(N__69378),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin23_pad_iopad.PULLUP=1'b0;
    IO_PAD pin23_pad_iopad (
            .OE(N__69371),
            .DIN(N__69370),
            .DOUT(N__69369),
            .PACKAGEPIN(pin23));
    defparam pin23_pad_preio.PIN_TYPE=6'b101001;
    defparam pin23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin23_pad_preio (
            .PADOEN(N__69371),
            .PADOUT(N__69370),
            .PADIN(N__69369),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin24_pad_iopad.PULLUP=1'b0;
    IO_PAD pin24_pad_iopad (
            .OE(N__69362),
            .DIN(N__69361),
            .DOUT(N__69360),
            .PACKAGEPIN(pin24));
    defparam pin24_pad_preio.PIN_TYPE=6'b101001;
    defparam pin24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin24_pad_preio (
            .PADOEN(N__69362),
            .PADOUT(N__69361),
            .PADIN(N__69360),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin2_usb_dn_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin2_usb_dn_pad_iopad.PULLUP=1'b0;
    IO_PAD pin2_usb_dn_pad_iopad (
            .OE(N__69353),
            .DIN(N__69352),
            .DOUT(N__69351),
            .PACKAGEPIN(pin2_usb_dn));
    defparam pin2_usb_dn_pad_preio.PIN_TYPE=6'b101001;
    defparam pin2_usb_dn_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin2_usb_dn_pad_preio (
            .PADOEN(N__69353),
            .PADOUT(N__69352),
            .PADIN(N__69351),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin7_pad_iopad.PULLUP=1'b0;
    IO_PAD pin7_pad_iopad (
            .OE(N__69344),
            .DIN(N__69343),
            .DOUT(N__69342),
            .PACKAGEPIN(pin7));
    defparam pin7_pad_preio.PIN_TYPE=6'b101001;
    defparam pin7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin7_pad_preio (
            .PADOEN(N__69344),
            .PADOUT(N__69343),
            .PADIN(N__69342),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin8_pad_iopad.PULLUP=1'b0;
    IO_PAD pin8_pad_iopad (
            .OE(N__69335),
            .DIN(N__69334),
            .DOUT(N__69333),
            .PACKAGEPIN(pin8));
    defparam pin8_pad_preio.PIN_TYPE=6'b101001;
    defparam pin8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin8_pad_preio (
            .PADOEN(N__69335),
            .PADOUT(N__69334),
            .PADIN(N__69333),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin9_pad_iopad.PULLUP=1'b0;
    IO_PAD pin9_pad_iopad (
            .OE(N__69326),
            .DIN(N__69325),
            .DOUT(N__69324),
            .PACKAGEPIN(pin9));
    defparam pin9_pad_preio.PIN_TYPE=6'b101001;
    defparam pin9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin9_pad_preio (
            .PADOEN(N__69326),
            .PADOUT(N__69325),
            .PADIN(N__69324),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin3_clk_16mhz_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin3_clk_16mhz_pad_iopad.PULLUP=1'b0;
    IO_PAD pin3_clk_16mhz_pad_iopad (
            .OE(N__69317),
            .DIN(N__69316),
            .DOUT(N__69315),
            .PACKAGEPIN(pin3_clk_16mhz));
    defparam pin3_clk_16mhz_pad_preio.PIN_TYPE=6'b000001;
    defparam pin3_clk_16mhz_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin3_clk_16mhz_pad_preio (
            .PADOEN(N__69317),
            .PADOUT(N__69316),
            .PADIN(N__69315),
            .CLOCKENABLE(),
            .DIN0(pin3_clk_16mhz_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__15992 (
            .O(N__69298),
            .I(N__69295));
    InMux I__15991 (
            .O(N__69295),
            .I(N__69288));
    InMux I__15990 (
            .O(N__69294),
            .I(N__69288));
    InMux I__15989 (
            .O(N__69293),
            .I(N__69285));
    LocalMux I__15988 (
            .O(N__69288),
            .I(N__69282));
    LocalMux I__15987 (
            .O(N__69285),
            .I(N__69279));
    Sp12to4 I__15986 (
            .O(N__69282),
            .I(N__69276));
    Span4Mux_h I__15985 (
            .O(N__69279),
            .I(N__69273));
    Odrv12 I__15984 (
            .O(N__69276),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26 ));
    Odrv4 I__15983 (
            .O(N__69273),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26 ));
    InMux I__15982 (
            .O(N__69268),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15592 ));
    InMux I__15981 (
            .O(N__69265),
            .I(N__69262));
    LocalMux I__15980 (
            .O(N__69262),
            .I(N__69259));
    Span12Mux_v I__15979 (
            .O(N__69259),
            .I(N__69256));
    Odrv12 I__15978 (
            .O(N__69256),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26 ));
    InMux I__15977 (
            .O(N__69253),
            .I(N__69246));
    InMux I__15976 (
            .O(N__69252),
            .I(N__69246));
    InMux I__15975 (
            .O(N__69251),
            .I(N__69243));
    LocalMux I__15974 (
            .O(N__69246),
            .I(N__69240));
    LocalMux I__15973 (
            .O(N__69243),
            .I(N__69237));
    Span12Mux_v I__15972 (
            .O(N__69240),
            .I(N__69234));
    Span4Mux_h I__15971 (
            .O(N__69237),
            .I(N__69231));
    Odrv12 I__15970 (
            .O(N__69234),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27 ));
    Odrv4 I__15969 (
            .O(N__69231),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27 ));
    InMux I__15968 (
            .O(N__69226),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15593 ));
    CascadeMux I__15967 (
            .O(N__69223),
            .I(N__69220));
    InMux I__15966 (
            .O(N__69220),
            .I(N__69217));
    LocalMux I__15965 (
            .O(N__69217),
            .I(N__69214));
    Span4Mux_v I__15964 (
            .O(N__69214),
            .I(N__69211));
    Odrv4 I__15963 (
            .O(N__69211),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27 ));
    InMux I__15962 (
            .O(N__69208),
            .I(N__69205));
    LocalMux I__15961 (
            .O(N__69205),
            .I(N__69200));
    InMux I__15960 (
            .O(N__69204),
            .I(N__69197));
    InMux I__15959 (
            .O(N__69203),
            .I(N__69194));
    Span4Mux_v I__15958 (
            .O(N__69200),
            .I(N__69191));
    LocalMux I__15957 (
            .O(N__69197),
            .I(N__69186));
    LocalMux I__15956 (
            .O(N__69194),
            .I(N__69186));
    Span4Mux_h I__15955 (
            .O(N__69191),
            .I(N__69183));
    Span4Mux_v I__15954 (
            .O(N__69186),
            .I(N__69180));
    Odrv4 I__15953 (
            .O(N__69183),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28 ));
    Odrv4 I__15952 (
            .O(N__69180),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28 ));
    InMux I__15951 (
            .O(N__69175),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15594 ));
    InMux I__15950 (
            .O(N__69172),
            .I(N__69169));
    LocalMux I__15949 (
            .O(N__69169),
            .I(N__69166));
    Span4Mux_v I__15948 (
            .O(N__69166),
            .I(N__69163));
    Span4Mux_h I__15947 (
            .O(N__69163),
            .I(N__69160));
    Odrv4 I__15946 (
            .O(N__69160),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28 ));
    InMux I__15945 (
            .O(N__69157),
            .I(N__69150));
    InMux I__15944 (
            .O(N__69156),
            .I(N__69150));
    CascadeMux I__15943 (
            .O(N__69155),
            .I(N__69147));
    LocalMux I__15942 (
            .O(N__69150),
            .I(N__69144));
    InMux I__15941 (
            .O(N__69147),
            .I(N__69141));
    Span4Mux_h I__15940 (
            .O(N__69144),
            .I(N__69136));
    LocalMux I__15939 (
            .O(N__69141),
            .I(N__69136));
    Sp12to4 I__15938 (
            .O(N__69136),
            .I(N__69133));
    Odrv12 I__15937 (
            .O(N__69133),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29 ));
    InMux I__15936 (
            .O(N__69130),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15595 ));
    CascadeMux I__15935 (
            .O(N__69127),
            .I(N__69124));
    InMux I__15934 (
            .O(N__69124),
            .I(N__69121));
    LocalMux I__15933 (
            .O(N__69121),
            .I(N__69118));
    Span4Mux_h I__15932 (
            .O(N__69118),
            .I(N__69115));
    Span4Mux_v I__15931 (
            .O(N__69115),
            .I(N__69112));
    Odrv4 I__15930 (
            .O(N__69112),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29 ));
    InMux I__15929 (
            .O(N__69109),
            .I(N__69102));
    InMux I__15928 (
            .O(N__69108),
            .I(N__69102));
    InMux I__15927 (
            .O(N__69107),
            .I(N__69099));
    LocalMux I__15926 (
            .O(N__69102),
            .I(N__69096));
    LocalMux I__15925 (
            .O(N__69099),
            .I(N__69093));
    Span4Mux_h I__15924 (
            .O(N__69096),
            .I(N__69090));
    Span4Mux_h I__15923 (
            .O(N__69093),
            .I(N__69087));
    Span4Mux_v I__15922 (
            .O(N__69090),
            .I(N__69084));
    Span4Mux_v I__15921 (
            .O(N__69087),
            .I(N__69081));
    Odrv4 I__15920 (
            .O(N__69084),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30 ));
    Odrv4 I__15919 (
            .O(N__69081),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30 ));
    InMux I__15918 (
            .O(N__69076),
            .I(bfn_24_20_0_));
    CascadeMux I__15917 (
            .O(N__69073),
            .I(N__69068));
    CascadeMux I__15916 (
            .O(N__69072),
            .I(N__69064));
    CascadeMux I__15915 (
            .O(N__69071),
            .I(N__69060));
    InMux I__15914 (
            .O(N__69068),
            .I(N__69046));
    InMux I__15913 (
            .O(N__69067),
            .I(N__69046));
    InMux I__15912 (
            .O(N__69064),
            .I(N__69046));
    InMux I__15911 (
            .O(N__69063),
            .I(N__69046));
    InMux I__15910 (
            .O(N__69060),
            .I(N__69046));
    InMux I__15909 (
            .O(N__69059),
            .I(N__69046));
    LocalMux I__15908 (
            .O(N__69046),
            .I(N__69040));
    InMux I__15907 (
            .O(N__69045),
            .I(N__69037));
    InMux I__15906 (
            .O(N__69044),
            .I(N__69032));
    InMux I__15905 (
            .O(N__69043),
            .I(N__69032));
    Odrv4 I__15904 (
            .O(N__69040),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31 ));
    LocalMux I__15903 (
            .O(N__69037),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31 ));
    LocalMux I__15902 (
            .O(N__69032),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31 ));
    InMux I__15901 (
            .O(N__69025),
            .I(N__69022));
    LocalMux I__15900 (
            .O(N__69022),
            .I(N__69019));
    Span4Mux_v I__15899 (
            .O(N__69019),
            .I(N__69016));
    Odrv4 I__15898 (
            .O(N__69016),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30 ));
    InMux I__15897 (
            .O(N__69013),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15597 ));
    CascadeMux I__15896 (
            .O(N__69010),
            .I(N__69007));
    InMux I__15895 (
            .O(N__69007),
            .I(N__69003));
    CascadeMux I__15894 (
            .O(N__69006),
            .I(N__69000));
    LocalMux I__15893 (
            .O(N__69003),
            .I(N__68997));
    InMux I__15892 (
            .O(N__69000),
            .I(N__68994));
    Span4Mux_v I__15891 (
            .O(N__68997),
            .I(N__68991));
    LocalMux I__15890 (
            .O(N__68994),
            .I(N__68988));
    Span4Mux_h I__15889 (
            .O(N__68991),
            .I(N__68983));
    Span4Mux_v I__15888 (
            .O(N__68988),
            .I(N__68983));
    Span4Mux_v I__15887 (
            .O(N__68983),
            .I(N__68980));
    Odrv4 I__15886 (
            .O(N__68980),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31 ));
    InMux I__15885 (
            .O(N__68977),
            .I(N__68974));
    LocalMux I__15884 (
            .O(N__68974),
            .I(N__68971));
    Span4Mux_v I__15883 (
            .O(N__68971),
            .I(N__68968));
    Odrv4 I__15882 (
            .O(N__68968),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18 ));
    InMux I__15881 (
            .O(N__68965),
            .I(N__68962));
    LocalMux I__15880 (
            .O(N__68962),
            .I(N__68958));
    CascadeMux I__15879 (
            .O(N__68961),
            .I(N__68955));
    Sp12to4 I__15878 (
            .O(N__68958),
            .I(N__68952));
    InMux I__15877 (
            .O(N__68955),
            .I(N__68949));
    Odrv12 I__15876 (
            .O(N__68952),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26 ));
    LocalMux I__15875 (
            .O(N__68949),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26 ));
    InMux I__15874 (
            .O(N__68944),
            .I(N__68937));
    InMux I__15873 (
            .O(N__68943),
            .I(N__68937));
    InMux I__15872 (
            .O(N__68942),
            .I(N__68933));
    LocalMux I__15871 (
            .O(N__68937),
            .I(N__68930));
    InMux I__15870 (
            .O(N__68936),
            .I(N__68927));
    LocalMux I__15869 (
            .O(N__68933),
            .I(N__68924));
    Span4Mux_h I__15868 (
            .O(N__68930),
            .I(N__68919));
    LocalMux I__15867 (
            .O(N__68927),
            .I(N__68919));
    Odrv12 I__15866 (
            .O(N__68924),
            .I(\foc.preSatVoltage_19_adj_2329 ));
    Odrv4 I__15865 (
            .O(N__68919),
            .I(\foc.preSatVoltage_19_adj_2329 ));
    InMux I__15864 (
            .O(N__68914),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15585 ));
    InMux I__15863 (
            .O(N__68911),
            .I(N__68907));
    InMux I__15862 (
            .O(N__68910),
            .I(N__68904));
    LocalMux I__15861 (
            .O(N__68907),
            .I(N__68901));
    LocalMux I__15860 (
            .O(N__68904),
            .I(N__68898));
    Span4Mux_v I__15859 (
            .O(N__68901),
            .I(N__68895));
    Odrv12 I__15858 (
            .O(N__68898),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27 ));
    Odrv4 I__15857 (
            .O(N__68895),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27 ));
    CascadeMux I__15856 (
            .O(N__68890),
            .I(N__68887));
    InMux I__15855 (
            .O(N__68887),
            .I(N__68884));
    LocalMux I__15854 (
            .O(N__68884),
            .I(N__68881));
    Span4Mux_v I__15853 (
            .O(N__68881),
            .I(N__68878));
    Span4Mux_h I__15852 (
            .O(N__68878),
            .I(N__68875));
    Odrv4 I__15851 (
            .O(N__68875),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19 ));
    InMux I__15850 (
            .O(N__68872),
            .I(N__68866));
    InMux I__15849 (
            .O(N__68871),
            .I(N__68866));
    LocalMux I__15848 (
            .O(N__68866),
            .I(N__68863));
    Span4Mux_h I__15847 (
            .O(N__68863),
            .I(N__68858));
    InMux I__15846 (
            .O(N__68862),
            .I(N__68855));
    InMux I__15845 (
            .O(N__68861),
            .I(N__68852));
    Sp12to4 I__15844 (
            .O(N__68858),
            .I(N__68845));
    LocalMux I__15843 (
            .O(N__68855),
            .I(N__68845));
    LocalMux I__15842 (
            .O(N__68852),
            .I(N__68845));
    Odrv12 I__15841 (
            .O(N__68845),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20 ));
    InMux I__15840 (
            .O(N__68842),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15586 ));
    CascadeMux I__15839 (
            .O(N__68839),
            .I(N__68836));
    InMux I__15838 (
            .O(N__68836),
            .I(N__68833));
    LocalMux I__15837 (
            .O(N__68833),
            .I(N__68830));
    Span4Mux_v I__15836 (
            .O(N__68830),
            .I(N__68826));
    InMux I__15835 (
            .O(N__68829),
            .I(N__68823));
    Odrv4 I__15834 (
            .O(N__68826),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28 ));
    LocalMux I__15833 (
            .O(N__68823),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28 ));
    CascadeMux I__15832 (
            .O(N__68818),
            .I(N__68815));
    InMux I__15831 (
            .O(N__68815),
            .I(N__68812));
    LocalMux I__15830 (
            .O(N__68812),
            .I(N__68809));
    Span4Mux_h I__15829 (
            .O(N__68809),
            .I(N__68806));
    Span4Mux_v I__15828 (
            .O(N__68806),
            .I(N__68803));
    Odrv4 I__15827 (
            .O(N__68803),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20 ));
    InMux I__15826 (
            .O(N__68800),
            .I(N__68794));
    InMux I__15825 (
            .O(N__68799),
            .I(N__68794));
    LocalMux I__15824 (
            .O(N__68794),
            .I(N__68789));
    InMux I__15823 (
            .O(N__68793),
            .I(N__68786));
    InMux I__15822 (
            .O(N__68792),
            .I(N__68783));
    Span12Mux_h I__15821 (
            .O(N__68789),
            .I(N__68776));
    LocalMux I__15820 (
            .O(N__68786),
            .I(N__68776));
    LocalMux I__15819 (
            .O(N__68783),
            .I(N__68776));
    Odrv12 I__15818 (
            .O(N__68776),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21 ));
    InMux I__15817 (
            .O(N__68773),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15587 ));
    CascadeMux I__15816 (
            .O(N__68770),
            .I(N__68766));
    InMux I__15815 (
            .O(N__68769),
            .I(N__68763));
    InMux I__15814 (
            .O(N__68766),
            .I(N__68760));
    LocalMux I__15813 (
            .O(N__68763),
            .I(N__68757));
    LocalMux I__15812 (
            .O(N__68760),
            .I(N__68754));
    Span4Mux_v I__15811 (
            .O(N__68757),
            .I(N__68751));
    Odrv12 I__15810 (
            .O(N__68754),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29 ));
    Odrv4 I__15809 (
            .O(N__68751),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29 ));
    CascadeMux I__15808 (
            .O(N__68746),
            .I(N__68743));
    InMux I__15807 (
            .O(N__68743),
            .I(N__68740));
    LocalMux I__15806 (
            .O(N__68740),
            .I(N__68737));
    Span4Mux_v I__15805 (
            .O(N__68737),
            .I(N__68734));
    Span4Mux_h I__15804 (
            .O(N__68734),
            .I(N__68731));
    Odrv4 I__15803 (
            .O(N__68731),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21 ));
    InMux I__15802 (
            .O(N__68728),
            .I(N__68722));
    InMux I__15801 (
            .O(N__68727),
            .I(N__68722));
    LocalMux I__15800 (
            .O(N__68722),
            .I(N__68717));
    InMux I__15799 (
            .O(N__68721),
            .I(N__68714));
    InMux I__15798 (
            .O(N__68720),
            .I(N__68711));
    Sp12to4 I__15797 (
            .O(N__68717),
            .I(N__68704));
    LocalMux I__15796 (
            .O(N__68714),
            .I(N__68704));
    LocalMux I__15795 (
            .O(N__68711),
            .I(N__68704));
    Odrv12 I__15794 (
            .O(N__68704),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22 ));
    InMux I__15793 (
            .O(N__68701),
            .I(bfn_24_19_0_));
    InMux I__15792 (
            .O(N__68698),
            .I(N__68694));
    InMux I__15791 (
            .O(N__68697),
            .I(N__68691));
    LocalMux I__15790 (
            .O(N__68694),
            .I(N__68688));
    LocalMux I__15789 (
            .O(N__68691),
            .I(N__68685));
    Span4Mux_v I__15788 (
            .O(N__68688),
            .I(N__68682));
    Span4Mux_v I__15787 (
            .O(N__68685),
            .I(N__68679));
    Odrv4 I__15786 (
            .O(N__68682),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30 ));
    Odrv4 I__15785 (
            .O(N__68679),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30 ));
    CascadeMux I__15784 (
            .O(N__68674),
            .I(N__68671));
    InMux I__15783 (
            .O(N__68671),
            .I(N__68668));
    LocalMux I__15782 (
            .O(N__68668),
            .I(N__68665));
    Span4Mux_v I__15781 (
            .O(N__68665),
            .I(N__68662));
    Odrv4 I__15780 (
            .O(N__68662),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22 ));
    InMux I__15779 (
            .O(N__68659),
            .I(N__68653));
    InMux I__15778 (
            .O(N__68658),
            .I(N__68653));
    LocalMux I__15777 (
            .O(N__68653),
            .I(N__68650));
    Span4Mux_v I__15776 (
            .O(N__68650),
            .I(N__68645));
    InMux I__15775 (
            .O(N__68649),
            .I(N__68642));
    InMux I__15774 (
            .O(N__68648),
            .I(N__68639));
    Span4Mux_v I__15773 (
            .O(N__68645),
            .I(N__68636));
    LocalMux I__15772 (
            .O(N__68642),
            .I(N__68631));
    LocalMux I__15771 (
            .O(N__68639),
            .I(N__68631));
    Odrv4 I__15770 (
            .O(N__68636),
            .I(\foc.preSatVoltage_23_adj_2328 ));
    Odrv12 I__15769 (
            .O(N__68631),
            .I(\foc.preSatVoltage_23_adj_2328 ));
    InMux I__15768 (
            .O(N__68626),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15589 ));
    CascadeMux I__15767 (
            .O(N__68623),
            .I(N__68620));
    InMux I__15766 (
            .O(N__68620),
            .I(N__68617));
    LocalMux I__15765 (
            .O(N__68617),
            .I(N__68614));
    Span4Mux_v I__15764 (
            .O(N__68614),
            .I(N__68611));
    Odrv4 I__15763 (
            .O(N__68611),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23 ));
    InMux I__15762 (
            .O(N__68608),
            .I(N__68602));
    InMux I__15761 (
            .O(N__68607),
            .I(N__68602));
    LocalMux I__15760 (
            .O(N__68602),
            .I(N__68598));
    InMux I__15759 (
            .O(N__68601),
            .I(N__68595));
    Span4Mux_v I__15758 (
            .O(N__68598),
            .I(N__68591));
    LocalMux I__15757 (
            .O(N__68595),
            .I(N__68588));
    InMux I__15756 (
            .O(N__68594),
            .I(N__68585));
    Span4Mux_h I__15755 (
            .O(N__68591),
            .I(N__68582));
    Sp12to4 I__15754 (
            .O(N__68588),
            .I(N__68577));
    LocalMux I__15753 (
            .O(N__68585),
            .I(N__68577));
    Odrv4 I__15752 (
            .O(N__68582),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24 ));
    Odrv12 I__15751 (
            .O(N__68577),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24 ));
    InMux I__15750 (
            .O(N__68572),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15590 ));
    InMux I__15749 (
            .O(N__68569),
            .I(N__68566));
    LocalMux I__15748 (
            .O(N__68566),
            .I(N__68563));
    Span4Mux_v I__15747 (
            .O(N__68563),
            .I(N__68560));
    Odrv4 I__15746 (
            .O(N__68560),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24 ));
    CascadeMux I__15745 (
            .O(N__68557),
            .I(N__68554));
    InMux I__15744 (
            .O(N__68554),
            .I(N__68551));
    LocalMux I__15743 (
            .O(N__68551),
            .I(N__68546));
    InMux I__15742 (
            .O(N__68550),
            .I(N__68543));
    CascadeMux I__15741 (
            .O(N__68549),
            .I(N__68540));
    Span4Mux_v I__15740 (
            .O(N__68546),
            .I(N__68537));
    LocalMux I__15739 (
            .O(N__68543),
            .I(N__68534));
    InMux I__15738 (
            .O(N__68540),
            .I(N__68531));
    Span4Mux_h I__15737 (
            .O(N__68537),
            .I(N__68528));
    Sp12to4 I__15736 (
            .O(N__68534),
            .I(N__68523));
    LocalMux I__15735 (
            .O(N__68531),
            .I(N__68523));
    Odrv4 I__15734 (
            .O(N__68528),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25 ));
    Odrv12 I__15733 (
            .O(N__68523),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25 ));
    InMux I__15732 (
            .O(N__68518),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15591 ));
    CascadeMux I__15731 (
            .O(N__68515),
            .I(N__68512));
    InMux I__15730 (
            .O(N__68512),
            .I(N__68509));
    LocalMux I__15729 (
            .O(N__68509),
            .I(N__68506));
    Span4Mux_v I__15728 (
            .O(N__68506),
            .I(N__68503));
    Odrv4 I__15727 (
            .O(N__68503),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25 ));
    CascadeMux I__15726 (
            .O(N__68500),
            .I(N__68497));
    InMux I__15725 (
            .O(N__68497),
            .I(N__68493));
    InMux I__15724 (
            .O(N__68496),
            .I(N__68490));
    LocalMux I__15723 (
            .O(N__68493),
            .I(N__68487));
    LocalMux I__15722 (
            .O(N__68490),
            .I(N__68484));
    Odrv12 I__15721 (
            .O(N__68487),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20 ));
    Odrv12 I__15720 (
            .O(N__68484),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20 ));
    CascadeMux I__15719 (
            .O(N__68479),
            .I(N__68476));
    InMux I__15718 (
            .O(N__68476),
            .I(N__68473));
    LocalMux I__15717 (
            .O(N__68473),
            .I(N__68470));
    Span4Mux_v I__15716 (
            .O(N__68470),
            .I(N__68467));
    Odrv4 I__15715 (
            .O(N__68467),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12 ));
    InMux I__15714 (
            .O(N__68464),
            .I(N__68461));
    LocalMux I__15713 (
            .O(N__68461),
            .I(N__68456));
    InMux I__15712 (
            .O(N__68460),
            .I(N__68453));
    InMux I__15711 (
            .O(N__68459),
            .I(N__68450));
    Span4Mux_h I__15710 (
            .O(N__68456),
            .I(N__68445));
    LocalMux I__15709 (
            .O(N__68453),
            .I(N__68445));
    LocalMux I__15708 (
            .O(N__68450),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13 ));
    Odrv4 I__15707 (
            .O(N__68445),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13 ));
    InMux I__15706 (
            .O(N__68440),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15579 ));
    InMux I__15705 (
            .O(N__68437),
            .I(N__68429));
    InMux I__15704 (
            .O(N__68436),
            .I(N__68429));
    InMux I__15703 (
            .O(N__68435),
            .I(N__68423));
    CascadeMux I__15702 (
            .O(N__68434),
            .I(N__68419));
    LocalMux I__15701 (
            .O(N__68429),
            .I(N__68415));
    InMux I__15700 (
            .O(N__68428),
            .I(N__68412));
    CascadeMux I__15699 (
            .O(N__68427),
            .I(N__68408));
    CascadeMux I__15698 (
            .O(N__68426),
            .I(N__68404));
    LocalMux I__15697 (
            .O(N__68423),
            .I(N__68387));
    InMux I__15696 (
            .O(N__68422),
            .I(N__68384));
    InMux I__15695 (
            .O(N__68419),
            .I(N__68379));
    InMux I__15694 (
            .O(N__68418),
            .I(N__68379));
    Span4Mux_v I__15693 (
            .O(N__68415),
            .I(N__68374));
    LocalMux I__15692 (
            .O(N__68412),
            .I(N__68374));
    InMux I__15691 (
            .O(N__68411),
            .I(N__68365));
    InMux I__15690 (
            .O(N__68408),
            .I(N__68365));
    InMux I__15689 (
            .O(N__68407),
            .I(N__68365));
    InMux I__15688 (
            .O(N__68404),
            .I(N__68365));
    CascadeMux I__15687 (
            .O(N__68403),
            .I(N__68361));
    CascadeMux I__15686 (
            .O(N__68402),
            .I(N__68357));
    CascadeMux I__15685 (
            .O(N__68401),
            .I(N__68353));
    CascadeMux I__15684 (
            .O(N__68400),
            .I(N__68349));
    CascadeMux I__15683 (
            .O(N__68399),
            .I(N__68345));
    CascadeMux I__15682 (
            .O(N__68398),
            .I(N__68341));
    CascadeMux I__15681 (
            .O(N__68397),
            .I(N__68337));
    CascadeMux I__15680 (
            .O(N__68396),
            .I(N__68333));
    CascadeMux I__15679 (
            .O(N__68395),
            .I(N__68329));
    CascadeMux I__15678 (
            .O(N__68394),
            .I(N__68326));
    CascadeMux I__15677 (
            .O(N__68393),
            .I(N__68323));
    CascadeMux I__15676 (
            .O(N__68392),
            .I(N__68320));
    CascadeMux I__15675 (
            .O(N__68391),
            .I(N__68317));
    CascadeMux I__15674 (
            .O(N__68390),
            .I(N__68314));
    Span4Mux_v I__15673 (
            .O(N__68387),
            .I(N__68311));
    LocalMux I__15672 (
            .O(N__68384),
            .I(N__68306));
    LocalMux I__15671 (
            .O(N__68379),
            .I(N__68306));
    Span4Mux_v I__15670 (
            .O(N__68374),
            .I(N__68303));
    LocalMux I__15669 (
            .O(N__68365),
            .I(N__68300));
    InMux I__15668 (
            .O(N__68364),
            .I(N__68283));
    InMux I__15667 (
            .O(N__68361),
            .I(N__68283));
    InMux I__15666 (
            .O(N__68360),
            .I(N__68283));
    InMux I__15665 (
            .O(N__68357),
            .I(N__68283));
    InMux I__15664 (
            .O(N__68356),
            .I(N__68283));
    InMux I__15663 (
            .O(N__68353),
            .I(N__68283));
    InMux I__15662 (
            .O(N__68352),
            .I(N__68283));
    InMux I__15661 (
            .O(N__68349),
            .I(N__68283));
    InMux I__15660 (
            .O(N__68348),
            .I(N__68266));
    InMux I__15659 (
            .O(N__68345),
            .I(N__68266));
    InMux I__15658 (
            .O(N__68344),
            .I(N__68266));
    InMux I__15657 (
            .O(N__68341),
            .I(N__68266));
    InMux I__15656 (
            .O(N__68340),
            .I(N__68266));
    InMux I__15655 (
            .O(N__68337),
            .I(N__68266));
    InMux I__15654 (
            .O(N__68336),
            .I(N__68266));
    InMux I__15653 (
            .O(N__68333),
            .I(N__68266));
    InMux I__15652 (
            .O(N__68332),
            .I(N__68257));
    InMux I__15651 (
            .O(N__68329),
            .I(N__68257));
    InMux I__15650 (
            .O(N__68326),
            .I(N__68257));
    InMux I__15649 (
            .O(N__68323),
            .I(N__68257));
    InMux I__15648 (
            .O(N__68320),
            .I(N__68250));
    InMux I__15647 (
            .O(N__68317),
            .I(N__68250));
    InMux I__15646 (
            .O(N__68314),
            .I(N__68250));
    Span4Mux_v I__15645 (
            .O(N__68311),
            .I(N__68247));
    Span4Mux_v I__15644 (
            .O(N__68306),
            .I(N__68244));
    Span4Mux_h I__15643 (
            .O(N__68303),
            .I(N__68231));
    Span4Mux_v I__15642 (
            .O(N__68300),
            .I(N__68231));
    LocalMux I__15641 (
            .O(N__68283),
            .I(N__68231));
    LocalMux I__15640 (
            .O(N__68266),
            .I(N__68231));
    LocalMux I__15639 (
            .O(N__68257),
            .I(N__68231));
    LocalMux I__15638 (
            .O(N__68250),
            .I(N__68231));
    Span4Mux_v I__15637 (
            .O(N__68247),
            .I(N__68226));
    Span4Mux_h I__15636 (
            .O(N__68244),
            .I(N__68226));
    Span4Mux_v I__15635 (
            .O(N__68231),
            .I(N__68223));
    Odrv4 I__15634 (
            .O(N__68226),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__15633 (
            .O(N__68223),
            .I(CONSTANT_ONE_NET));
    InMux I__15632 (
            .O(N__68218),
            .I(N__68215));
    LocalMux I__15631 (
            .O(N__68215),
            .I(N__68211));
    InMux I__15630 (
            .O(N__68214),
            .I(N__68208));
    Odrv4 I__15629 (
            .O(N__68211),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21 ));
    LocalMux I__15628 (
            .O(N__68208),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21 ));
    CascadeMux I__15627 (
            .O(N__68203),
            .I(N__68200));
    InMux I__15626 (
            .O(N__68200),
            .I(N__68197));
    LocalMux I__15625 (
            .O(N__68197),
            .I(N__68194));
    Span4Mux_v I__15624 (
            .O(N__68194),
            .I(N__68191));
    Odrv4 I__15623 (
            .O(N__68191),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13 ));
    InMux I__15622 (
            .O(N__68188),
            .I(N__68184));
    InMux I__15621 (
            .O(N__68187),
            .I(N__68181));
    LocalMux I__15620 (
            .O(N__68184),
            .I(N__68174));
    LocalMux I__15619 (
            .O(N__68181),
            .I(N__68174));
    CascadeMux I__15618 (
            .O(N__68180),
            .I(N__68171));
    CascadeMux I__15617 (
            .O(N__68179),
            .I(N__68168));
    Span4Mux_v I__15616 (
            .O(N__68174),
            .I(N__68165));
    InMux I__15615 (
            .O(N__68171),
            .I(N__68162));
    InMux I__15614 (
            .O(N__68168),
            .I(N__68159));
    Span4Mux_v I__15613 (
            .O(N__68165),
            .I(N__68156));
    LocalMux I__15612 (
            .O(N__68162),
            .I(N__68151));
    LocalMux I__15611 (
            .O(N__68159),
            .I(N__68151));
    Odrv4 I__15610 (
            .O(N__68156),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14 ));
    Odrv12 I__15609 (
            .O(N__68151),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14 ));
    InMux I__15608 (
            .O(N__68146),
            .I(bfn_24_18_0_));
    CascadeMux I__15607 (
            .O(N__68143),
            .I(N__68140));
    InMux I__15606 (
            .O(N__68140),
            .I(N__68137));
    LocalMux I__15605 (
            .O(N__68137),
            .I(N__68133));
    InMux I__15604 (
            .O(N__68136),
            .I(N__68130));
    Odrv4 I__15603 (
            .O(N__68133),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22 ));
    LocalMux I__15602 (
            .O(N__68130),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22 ));
    CascadeMux I__15601 (
            .O(N__68125),
            .I(N__68122));
    InMux I__15600 (
            .O(N__68122),
            .I(N__68119));
    LocalMux I__15599 (
            .O(N__68119),
            .I(N__68116));
    Span4Mux_h I__15598 (
            .O(N__68116),
            .I(N__68113));
    Span4Mux_v I__15597 (
            .O(N__68113),
            .I(N__68110));
    Odrv4 I__15596 (
            .O(N__68110),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14 ));
    InMux I__15595 (
            .O(N__68107),
            .I(N__68101));
    InMux I__15594 (
            .O(N__68106),
            .I(N__68101));
    LocalMux I__15593 (
            .O(N__68101),
            .I(N__68096));
    InMux I__15592 (
            .O(N__68100),
            .I(N__68091));
    InMux I__15591 (
            .O(N__68099),
            .I(N__68091));
    Sp12to4 I__15590 (
            .O(N__68096),
            .I(N__68086));
    LocalMux I__15589 (
            .O(N__68091),
            .I(N__68086));
    Odrv12 I__15588 (
            .O(N__68086),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15 ));
    InMux I__15587 (
            .O(N__68083),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15581 ));
    InMux I__15586 (
            .O(N__68080),
            .I(N__68077));
    LocalMux I__15585 (
            .O(N__68077),
            .I(N__68073));
    InMux I__15584 (
            .O(N__68076),
            .I(N__68070));
    Odrv4 I__15583 (
            .O(N__68073),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23 ));
    LocalMux I__15582 (
            .O(N__68070),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23 ));
    CascadeMux I__15581 (
            .O(N__68065),
            .I(N__68062));
    InMux I__15580 (
            .O(N__68062),
            .I(N__68059));
    LocalMux I__15579 (
            .O(N__68059),
            .I(N__68056));
    Span4Mux_v I__15578 (
            .O(N__68056),
            .I(N__68053));
    Odrv4 I__15577 (
            .O(N__68053),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15 ));
    InMux I__15576 (
            .O(N__68050),
            .I(N__68042));
    InMux I__15575 (
            .O(N__68049),
            .I(N__68042));
    InMux I__15574 (
            .O(N__68048),
            .I(N__68037));
    InMux I__15573 (
            .O(N__68047),
            .I(N__68037));
    LocalMux I__15572 (
            .O(N__68042),
            .I(N__68034));
    LocalMux I__15571 (
            .O(N__68037),
            .I(N__68031));
    Sp12to4 I__15570 (
            .O(N__68034),
            .I(N__68028));
    Span4Mux_v I__15569 (
            .O(N__68031),
            .I(N__68025));
    Odrv12 I__15568 (
            .O(N__68028),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16 ));
    Odrv4 I__15567 (
            .O(N__68025),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16 ));
    InMux I__15566 (
            .O(N__68020),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15582 ));
    InMux I__15565 (
            .O(N__68017),
            .I(N__68014));
    LocalMux I__15564 (
            .O(N__68014),
            .I(N__68010));
    InMux I__15563 (
            .O(N__68013),
            .I(N__68007));
    Span4Mux_v I__15562 (
            .O(N__68010),
            .I(N__68004));
    LocalMux I__15561 (
            .O(N__68007),
            .I(N__68001));
    Odrv4 I__15560 (
            .O(N__68004),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24 ));
    Odrv4 I__15559 (
            .O(N__68001),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24 ));
    CascadeMux I__15558 (
            .O(N__67996),
            .I(N__67993));
    InMux I__15557 (
            .O(N__67993),
            .I(N__67990));
    LocalMux I__15556 (
            .O(N__67990),
            .I(N__67987));
    Span4Mux_v I__15555 (
            .O(N__67987),
            .I(N__67984));
    Span4Mux_h I__15554 (
            .O(N__67984),
            .I(N__67981));
    Odrv4 I__15553 (
            .O(N__67981),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16 ));
    InMux I__15552 (
            .O(N__67978),
            .I(N__67974));
    InMux I__15551 (
            .O(N__67977),
            .I(N__67971));
    LocalMux I__15550 (
            .O(N__67974),
            .I(N__67965));
    LocalMux I__15549 (
            .O(N__67971),
            .I(N__67965));
    InMux I__15548 (
            .O(N__67970),
            .I(N__67961));
    Span4Mux_h I__15547 (
            .O(N__67965),
            .I(N__67958));
    InMux I__15546 (
            .O(N__67964),
            .I(N__67955));
    LocalMux I__15545 (
            .O(N__67961),
            .I(N__67952));
    Span4Mux_v I__15544 (
            .O(N__67958),
            .I(N__67949));
    LocalMux I__15543 (
            .O(N__67955),
            .I(N__67946));
    Span4Mux_v I__15542 (
            .O(N__67952),
            .I(N__67943));
    Odrv4 I__15541 (
            .O(N__67949),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17 ));
    Odrv12 I__15540 (
            .O(N__67946),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17 ));
    Odrv4 I__15539 (
            .O(N__67943),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17 ));
    InMux I__15538 (
            .O(N__67936),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15583 ));
    InMux I__15537 (
            .O(N__67933),
            .I(N__67930));
    LocalMux I__15536 (
            .O(N__67930),
            .I(N__67926));
    InMux I__15535 (
            .O(N__67929),
            .I(N__67923));
    Span4Mux_v I__15534 (
            .O(N__67926),
            .I(N__67918));
    LocalMux I__15533 (
            .O(N__67923),
            .I(N__67918));
    Odrv4 I__15532 (
            .O(N__67918),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25 ));
    CascadeMux I__15531 (
            .O(N__67915),
            .I(N__67912));
    InMux I__15530 (
            .O(N__67912),
            .I(N__67909));
    LocalMux I__15529 (
            .O(N__67909),
            .I(N__67906));
    Span4Mux_v I__15528 (
            .O(N__67906),
            .I(N__67903));
    Odrv4 I__15527 (
            .O(N__67903),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17 ));
    CascadeMux I__15526 (
            .O(N__67900),
            .I(N__67895));
    InMux I__15525 (
            .O(N__67899),
            .I(N__67892));
    InMux I__15524 (
            .O(N__67898),
            .I(N__67889));
    InMux I__15523 (
            .O(N__67895),
            .I(N__67886));
    LocalMux I__15522 (
            .O(N__67892),
            .I(N__67880));
    LocalMux I__15521 (
            .O(N__67889),
            .I(N__67880));
    LocalMux I__15520 (
            .O(N__67886),
            .I(N__67877));
    InMux I__15519 (
            .O(N__67885),
            .I(N__67874));
    Span4Mux_h I__15518 (
            .O(N__67880),
            .I(N__67867));
    Span4Mux_v I__15517 (
            .O(N__67877),
            .I(N__67867));
    LocalMux I__15516 (
            .O(N__67874),
            .I(N__67867));
    Odrv4 I__15515 (
            .O(N__67867),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18 ));
    InMux I__15514 (
            .O(N__67864),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15584 ));
    InMux I__15513 (
            .O(N__67861),
            .I(N__67858));
    LocalMux I__15512 (
            .O(N__67858),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20194 ));
    InMux I__15511 (
            .O(N__67855),
            .I(N__67852));
    LocalMux I__15510 (
            .O(N__67852),
            .I(N__67849));
    Span4Mux_v I__15509 (
            .O(N__67849),
            .I(N__67846));
    Odrv4 I__15508 (
            .O(N__67846),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6 ));
    InMux I__15507 (
            .O(N__67843),
            .I(N__67839));
    CascadeMux I__15506 (
            .O(N__67842),
            .I(N__67836));
    LocalMux I__15505 (
            .O(N__67839),
            .I(N__67833));
    InMux I__15504 (
            .O(N__67836),
            .I(N__67830));
    Odrv4 I__15503 (
            .O(N__67833),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14 ));
    LocalMux I__15502 (
            .O(N__67830),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14 ));
    InMux I__15501 (
            .O(N__67825),
            .I(bfn_24_17_0_));
    InMux I__15500 (
            .O(N__67822),
            .I(N__67819));
    LocalMux I__15499 (
            .O(N__67819),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20196 ));
    CascadeMux I__15498 (
            .O(N__67816),
            .I(N__67813));
    InMux I__15497 (
            .O(N__67813),
            .I(N__67810));
    LocalMux I__15496 (
            .O(N__67810),
            .I(N__67806));
    InMux I__15495 (
            .O(N__67809),
            .I(N__67803));
    Odrv4 I__15494 (
            .O(N__67806),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15 ));
    LocalMux I__15493 (
            .O(N__67803),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15 ));
    CascadeMux I__15492 (
            .O(N__67798),
            .I(N__67795));
    InMux I__15491 (
            .O(N__67795),
            .I(N__67792));
    LocalMux I__15490 (
            .O(N__67792),
            .I(N__67789));
    Span4Mux_v I__15489 (
            .O(N__67789),
            .I(N__67786));
    Odrv4 I__15488 (
            .O(N__67786),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7 ));
    InMux I__15487 (
            .O(N__67783),
            .I(N__67780));
    LocalMux I__15486 (
            .O(N__67780),
            .I(N__67776));
    InMux I__15485 (
            .O(N__67779),
            .I(N__67773));
    Odrv4 I__15484 (
            .O(N__67776),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20198 ));
    LocalMux I__15483 (
            .O(N__67773),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20198 ));
    InMux I__15482 (
            .O(N__67768),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15574 ));
    InMux I__15481 (
            .O(N__67765),
            .I(N__67762));
    LocalMux I__15480 (
            .O(N__67762),
            .I(N__67759));
    Span4Mux_v I__15479 (
            .O(N__67759),
            .I(N__67755));
    InMux I__15478 (
            .O(N__67758),
            .I(N__67752));
    Odrv4 I__15477 (
            .O(N__67755),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16 ));
    LocalMux I__15476 (
            .O(N__67752),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16 ));
    CascadeMux I__15475 (
            .O(N__67747),
            .I(N__67744));
    InMux I__15474 (
            .O(N__67744),
            .I(N__67741));
    LocalMux I__15473 (
            .O(N__67741),
            .I(N__67738));
    Span4Mux_v I__15472 (
            .O(N__67738),
            .I(N__67735));
    Odrv4 I__15471 (
            .O(N__67735),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8 ));
    InMux I__15470 (
            .O(N__67732),
            .I(N__67729));
    LocalMux I__15469 (
            .O(N__67729),
            .I(N__67725));
    InMux I__15468 (
            .O(N__67728),
            .I(N__67722));
    Odrv4 I__15467 (
            .O(N__67725),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9 ));
    LocalMux I__15466 (
            .O(N__67722),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9 ));
    InMux I__15465 (
            .O(N__67717),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15575 ));
    InMux I__15464 (
            .O(N__67714),
            .I(N__67711));
    LocalMux I__15463 (
            .O(N__67711),
            .I(N__67708));
    Span4Mux_v I__15462 (
            .O(N__67708),
            .I(N__67705));
    Odrv4 I__15461 (
            .O(N__67705),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9 ));
    InMux I__15460 (
            .O(N__67702),
            .I(N__67699));
    LocalMux I__15459 (
            .O(N__67699),
            .I(N__67696));
    Span4Mux_v I__15458 (
            .O(N__67696),
            .I(N__67692));
    CascadeMux I__15457 (
            .O(N__67695),
            .I(N__67689));
    Sp12to4 I__15456 (
            .O(N__67692),
            .I(N__67686));
    InMux I__15455 (
            .O(N__67689),
            .I(N__67683));
    Odrv12 I__15454 (
            .O(N__67686),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17 ));
    LocalMux I__15453 (
            .O(N__67683),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17 ));
    InMux I__15452 (
            .O(N__67678),
            .I(N__67674));
    InMux I__15451 (
            .O(N__67677),
            .I(N__67670));
    LocalMux I__15450 (
            .O(N__67674),
            .I(N__67667));
    InMux I__15449 (
            .O(N__67673),
            .I(N__67664));
    LocalMux I__15448 (
            .O(N__67670),
            .I(N__67661));
    Odrv4 I__15447 (
            .O(N__67667),
            .I(\foc.preSatVoltage_10_adj_2311 ));
    LocalMux I__15446 (
            .O(N__67664),
            .I(\foc.preSatVoltage_10_adj_2311 ));
    Odrv4 I__15445 (
            .O(N__67661),
            .I(\foc.preSatVoltage_10_adj_2311 ));
    InMux I__15444 (
            .O(N__67654),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15576 ));
    InMux I__15443 (
            .O(N__67651),
            .I(N__67647));
    InMux I__15442 (
            .O(N__67650),
            .I(N__67644));
    LocalMux I__15441 (
            .O(N__67647),
            .I(N__67641));
    LocalMux I__15440 (
            .O(N__67644),
            .I(N__67638));
    Odrv12 I__15439 (
            .O(N__67641),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18 ));
    Odrv4 I__15438 (
            .O(N__67638),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18 ));
    CascadeMux I__15437 (
            .O(N__67633),
            .I(N__67630));
    InMux I__15436 (
            .O(N__67630),
            .I(N__67627));
    LocalMux I__15435 (
            .O(N__67627),
            .I(N__67624));
    Span4Mux_v I__15434 (
            .O(N__67624),
            .I(N__67621));
    Odrv4 I__15433 (
            .O(N__67621),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10 ));
    InMux I__15432 (
            .O(N__67618),
            .I(N__67612));
    InMux I__15431 (
            .O(N__67617),
            .I(N__67612));
    LocalMux I__15430 (
            .O(N__67612),
            .I(N__67607));
    InMux I__15429 (
            .O(N__67611),
            .I(N__67604));
    InMux I__15428 (
            .O(N__67610),
            .I(N__67601));
    Span4Mux_h I__15427 (
            .O(N__67607),
            .I(N__67596));
    LocalMux I__15426 (
            .O(N__67604),
            .I(N__67596));
    LocalMux I__15425 (
            .O(N__67601),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11 ));
    Odrv4 I__15424 (
            .O(N__67596),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11 ));
    InMux I__15423 (
            .O(N__67591),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15577 ));
    CascadeMux I__15422 (
            .O(N__67588),
            .I(N__67585));
    InMux I__15421 (
            .O(N__67585),
            .I(N__67582));
    LocalMux I__15420 (
            .O(N__67582),
            .I(N__67578));
    InMux I__15419 (
            .O(N__67581),
            .I(N__67575));
    Odrv4 I__15418 (
            .O(N__67578),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19 ));
    LocalMux I__15417 (
            .O(N__67575),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19 ));
    CascadeMux I__15416 (
            .O(N__67570),
            .I(N__67567));
    InMux I__15415 (
            .O(N__67567),
            .I(N__67564));
    LocalMux I__15414 (
            .O(N__67564),
            .I(N__67561));
    Span4Mux_v I__15413 (
            .O(N__67561),
            .I(N__67558));
    Odrv4 I__15412 (
            .O(N__67558),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11 ));
    InMux I__15411 (
            .O(N__67555),
            .I(N__67549));
    InMux I__15410 (
            .O(N__67554),
            .I(N__67549));
    LocalMux I__15409 (
            .O(N__67549),
            .I(N__67544));
    InMux I__15408 (
            .O(N__67548),
            .I(N__67541));
    InMux I__15407 (
            .O(N__67547),
            .I(N__67538));
    Span4Mux_v I__15406 (
            .O(N__67544),
            .I(N__67535));
    LocalMux I__15405 (
            .O(N__67541),
            .I(N__67530));
    LocalMux I__15404 (
            .O(N__67538),
            .I(N__67530));
    Odrv4 I__15403 (
            .O(N__67535),
            .I(\foc.preSatVoltage_12_adj_2330 ));
    Odrv4 I__15402 (
            .O(N__67530),
            .I(\foc.preSatVoltage_12_adj_2330 ));
    InMux I__15401 (
            .O(N__67525),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15578 ));
    InMux I__15400 (
            .O(N__67522),
            .I(N__67519));
    LocalMux I__15399 (
            .O(N__67519),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455 ));
    InMux I__15398 (
            .O(N__67516),
            .I(N__67513));
    LocalMux I__15397 (
            .O(N__67513),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690 ));
    CascadeMux I__15396 (
            .O(N__67510),
            .I(N__67507));
    InMux I__15395 (
            .O(N__67507),
            .I(N__67504));
    LocalMux I__15394 (
            .O(N__67504),
            .I(N__67500));
    InMux I__15393 (
            .O(N__67503),
            .I(N__67497));
    Odrv4 I__15392 (
            .O(N__67500),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0 ));
    LocalMux I__15391 (
            .O(N__67497),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0 ));
    InMux I__15390 (
            .O(N__67492),
            .I(N__67489));
    LocalMux I__15389 (
            .O(N__67489),
            .I(N__67486));
    Span12Mux_h I__15388 (
            .O(N__67486),
            .I(N__67482));
    InMux I__15387 (
            .O(N__67485),
            .I(N__67479));
    Odrv12 I__15386 (
            .O(N__67482),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8 ));
    LocalMux I__15385 (
            .O(N__67479),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8 ));
    CascadeMux I__15384 (
            .O(N__67474),
            .I(N__67471));
    InMux I__15383 (
            .O(N__67471),
            .I(N__67468));
    LocalMux I__15382 (
            .O(N__67468),
            .I(N__67452));
    CascadeMux I__15381 (
            .O(N__67467),
            .I(N__67449));
    CascadeMux I__15380 (
            .O(N__67466),
            .I(N__67446));
    CascadeMux I__15379 (
            .O(N__67465),
            .I(N__67443));
    CascadeMux I__15378 (
            .O(N__67464),
            .I(N__67439));
    CascadeMux I__15377 (
            .O(N__67463),
            .I(N__67436));
    CascadeMux I__15376 (
            .O(N__67462),
            .I(N__67433));
    CascadeMux I__15375 (
            .O(N__67461),
            .I(N__67430));
    CascadeMux I__15374 (
            .O(N__67460),
            .I(N__67427));
    CascadeMux I__15373 (
            .O(N__67459),
            .I(N__67422));
    CascadeMux I__15372 (
            .O(N__67458),
            .I(N__67418));
    CascadeMux I__15371 (
            .O(N__67457),
            .I(N__67414));
    CascadeMux I__15370 (
            .O(N__67456),
            .I(N__67410));
    CascadeMux I__15369 (
            .O(N__67455),
            .I(N__67406));
    Span4Mux_v I__15368 (
            .O(N__67452),
            .I(N__67401));
    InMux I__15367 (
            .O(N__67449),
            .I(N__67398));
    InMux I__15366 (
            .O(N__67446),
            .I(N__67392));
    InMux I__15365 (
            .O(N__67443),
            .I(N__67389));
    CascadeMux I__15364 (
            .O(N__67442),
            .I(N__67386));
    InMux I__15363 (
            .O(N__67439),
            .I(N__67381));
    InMux I__15362 (
            .O(N__67436),
            .I(N__67381));
    InMux I__15361 (
            .O(N__67433),
            .I(N__67372));
    InMux I__15360 (
            .O(N__67430),
            .I(N__67372));
    InMux I__15359 (
            .O(N__67427),
            .I(N__67372));
    InMux I__15358 (
            .O(N__67426),
            .I(N__67372));
    InMux I__15357 (
            .O(N__67425),
            .I(N__67355));
    InMux I__15356 (
            .O(N__67422),
            .I(N__67355));
    InMux I__15355 (
            .O(N__67421),
            .I(N__67355));
    InMux I__15354 (
            .O(N__67418),
            .I(N__67355));
    InMux I__15353 (
            .O(N__67417),
            .I(N__67355));
    InMux I__15352 (
            .O(N__67414),
            .I(N__67355));
    InMux I__15351 (
            .O(N__67413),
            .I(N__67355));
    InMux I__15350 (
            .O(N__67410),
            .I(N__67355));
    CascadeMux I__15349 (
            .O(N__67409),
            .I(N__67352));
    InMux I__15348 (
            .O(N__67406),
            .I(N__67348));
    CascadeMux I__15347 (
            .O(N__67405),
            .I(N__67345));
    CascadeMux I__15346 (
            .O(N__67404),
            .I(N__67342));
    Span4Mux_h I__15345 (
            .O(N__67401),
            .I(N__67337));
    LocalMux I__15344 (
            .O(N__67398),
            .I(N__67337));
    CascadeMux I__15343 (
            .O(N__67397),
            .I(N__67334));
    CascadeMux I__15342 (
            .O(N__67396),
            .I(N__67331));
    CascadeMux I__15341 (
            .O(N__67395),
            .I(N__67328));
    LocalMux I__15340 (
            .O(N__67392),
            .I(N__67323));
    LocalMux I__15339 (
            .O(N__67389),
            .I(N__67323));
    InMux I__15338 (
            .O(N__67386),
            .I(N__67320));
    LocalMux I__15337 (
            .O(N__67381),
            .I(N__67315));
    LocalMux I__15336 (
            .O(N__67372),
            .I(N__67315));
    LocalMux I__15335 (
            .O(N__67355),
            .I(N__67312));
    InMux I__15334 (
            .O(N__67352),
            .I(N__67309));
    CascadeMux I__15333 (
            .O(N__67351),
            .I(N__67306));
    LocalMux I__15332 (
            .O(N__67348),
            .I(N__67303));
    InMux I__15331 (
            .O(N__67345),
            .I(N__67300));
    InMux I__15330 (
            .O(N__67342),
            .I(N__67297));
    Span4Mux_v I__15329 (
            .O(N__67337),
            .I(N__67293));
    InMux I__15328 (
            .O(N__67334),
            .I(N__67290));
    InMux I__15327 (
            .O(N__67331),
            .I(N__67287));
    InMux I__15326 (
            .O(N__67328),
            .I(N__67284));
    Span4Mux_v I__15325 (
            .O(N__67323),
            .I(N__67279));
    LocalMux I__15324 (
            .O(N__67320),
            .I(N__67279));
    Span4Mux_v I__15323 (
            .O(N__67315),
            .I(N__67272));
    Span4Mux_v I__15322 (
            .O(N__67312),
            .I(N__67272));
    LocalMux I__15321 (
            .O(N__67309),
            .I(N__67272));
    InMux I__15320 (
            .O(N__67306),
            .I(N__67269));
    Span4Mux_v I__15319 (
            .O(N__67303),
            .I(N__67262));
    LocalMux I__15318 (
            .O(N__67300),
            .I(N__67262));
    LocalMux I__15317 (
            .O(N__67297),
            .I(N__67262));
    CascadeMux I__15316 (
            .O(N__67296),
            .I(N__67259));
    Span4Mux_h I__15315 (
            .O(N__67293),
            .I(N__67254));
    LocalMux I__15314 (
            .O(N__67290),
            .I(N__67254));
    LocalMux I__15313 (
            .O(N__67287),
            .I(N__67243));
    LocalMux I__15312 (
            .O(N__67284),
            .I(N__67243));
    Span4Mux_h I__15311 (
            .O(N__67279),
            .I(N__67243));
    Span4Mux_h I__15310 (
            .O(N__67272),
            .I(N__67243));
    LocalMux I__15309 (
            .O(N__67269),
            .I(N__67243));
    Span4Mux_v I__15308 (
            .O(N__67262),
            .I(N__67240));
    InMux I__15307 (
            .O(N__67259),
            .I(N__67237));
    Span4Mux_v I__15306 (
            .O(N__67254),
            .I(N__67234));
    Span4Mux_v I__15305 (
            .O(N__67243),
            .I(N__67227));
    Span4Mux_v I__15304 (
            .O(N__67240),
            .I(N__67227));
    LocalMux I__15303 (
            .O(N__67237),
            .I(N__67227));
    Span4Mux_v I__15302 (
            .O(N__67234),
            .I(N__67224));
    Span4Mux_v I__15301 (
            .O(N__67227),
            .I(N__67221));
    Odrv4 I__15300 (
            .O(N__67224),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0 ));
    Odrv4 I__15299 (
            .O(N__67221),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0 ));
    InMux I__15298 (
            .O(N__67216),
            .I(N__67213));
    LocalMux I__15297 (
            .O(N__67213),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20184 ));
    InMux I__15296 (
            .O(N__67210),
            .I(N__67207));
    LocalMux I__15295 (
            .O(N__67207),
            .I(N__67204));
    Span4Mux_v I__15294 (
            .O(N__67204),
            .I(N__67200));
    InMux I__15293 (
            .O(N__67203),
            .I(N__67197));
    Odrv4 I__15292 (
            .O(N__67200),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9 ));
    LocalMux I__15291 (
            .O(N__67197),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9 ));
    CascadeMux I__15290 (
            .O(N__67192),
            .I(N__67189));
    InMux I__15289 (
            .O(N__67189),
            .I(N__67186));
    LocalMux I__15288 (
            .O(N__67186),
            .I(N__67183));
    Span4Mux_v I__15287 (
            .O(N__67183),
            .I(N__67180));
    Odrv4 I__15286 (
            .O(N__67180),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1 ));
    InMux I__15285 (
            .O(N__67177),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15568 ));
    InMux I__15284 (
            .O(N__67174),
            .I(N__67171));
    LocalMux I__15283 (
            .O(N__67171),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20186 ));
    InMux I__15282 (
            .O(N__67168),
            .I(N__67165));
    LocalMux I__15281 (
            .O(N__67165),
            .I(N__67162));
    Span4Mux_v I__15280 (
            .O(N__67162),
            .I(N__67158));
    InMux I__15279 (
            .O(N__67161),
            .I(N__67155));
    Odrv4 I__15278 (
            .O(N__67158),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10 ));
    LocalMux I__15277 (
            .O(N__67155),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10 ));
    CascadeMux I__15276 (
            .O(N__67150),
            .I(N__67147));
    InMux I__15275 (
            .O(N__67147),
            .I(N__67144));
    LocalMux I__15274 (
            .O(N__67144),
            .I(N__67141));
    Span4Mux_v I__15273 (
            .O(N__67141),
            .I(N__67138));
    Odrv4 I__15272 (
            .O(N__67138),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2 ));
    InMux I__15271 (
            .O(N__67135),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15569 ));
    InMux I__15270 (
            .O(N__67132),
            .I(N__67129));
    LocalMux I__15269 (
            .O(N__67129),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20188 ));
    CascadeMux I__15268 (
            .O(N__67126),
            .I(N__67123));
    InMux I__15267 (
            .O(N__67123),
            .I(N__67120));
    LocalMux I__15266 (
            .O(N__67120),
            .I(N__67117));
    Span4Mux_v I__15265 (
            .O(N__67117),
            .I(N__67113));
    InMux I__15264 (
            .O(N__67116),
            .I(N__67110));
    Odrv4 I__15263 (
            .O(N__67113),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11 ));
    LocalMux I__15262 (
            .O(N__67110),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11 ));
    CascadeMux I__15261 (
            .O(N__67105),
            .I(N__67102));
    InMux I__15260 (
            .O(N__67102),
            .I(N__67099));
    LocalMux I__15259 (
            .O(N__67099),
            .I(N__67096));
    Span4Mux_v I__15258 (
            .O(N__67096),
            .I(N__67093));
    Odrv4 I__15257 (
            .O(N__67093),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3 ));
    InMux I__15256 (
            .O(N__67090),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15570 ));
    InMux I__15255 (
            .O(N__67087),
            .I(N__67084));
    LocalMux I__15254 (
            .O(N__67084),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20190 ));
    InMux I__15253 (
            .O(N__67081),
            .I(N__67078));
    LocalMux I__15252 (
            .O(N__67078),
            .I(N__67074));
    InMux I__15251 (
            .O(N__67077),
            .I(N__67071));
    Odrv4 I__15250 (
            .O(N__67074),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12 ));
    LocalMux I__15249 (
            .O(N__67071),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12 ));
    CascadeMux I__15248 (
            .O(N__67066),
            .I(N__67063));
    InMux I__15247 (
            .O(N__67063),
            .I(N__67060));
    LocalMux I__15246 (
            .O(N__67060),
            .I(N__67057));
    Span4Mux_v I__15245 (
            .O(N__67057),
            .I(N__67054));
    Odrv4 I__15244 (
            .O(N__67054),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4 ));
    InMux I__15243 (
            .O(N__67051),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15571 ));
    InMux I__15242 (
            .O(N__67048),
            .I(N__67045));
    LocalMux I__15241 (
            .O(N__67045),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20192 ));
    InMux I__15240 (
            .O(N__67042),
            .I(N__67039));
    LocalMux I__15239 (
            .O(N__67039),
            .I(N__67036));
    Span4Mux_h I__15238 (
            .O(N__67036),
            .I(N__67033));
    Span4Mux_v I__15237 (
            .O(N__67033),
            .I(N__67029));
    InMux I__15236 (
            .O(N__67032),
            .I(N__67026));
    Odrv4 I__15235 (
            .O(N__67029),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13 ));
    LocalMux I__15234 (
            .O(N__67026),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13 ));
    CascadeMux I__15233 (
            .O(N__67021),
            .I(N__67018));
    InMux I__15232 (
            .O(N__67018),
            .I(N__67015));
    LocalMux I__15231 (
            .O(N__67015),
            .I(N__67012));
    Span4Mux_v I__15230 (
            .O(N__67012),
            .I(N__67009));
    Span4Mux_h I__15229 (
            .O(N__67009),
            .I(N__67006));
    Odrv4 I__15228 (
            .O(N__67006),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5 ));
    InMux I__15227 (
            .O(N__67003),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15572 ));
    InMux I__15226 (
            .O(N__67000),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18277 ));
    InMux I__15225 (
            .O(N__66997),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767 ));
    CascadeMux I__15224 (
            .O(N__66994),
            .I(N__66991));
    InMux I__15223 (
            .O(N__66991),
            .I(N__66988));
    LocalMux I__15222 (
            .O(N__66988),
            .I(N__66985));
    Span4Mux_h I__15221 (
            .O(N__66985),
            .I(N__66982));
    Span4Mux_v I__15220 (
            .O(N__66982),
            .I(N__66979));
    Odrv4 I__15219 (
            .O(N__66979),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO ));
    InMux I__15218 (
            .O(N__66976),
            .I(N__66973));
    LocalMux I__15217 (
            .O(N__66973),
            .I(N__66970));
    Odrv4 I__15216 (
            .O(N__66970),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926 ));
    CascadeMux I__15215 (
            .O(N__66967),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_ ));
    InMux I__15214 (
            .O(N__66964),
            .I(N__66961));
    LocalMux I__15213 (
            .O(N__66961),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098 ));
    CascadeMux I__15212 (
            .O(N__66958),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_ ));
    CascadeMux I__15211 (
            .O(N__66955),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_ ));
    CascadeMux I__15210 (
            .O(N__66952),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_ ));
    InMux I__15209 (
            .O(N__66949),
            .I(N__66946));
    LocalMux I__15208 (
            .O(N__66946),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424 ));
    InMux I__15207 (
            .O(N__66943),
            .I(N__66940));
    LocalMux I__15206 (
            .O(N__66940),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851 ));
    InMux I__15205 (
            .O(N__66937),
            .I(N__66934));
    LocalMux I__15204 (
            .O(N__66934),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n369 ));
    CascadeMux I__15203 (
            .O(N__66931),
            .I(N__66917));
    CascadeMux I__15202 (
            .O(N__66930),
            .I(N__66914));
    CascadeMux I__15201 (
            .O(N__66929),
            .I(N__66910));
    CascadeMux I__15200 (
            .O(N__66928),
            .I(N__66907));
    CascadeMux I__15199 (
            .O(N__66927),
            .I(N__66904));
    CascadeMux I__15198 (
            .O(N__66926),
            .I(N__66901));
    CascadeMux I__15197 (
            .O(N__66925),
            .I(N__66898));
    CascadeMux I__15196 (
            .O(N__66924),
            .I(N__66895));
    CascadeMux I__15195 (
            .O(N__66923),
            .I(N__66892));
    InMux I__15194 (
            .O(N__66922),
            .I(N__66885));
    CascadeMux I__15193 (
            .O(N__66921),
            .I(N__66881));
    CascadeMux I__15192 (
            .O(N__66920),
            .I(N__66877));
    InMux I__15191 (
            .O(N__66917),
            .I(N__66870));
    InMux I__15190 (
            .O(N__66914),
            .I(N__66870));
    InMux I__15189 (
            .O(N__66913),
            .I(N__66861));
    InMux I__15188 (
            .O(N__66910),
            .I(N__66861));
    InMux I__15187 (
            .O(N__66907),
            .I(N__66861));
    InMux I__15186 (
            .O(N__66904),
            .I(N__66861));
    InMux I__15185 (
            .O(N__66901),
            .I(N__66852));
    InMux I__15184 (
            .O(N__66898),
            .I(N__66852));
    InMux I__15183 (
            .O(N__66895),
            .I(N__66852));
    InMux I__15182 (
            .O(N__66892),
            .I(N__66852));
    CascadeMux I__15181 (
            .O(N__66891),
            .I(N__66849));
    CascadeMux I__15180 (
            .O(N__66890),
            .I(N__66846));
    CascadeMux I__15179 (
            .O(N__66889),
            .I(N__66843));
    CascadeMux I__15178 (
            .O(N__66888),
            .I(N__66840));
    LocalMux I__15177 (
            .O(N__66885),
            .I(N__66837));
    InMux I__15176 (
            .O(N__66884),
            .I(N__66834));
    InMux I__15175 (
            .O(N__66881),
            .I(N__66831));
    CascadeMux I__15174 (
            .O(N__66880),
            .I(N__66825));
    InMux I__15173 (
            .O(N__66877),
            .I(N__66819));
    CascadeMux I__15172 (
            .O(N__66876),
            .I(N__66816));
    CascadeMux I__15171 (
            .O(N__66875),
            .I(N__66813));
    LocalMux I__15170 (
            .O(N__66870),
            .I(N__66808));
    LocalMux I__15169 (
            .O(N__66861),
            .I(N__66808));
    LocalMux I__15168 (
            .O(N__66852),
            .I(N__66805));
    InMux I__15167 (
            .O(N__66849),
            .I(N__66796));
    InMux I__15166 (
            .O(N__66846),
            .I(N__66796));
    InMux I__15165 (
            .O(N__66843),
            .I(N__66796));
    InMux I__15164 (
            .O(N__66840),
            .I(N__66796));
    Span4Mux_h I__15163 (
            .O(N__66837),
            .I(N__66789));
    LocalMux I__15162 (
            .O(N__66834),
            .I(N__66789));
    LocalMux I__15161 (
            .O(N__66831),
            .I(N__66789));
    CascadeMux I__15160 (
            .O(N__66830),
            .I(N__66786));
    CascadeMux I__15159 (
            .O(N__66829),
            .I(N__66783));
    CascadeMux I__15158 (
            .O(N__66828),
            .I(N__66779));
    InMux I__15157 (
            .O(N__66825),
            .I(N__66776));
    CascadeMux I__15156 (
            .O(N__66824),
            .I(N__66773));
    CascadeMux I__15155 (
            .O(N__66823),
            .I(N__66770));
    InMux I__15154 (
            .O(N__66822),
            .I(N__66767));
    LocalMux I__15153 (
            .O(N__66819),
            .I(N__66764));
    InMux I__15152 (
            .O(N__66816),
            .I(N__66761));
    InMux I__15151 (
            .O(N__66813),
            .I(N__66757));
    Span4Mux_v I__15150 (
            .O(N__66808),
            .I(N__66750));
    Span4Mux_h I__15149 (
            .O(N__66805),
            .I(N__66750));
    LocalMux I__15148 (
            .O(N__66796),
            .I(N__66750));
    Span4Mux_h I__15147 (
            .O(N__66789),
            .I(N__66747));
    InMux I__15146 (
            .O(N__66786),
            .I(N__66744));
    InMux I__15145 (
            .O(N__66783),
            .I(N__66741));
    InMux I__15144 (
            .O(N__66782),
            .I(N__66738));
    InMux I__15143 (
            .O(N__66779),
            .I(N__66735));
    LocalMux I__15142 (
            .O(N__66776),
            .I(N__66732));
    InMux I__15141 (
            .O(N__66773),
            .I(N__66729));
    InMux I__15140 (
            .O(N__66770),
            .I(N__66726));
    LocalMux I__15139 (
            .O(N__66767),
            .I(N__66723));
    Span4Mux_h I__15138 (
            .O(N__66764),
            .I(N__66720));
    LocalMux I__15137 (
            .O(N__66761),
            .I(N__66717));
    InMux I__15136 (
            .O(N__66760),
            .I(N__66714));
    LocalMux I__15135 (
            .O(N__66757),
            .I(N__66711));
    Span4Mux_v I__15134 (
            .O(N__66750),
            .I(N__66708));
    Sp12to4 I__15133 (
            .O(N__66747),
            .I(N__66705));
    LocalMux I__15132 (
            .O(N__66744),
            .I(N__66698));
    LocalMux I__15131 (
            .O(N__66741),
            .I(N__66698));
    LocalMux I__15130 (
            .O(N__66738),
            .I(N__66698));
    LocalMux I__15129 (
            .O(N__66735),
            .I(N__66695));
    Span4Mux_v I__15128 (
            .O(N__66732),
            .I(N__66688));
    LocalMux I__15127 (
            .O(N__66729),
            .I(N__66688));
    LocalMux I__15126 (
            .O(N__66726),
            .I(N__66688));
    Span4Mux_v I__15125 (
            .O(N__66723),
            .I(N__66685));
    Span4Mux_v I__15124 (
            .O(N__66720),
            .I(N__66676));
    Span4Mux_v I__15123 (
            .O(N__66717),
            .I(N__66676));
    LocalMux I__15122 (
            .O(N__66714),
            .I(N__66676));
    Span4Mux_v I__15121 (
            .O(N__66711),
            .I(N__66676));
    Span4Mux_h I__15120 (
            .O(N__66708),
            .I(N__66673));
    Span12Mux_s7_v I__15119 (
            .O(N__66705),
            .I(N__66668));
    Span12Mux_h I__15118 (
            .O(N__66698),
            .I(N__66668));
    Span4Mux_v I__15117 (
            .O(N__66695),
            .I(N__66663));
    Span4Mux_v I__15116 (
            .O(N__66688),
            .I(N__66663));
    Span4Mux_h I__15115 (
            .O(N__66685),
            .I(N__66658));
    Span4Mux_h I__15114 (
            .O(N__66676),
            .I(N__66658));
    Odrv4 I__15113 (
            .O(N__66673),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ));
    Odrv12 I__15112 (
            .O(N__66668),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ));
    Odrv4 I__15111 (
            .O(N__66663),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ));
    Odrv4 I__15110 (
            .O(N__66658),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ));
    InMux I__15109 (
            .O(N__66649),
            .I(N__66646));
    LocalMux I__15108 (
            .O(N__66646),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n415 ));
    InMux I__15107 (
            .O(N__66643),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18270 ));
    CascadeMux I__15106 (
            .O(N__66640),
            .I(N__66635));
    CascadeMux I__15105 (
            .O(N__66639),
            .I(N__66632));
    InMux I__15104 (
            .O(N__66638),
            .I(N__66626));
    InMux I__15103 (
            .O(N__66635),
            .I(N__66622));
    InMux I__15102 (
            .O(N__66632),
            .I(N__66619));
    CascadeMux I__15101 (
            .O(N__66631),
            .I(N__66616));
    CascadeMux I__15100 (
            .O(N__66630),
            .I(N__66613));
    CascadeMux I__15099 (
            .O(N__66629),
            .I(N__66609));
    LocalMux I__15098 (
            .O(N__66626),
            .I(N__66605));
    CascadeMux I__15097 (
            .O(N__66625),
            .I(N__66601));
    LocalMux I__15096 (
            .O(N__66622),
            .I(N__66595));
    LocalMux I__15095 (
            .O(N__66619),
            .I(N__66592));
    InMux I__15094 (
            .O(N__66616),
            .I(N__66589));
    InMux I__15093 (
            .O(N__66613),
            .I(N__66586));
    InMux I__15092 (
            .O(N__66612),
            .I(N__66583));
    InMux I__15091 (
            .O(N__66609),
            .I(N__66580));
    CascadeMux I__15090 (
            .O(N__66608),
            .I(N__66577));
    Span4Mux_v I__15089 (
            .O(N__66605),
            .I(N__66571));
    CascadeMux I__15088 (
            .O(N__66604),
            .I(N__66568));
    InMux I__15087 (
            .O(N__66601),
            .I(N__66565));
    CascadeMux I__15086 (
            .O(N__66600),
            .I(N__66562));
    CascadeMux I__15085 (
            .O(N__66599),
            .I(N__66559));
    InMux I__15084 (
            .O(N__66598),
            .I(N__66556));
    Span4Mux_v I__15083 (
            .O(N__66595),
            .I(N__66549));
    Span4Mux_v I__15082 (
            .O(N__66592),
            .I(N__66549));
    LocalMux I__15081 (
            .O(N__66589),
            .I(N__66549));
    LocalMux I__15080 (
            .O(N__66586),
            .I(N__66542));
    LocalMux I__15079 (
            .O(N__66583),
            .I(N__66542));
    LocalMux I__15078 (
            .O(N__66580),
            .I(N__66542));
    InMux I__15077 (
            .O(N__66577),
            .I(N__66539));
    CascadeMux I__15076 (
            .O(N__66576),
            .I(N__66535));
    CascadeMux I__15075 (
            .O(N__66575),
            .I(N__66531));
    CascadeMux I__15074 (
            .O(N__66574),
            .I(N__66528));
    Span4Mux_h I__15073 (
            .O(N__66571),
            .I(N__66525));
    InMux I__15072 (
            .O(N__66568),
            .I(N__66522));
    LocalMux I__15071 (
            .O(N__66565),
            .I(N__66512));
    InMux I__15070 (
            .O(N__66562),
            .I(N__66509));
    InMux I__15069 (
            .O(N__66559),
            .I(N__66506));
    LocalMux I__15068 (
            .O(N__66556),
            .I(N__66503));
    Span4Mux_h I__15067 (
            .O(N__66549),
            .I(N__66496));
    Span4Mux_v I__15066 (
            .O(N__66542),
            .I(N__66496));
    LocalMux I__15065 (
            .O(N__66539),
            .I(N__66496));
    InMux I__15064 (
            .O(N__66538),
            .I(N__66493));
    InMux I__15063 (
            .O(N__66535),
            .I(N__66486));
    InMux I__15062 (
            .O(N__66534),
            .I(N__66486));
    InMux I__15061 (
            .O(N__66531),
            .I(N__66486));
    InMux I__15060 (
            .O(N__66528),
            .I(N__66483));
    Span4Mux_v I__15059 (
            .O(N__66525),
            .I(N__66478));
    LocalMux I__15058 (
            .O(N__66522),
            .I(N__66478));
    CascadeMux I__15057 (
            .O(N__66521),
            .I(N__66475));
    CascadeMux I__15056 (
            .O(N__66520),
            .I(N__66472));
    CascadeMux I__15055 (
            .O(N__66519),
            .I(N__66469));
    CascadeMux I__15054 (
            .O(N__66518),
            .I(N__66465));
    CascadeMux I__15053 (
            .O(N__66517),
            .I(N__66461));
    CascadeMux I__15052 (
            .O(N__66516),
            .I(N__66458));
    CascadeMux I__15051 (
            .O(N__66515),
            .I(N__66455));
    Span4Mux_v I__15050 (
            .O(N__66512),
            .I(N__66448));
    LocalMux I__15049 (
            .O(N__66509),
            .I(N__66448));
    LocalMux I__15048 (
            .O(N__66506),
            .I(N__66448));
    Sp12to4 I__15047 (
            .O(N__66503),
            .I(N__66445));
    Span4Mux_v I__15046 (
            .O(N__66496),
            .I(N__66442));
    LocalMux I__15045 (
            .O(N__66493),
            .I(N__66435));
    LocalMux I__15044 (
            .O(N__66486),
            .I(N__66435));
    LocalMux I__15043 (
            .O(N__66483),
            .I(N__66435));
    Span4Mux_v I__15042 (
            .O(N__66478),
            .I(N__66432));
    InMux I__15041 (
            .O(N__66475),
            .I(N__66429));
    InMux I__15040 (
            .O(N__66472),
            .I(N__66416));
    InMux I__15039 (
            .O(N__66469),
            .I(N__66416));
    InMux I__15038 (
            .O(N__66468),
            .I(N__66416));
    InMux I__15037 (
            .O(N__66465),
            .I(N__66416));
    InMux I__15036 (
            .O(N__66464),
            .I(N__66416));
    InMux I__15035 (
            .O(N__66461),
            .I(N__66416));
    InMux I__15034 (
            .O(N__66458),
            .I(N__66411));
    InMux I__15033 (
            .O(N__66455),
            .I(N__66411));
    Span4Mux_v I__15032 (
            .O(N__66448),
            .I(N__66408));
    Span12Mux_s10_v I__15031 (
            .O(N__66445),
            .I(N__66393));
    Sp12to4 I__15030 (
            .O(N__66442),
            .I(N__66393));
    Span12Mux_s10_v I__15029 (
            .O(N__66435),
            .I(N__66393));
    Sp12to4 I__15028 (
            .O(N__66432),
            .I(N__66393));
    LocalMux I__15027 (
            .O(N__66429),
            .I(N__66393));
    LocalMux I__15026 (
            .O(N__66416),
            .I(N__66393));
    LocalMux I__15025 (
            .O(N__66411),
            .I(N__66393));
    Odrv4 I__15024 (
            .O(N__66408),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n126 ));
    Odrv12 I__15023 (
            .O(N__66393),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n126 ));
    CascadeMux I__15022 (
            .O(N__66388),
            .I(N__66385));
    InMux I__15021 (
            .O(N__66385),
            .I(N__66382));
    LocalMux I__15020 (
            .O(N__66382),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n418 ));
    InMux I__15019 (
            .O(N__66379),
            .I(N__66376));
    LocalMux I__15018 (
            .O(N__66376),
            .I(N__66373));
    Odrv4 I__15017 (
            .O(N__66373),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n464 ));
    InMux I__15016 (
            .O(N__66370),
            .I(bfn_23_28_0_));
    InMux I__15015 (
            .O(N__66367),
            .I(N__66364));
    LocalMux I__15014 (
            .O(N__66364),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n467 ));
    CascadeMux I__15013 (
            .O(N__66361),
            .I(N__66356));
    CascadeMux I__15012 (
            .O(N__66360),
            .I(N__66353));
    CascadeMux I__15011 (
            .O(N__66359),
            .I(N__66350));
    InMux I__15010 (
            .O(N__66356),
            .I(N__66340));
    InMux I__15009 (
            .O(N__66353),
            .I(N__66337));
    InMux I__15008 (
            .O(N__66350),
            .I(N__66334));
    CascadeMux I__15007 (
            .O(N__66349),
            .I(N__66331));
    CascadeMux I__15006 (
            .O(N__66348),
            .I(N__66328));
    CascadeMux I__15005 (
            .O(N__66347),
            .I(N__66324));
    CascadeMux I__15004 (
            .O(N__66346),
            .I(N__66321));
    CascadeMux I__15003 (
            .O(N__66345),
            .I(N__66318));
    CascadeMux I__15002 (
            .O(N__66344),
            .I(N__66315));
    CascadeMux I__15001 (
            .O(N__66343),
            .I(N__66312));
    LocalMux I__15000 (
            .O(N__66340),
            .I(N__66307));
    LocalMux I__14999 (
            .O(N__66337),
            .I(N__66307));
    LocalMux I__14998 (
            .O(N__66334),
            .I(N__66304));
    InMux I__14997 (
            .O(N__66331),
            .I(N__66301));
    InMux I__14996 (
            .O(N__66328),
            .I(N__66298));
    CascadeMux I__14995 (
            .O(N__66327),
            .I(N__66295));
    InMux I__14994 (
            .O(N__66324),
            .I(N__66290));
    InMux I__14993 (
            .O(N__66321),
            .I(N__66287));
    InMux I__14992 (
            .O(N__66318),
            .I(N__66283));
    InMux I__14991 (
            .O(N__66315),
            .I(N__66280));
    InMux I__14990 (
            .O(N__66312),
            .I(N__66277));
    Span4Mux_v I__14989 (
            .O(N__66307),
            .I(N__66268));
    Span4Mux_v I__14988 (
            .O(N__66304),
            .I(N__66268));
    LocalMux I__14987 (
            .O(N__66301),
            .I(N__66268));
    LocalMux I__14986 (
            .O(N__66298),
            .I(N__66268));
    InMux I__14985 (
            .O(N__66295),
            .I(N__66265));
    CascadeMux I__14984 (
            .O(N__66294),
            .I(N__66262));
    CascadeMux I__14983 (
            .O(N__66293),
            .I(N__66256));
    LocalMux I__14982 (
            .O(N__66290),
            .I(N__66253));
    LocalMux I__14981 (
            .O(N__66287),
            .I(N__66250));
    CascadeMux I__14980 (
            .O(N__66286),
            .I(N__66247));
    LocalMux I__14979 (
            .O(N__66283),
            .I(N__66244));
    LocalMux I__14978 (
            .O(N__66280),
            .I(N__66235));
    LocalMux I__14977 (
            .O(N__66277),
            .I(N__66235));
    Span4Mux_h I__14976 (
            .O(N__66268),
            .I(N__66235));
    LocalMux I__14975 (
            .O(N__66265),
            .I(N__66235));
    InMux I__14974 (
            .O(N__66262),
            .I(N__66232));
    CascadeMux I__14973 (
            .O(N__66261),
            .I(N__66229));
    InMux I__14972 (
            .O(N__66260),
            .I(N__66226));
    InMux I__14971 (
            .O(N__66259),
            .I(N__66221));
    InMux I__14970 (
            .O(N__66256),
            .I(N__66221));
    Span4Mux_v I__14969 (
            .O(N__66253),
            .I(N__66214));
    Span4Mux_v I__14968 (
            .O(N__66250),
            .I(N__66211));
    InMux I__14967 (
            .O(N__66247),
            .I(N__66208));
    Span4Mux_h I__14966 (
            .O(N__66244),
            .I(N__66201));
    Span4Mux_v I__14965 (
            .O(N__66235),
            .I(N__66201));
    LocalMux I__14964 (
            .O(N__66232),
            .I(N__66201));
    InMux I__14963 (
            .O(N__66229),
            .I(N__66198));
    LocalMux I__14962 (
            .O(N__66226),
            .I(N__66193));
    LocalMux I__14961 (
            .O(N__66221),
            .I(N__66193));
    CascadeMux I__14960 (
            .O(N__66220),
            .I(N__66189));
    CascadeMux I__14959 (
            .O(N__66219),
            .I(N__66185));
    CascadeMux I__14958 (
            .O(N__66218),
            .I(N__66181));
    CascadeMux I__14957 (
            .O(N__66217),
            .I(N__66177));
    Span4Mux_h I__14956 (
            .O(N__66214),
            .I(N__66174));
    Span4Mux_v I__14955 (
            .O(N__66211),
            .I(N__66169));
    LocalMux I__14954 (
            .O(N__66208),
            .I(N__66169));
    Span4Mux_v I__14953 (
            .O(N__66201),
            .I(N__66166));
    LocalMux I__14952 (
            .O(N__66198),
            .I(N__66163));
    Span4Mux_v I__14951 (
            .O(N__66193),
            .I(N__66160));
    InMux I__14950 (
            .O(N__66192),
            .I(N__66143));
    InMux I__14949 (
            .O(N__66189),
            .I(N__66143));
    InMux I__14948 (
            .O(N__66188),
            .I(N__66143));
    InMux I__14947 (
            .O(N__66185),
            .I(N__66143));
    InMux I__14946 (
            .O(N__66184),
            .I(N__66143));
    InMux I__14945 (
            .O(N__66181),
            .I(N__66143));
    InMux I__14944 (
            .O(N__66180),
            .I(N__66143));
    InMux I__14943 (
            .O(N__66177),
            .I(N__66143));
    Span4Mux_v I__14942 (
            .O(N__66174),
            .I(N__66140));
    Span4Mux_v I__14941 (
            .O(N__66169),
            .I(N__66137));
    Span4Mux_h I__14940 (
            .O(N__66166),
            .I(N__66132));
    Span4Mux_h I__14939 (
            .O(N__66163),
            .I(N__66132));
    Sp12to4 I__14938 (
            .O(N__66160),
            .I(N__66127));
    LocalMux I__14937 (
            .O(N__66143),
            .I(N__66127));
    Odrv4 I__14936 (
            .O(N__66140),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ));
    Odrv4 I__14935 (
            .O(N__66137),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ));
    Odrv4 I__14934 (
            .O(N__66132),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ));
    Odrv12 I__14933 (
            .O(N__66127),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ));
    InMux I__14932 (
            .O(N__66118),
            .I(N__66115));
    LocalMux I__14931 (
            .O(N__66115),
            .I(N__66112));
    Odrv4 I__14930 (
            .O(N__66112),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n513 ));
    InMux I__14929 (
            .O(N__66109),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18272 ));
    InMux I__14928 (
            .O(N__66106),
            .I(N__66103));
    LocalMux I__14927 (
            .O(N__66103),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n516 ));
    CascadeMux I__14926 (
            .O(N__66100),
            .I(N__66095));
    CascadeMux I__14925 (
            .O(N__66099),
            .I(N__66087));
    CascadeMux I__14924 (
            .O(N__66098),
            .I(N__66083));
    InMux I__14923 (
            .O(N__66095),
            .I(N__66080));
    CascadeMux I__14922 (
            .O(N__66094),
            .I(N__66077));
    CascadeMux I__14921 (
            .O(N__66093),
            .I(N__66074));
    CascadeMux I__14920 (
            .O(N__66092),
            .I(N__66071));
    CascadeMux I__14919 (
            .O(N__66091),
            .I(N__66067));
    CascadeMux I__14918 (
            .O(N__66090),
            .I(N__66064));
    InMux I__14917 (
            .O(N__66087),
            .I(N__66060));
    CascadeMux I__14916 (
            .O(N__66086),
            .I(N__66057));
    InMux I__14915 (
            .O(N__66083),
            .I(N__66053));
    LocalMux I__14914 (
            .O(N__66080),
            .I(N__66050));
    InMux I__14913 (
            .O(N__66077),
            .I(N__66047));
    InMux I__14912 (
            .O(N__66074),
            .I(N__66044));
    InMux I__14911 (
            .O(N__66071),
            .I(N__66041));
    CascadeMux I__14910 (
            .O(N__66070),
            .I(N__66037));
    InMux I__14909 (
            .O(N__66067),
            .I(N__66033));
    InMux I__14908 (
            .O(N__66064),
            .I(N__66025));
    CascadeMux I__14907 (
            .O(N__66063),
            .I(N__66022));
    LocalMux I__14906 (
            .O(N__66060),
            .I(N__66019));
    InMux I__14905 (
            .O(N__66057),
            .I(N__66016));
    InMux I__14904 (
            .O(N__66056),
            .I(N__66013));
    LocalMux I__14903 (
            .O(N__66053),
            .I(N__66005));
    Span4Mux_v I__14902 (
            .O(N__66050),
            .I(N__66005));
    LocalMux I__14901 (
            .O(N__66047),
            .I(N__66005));
    LocalMux I__14900 (
            .O(N__66044),
            .I(N__66002));
    LocalMux I__14899 (
            .O(N__66041),
            .I(N__65999));
    InMux I__14898 (
            .O(N__66040),
            .I(N__65996));
    InMux I__14897 (
            .O(N__66037),
            .I(N__65993));
    CascadeMux I__14896 (
            .O(N__66036),
            .I(N__65990));
    LocalMux I__14895 (
            .O(N__66033),
            .I(N__65987));
    CascadeMux I__14894 (
            .O(N__66032),
            .I(N__65984));
    CascadeMux I__14893 (
            .O(N__66031),
            .I(N__65980));
    CascadeMux I__14892 (
            .O(N__66030),
            .I(N__65976));
    CascadeMux I__14891 (
            .O(N__66029),
            .I(N__65972));
    CascadeMux I__14890 (
            .O(N__66028),
            .I(N__65969));
    LocalMux I__14889 (
            .O(N__66025),
            .I(N__65966));
    InMux I__14888 (
            .O(N__66022),
            .I(N__65963));
    Span4Mux_h I__14887 (
            .O(N__66019),
            .I(N__65958));
    LocalMux I__14886 (
            .O(N__66016),
            .I(N__65958));
    LocalMux I__14885 (
            .O(N__66013),
            .I(N__65955));
    CascadeMux I__14884 (
            .O(N__66012),
            .I(N__65952));
    Span4Mux_h I__14883 (
            .O(N__66005),
            .I(N__65941));
    Span4Mux_h I__14882 (
            .O(N__66002),
            .I(N__65941));
    Span4Mux_h I__14881 (
            .O(N__65999),
            .I(N__65941));
    LocalMux I__14880 (
            .O(N__65996),
            .I(N__65941));
    LocalMux I__14879 (
            .O(N__65993),
            .I(N__65941));
    InMux I__14878 (
            .O(N__65990),
            .I(N__65938));
    Span4Mux_v I__14877 (
            .O(N__65987),
            .I(N__65935));
    InMux I__14876 (
            .O(N__65984),
            .I(N__65928));
    InMux I__14875 (
            .O(N__65983),
            .I(N__65928));
    InMux I__14874 (
            .O(N__65980),
            .I(N__65928));
    InMux I__14873 (
            .O(N__65979),
            .I(N__65917));
    InMux I__14872 (
            .O(N__65976),
            .I(N__65917));
    InMux I__14871 (
            .O(N__65975),
            .I(N__65917));
    InMux I__14870 (
            .O(N__65972),
            .I(N__65917));
    InMux I__14869 (
            .O(N__65969),
            .I(N__65917));
    Span4Mux_h I__14868 (
            .O(N__65966),
            .I(N__65914));
    LocalMux I__14867 (
            .O(N__65963),
            .I(N__65911));
    Sp12to4 I__14866 (
            .O(N__65958),
            .I(N__65908));
    Span4Mux_v I__14865 (
            .O(N__65955),
            .I(N__65905));
    InMux I__14864 (
            .O(N__65952),
            .I(N__65902));
    Span4Mux_v I__14863 (
            .O(N__65941),
            .I(N__65897));
    LocalMux I__14862 (
            .O(N__65938),
            .I(N__65897));
    Span4Mux_h I__14861 (
            .O(N__65935),
            .I(N__65890));
    LocalMux I__14860 (
            .O(N__65928),
            .I(N__65890));
    LocalMux I__14859 (
            .O(N__65917),
            .I(N__65890));
    Span4Mux_v I__14858 (
            .O(N__65914),
            .I(N__65887));
    Span4Mux_v I__14857 (
            .O(N__65911),
            .I(N__65884));
    Span12Mux_s10_v I__14856 (
            .O(N__65908),
            .I(N__65877));
    Sp12to4 I__14855 (
            .O(N__65905),
            .I(N__65877));
    LocalMux I__14854 (
            .O(N__65902),
            .I(N__65877));
    Span4Mux_h I__14853 (
            .O(N__65897),
            .I(N__65872));
    Span4Mux_h I__14852 (
            .O(N__65890),
            .I(N__65872));
    Odrv4 I__14851 (
            .O(N__65887),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ));
    Odrv4 I__14850 (
            .O(N__65884),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ));
    Odrv12 I__14849 (
            .O(N__65877),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ));
    Odrv4 I__14848 (
            .O(N__65872),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ));
    InMux I__14847 (
            .O(N__65863),
            .I(N__65860));
    LocalMux I__14846 (
            .O(N__65860),
            .I(N__65857));
    Odrv12 I__14845 (
            .O(N__65857),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n562 ));
    InMux I__14844 (
            .O(N__65854),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18273 ));
    InMux I__14843 (
            .O(N__65851),
            .I(N__65848));
    LocalMux I__14842 (
            .O(N__65848),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n565 ));
    CascadeMux I__14841 (
            .O(N__65845),
            .I(N__65840));
    CascadeMux I__14840 (
            .O(N__65844),
            .I(N__65836));
    CascadeMux I__14839 (
            .O(N__65843),
            .I(N__65833));
    InMux I__14838 (
            .O(N__65840),
            .I(N__65825));
    CascadeMux I__14837 (
            .O(N__65839),
            .I(N__65822));
    InMux I__14836 (
            .O(N__65836),
            .I(N__65819));
    InMux I__14835 (
            .O(N__65833),
            .I(N__65816));
    CascadeMux I__14834 (
            .O(N__65832),
            .I(N__65813));
    CascadeMux I__14833 (
            .O(N__65831),
            .I(N__65810));
    CascadeMux I__14832 (
            .O(N__65830),
            .I(N__65804));
    CascadeMux I__14831 (
            .O(N__65829),
            .I(N__65801));
    CascadeMux I__14830 (
            .O(N__65828),
            .I(N__65798));
    LocalMux I__14829 (
            .O(N__65825),
            .I(N__65795));
    InMux I__14828 (
            .O(N__65822),
            .I(N__65792));
    LocalMux I__14827 (
            .O(N__65819),
            .I(N__65786));
    LocalMux I__14826 (
            .O(N__65816),
            .I(N__65786));
    InMux I__14825 (
            .O(N__65813),
            .I(N__65783));
    InMux I__14824 (
            .O(N__65810),
            .I(N__65780));
    CascadeMux I__14823 (
            .O(N__65809),
            .I(N__65777));
    CascadeMux I__14822 (
            .O(N__65808),
            .I(N__65773));
    CascadeMux I__14821 (
            .O(N__65807),
            .I(N__65770));
    InMux I__14820 (
            .O(N__65804),
            .I(N__65767));
    InMux I__14819 (
            .O(N__65801),
            .I(N__65764));
    InMux I__14818 (
            .O(N__65798),
            .I(N__65761));
    Span4Mux_v I__14817 (
            .O(N__65795),
            .I(N__65756));
    LocalMux I__14816 (
            .O(N__65792),
            .I(N__65756));
    CascadeMux I__14815 (
            .O(N__65791),
            .I(N__65753));
    Span4Mux_v I__14814 (
            .O(N__65786),
            .I(N__65746));
    LocalMux I__14813 (
            .O(N__65783),
            .I(N__65746));
    LocalMux I__14812 (
            .O(N__65780),
            .I(N__65746));
    InMux I__14811 (
            .O(N__65777),
            .I(N__65743));
    CascadeMux I__14810 (
            .O(N__65776),
            .I(N__65740));
    InMux I__14809 (
            .O(N__65773),
            .I(N__65731));
    InMux I__14808 (
            .O(N__65770),
            .I(N__65728));
    LocalMux I__14807 (
            .O(N__65767),
            .I(N__65725));
    LocalMux I__14806 (
            .O(N__65764),
            .I(N__65718));
    LocalMux I__14805 (
            .O(N__65761),
            .I(N__65718));
    Span4Mux_h I__14804 (
            .O(N__65756),
            .I(N__65718));
    InMux I__14803 (
            .O(N__65753),
            .I(N__65715));
    Span4Mux_h I__14802 (
            .O(N__65746),
            .I(N__65710));
    LocalMux I__14801 (
            .O(N__65743),
            .I(N__65710));
    InMux I__14800 (
            .O(N__65740),
            .I(N__65707));
    InMux I__14799 (
            .O(N__65739),
            .I(N__65704));
    CascadeMux I__14798 (
            .O(N__65738),
            .I(N__65701));
    CascadeMux I__14797 (
            .O(N__65737),
            .I(N__65698));
    CascadeMux I__14796 (
            .O(N__65736),
            .I(N__65694));
    CascadeMux I__14795 (
            .O(N__65735),
            .I(N__65691));
    CascadeMux I__14794 (
            .O(N__65734),
            .I(N__65688));
    LocalMux I__14793 (
            .O(N__65731),
            .I(N__65683));
    LocalMux I__14792 (
            .O(N__65728),
            .I(N__65683));
    Span4Mux_h I__14791 (
            .O(N__65725),
            .I(N__65680));
    Span4Mux_v I__14790 (
            .O(N__65718),
            .I(N__65675));
    LocalMux I__14789 (
            .O(N__65715),
            .I(N__65675));
    Span4Mux_v I__14788 (
            .O(N__65710),
            .I(N__65670));
    LocalMux I__14787 (
            .O(N__65707),
            .I(N__65670));
    LocalMux I__14786 (
            .O(N__65704),
            .I(N__65667));
    InMux I__14785 (
            .O(N__65701),
            .I(N__65662));
    InMux I__14784 (
            .O(N__65698),
            .I(N__65662));
    InMux I__14783 (
            .O(N__65697),
            .I(N__65653));
    InMux I__14782 (
            .O(N__65694),
            .I(N__65653));
    InMux I__14781 (
            .O(N__65691),
            .I(N__65653));
    InMux I__14780 (
            .O(N__65688),
            .I(N__65653));
    Span4Mux_v I__14779 (
            .O(N__65683),
            .I(N__65648));
    Span4Mux_h I__14778 (
            .O(N__65680),
            .I(N__65648));
    Span4Mux_h I__14777 (
            .O(N__65675),
            .I(N__65645));
    Span4Mux_v I__14776 (
            .O(N__65670),
            .I(N__65636));
    Span4Mux_h I__14775 (
            .O(N__65667),
            .I(N__65636));
    LocalMux I__14774 (
            .O(N__65662),
            .I(N__65636));
    LocalMux I__14773 (
            .O(N__65653),
            .I(N__65636));
    Odrv4 I__14772 (
            .O(N__65648),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n135 ));
    Odrv4 I__14771 (
            .O(N__65645),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n135 ));
    Odrv4 I__14770 (
            .O(N__65636),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n135 ));
    InMux I__14769 (
            .O(N__65629),
            .I(N__65626));
    LocalMux I__14768 (
            .O(N__65626),
            .I(N__65623));
    Odrv4 I__14767 (
            .O(N__65623),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n611 ));
    InMux I__14766 (
            .O(N__65620),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18274 ));
    InMux I__14765 (
            .O(N__65617),
            .I(N__65614));
    LocalMux I__14764 (
            .O(N__65614),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n614 ));
    CascadeMux I__14763 (
            .O(N__65611),
            .I(N__65606));
    CascadeMux I__14762 (
            .O(N__65610),
            .I(N__65603));
    CascadeMux I__14761 (
            .O(N__65609),
            .I(N__65597));
    InMux I__14760 (
            .O(N__65606),
            .I(N__65592));
    InMux I__14759 (
            .O(N__65603),
            .I(N__65589));
    CascadeMux I__14758 (
            .O(N__65602),
            .I(N__65586));
    CascadeMux I__14757 (
            .O(N__65601),
            .I(N__65583));
    CascadeMux I__14756 (
            .O(N__65600),
            .I(N__65577));
    InMux I__14755 (
            .O(N__65597),
            .I(N__65574));
    CascadeMux I__14754 (
            .O(N__65596),
            .I(N__65571));
    InMux I__14753 (
            .O(N__65595),
            .I(N__65567));
    LocalMux I__14752 (
            .O(N__65592),
            .I(N__65562));
    LocalMux I__14751 (
            .O(N__65589),
            .I(N__65562));
    InMux I__14750 (
            .O(N__65586),
            .I(N__65559));
    InMux I__14749 (
            .O(N__65583),
            .I(N__65556));
    CascadeMux I__14748 (
            .O(N__65582),
            .I(N__65553));
    CascadeMux I__14747 (
            .O(N__65581),
            .I(N__65550));
    CascadeMux I__14746 (
            .O(N__65580),
            .I(N__65547));
    InMux I__14745 (
            .O(N__65577),
            .I(N__65543));
    LocalMux I__14744 (
            .O(N__65574),
            .I(N__65540));
    InMux I__14743 (
            .O(N__65571),
            .I(N__65537));
    CascadeMux I__14742 (
            .O(N__65570),
            .I(N__65534));
    LocalMux I__14741 (
            .O(N__65567),
            .I(N__65531));
    Span4Mux_v I__14740 (
            .O(N__65562),
            .I(N__65524));
    LocalMux I__14739 (
            .O(N__65559),
            .I(N__65524));
    LocalMux I__14738 (
            .O(N__65556),
            .I(N__65524));
    InMux I__14737 (
            .O(N__65553),
            .I(N__65521));
    InMux I__14736 (
            .O(N__65550),
            .I(N__65518));
    InMux I__14735 (
            .O(N__65547),
            .I(N__65515));
    CascadeMux I__14734 (
            .O(N__65546),
            .I(N__65512));
    LocalMux I__14733 (
            .O(N__65543),
            .I(N__65504));
    Span4Mux_h I__14732 (
            .O(N__65540),
            .I(N__65499));
    LocalMux I__14731 (
            .O(N__65537),
            .I(N__65499));
    InMux I__14730 (
            .O(N__65534),
            .I(N__65496));
    Span4Mux_v I__14729 (
            .O(N__65531),
            .I(N__65493));
    Span4Mux_h I__14728 (
            .O(N__65524),
            .I(N__65483));
    LocalMux I__14727 (
            .O(N__65521),
            .I(N__65483));
    LocalMux I__14726 (
            .O(N__65518),
            .I(N__65483));
    LocalMux I__14725 (
            .O(N__65515),
            .I(N__65483));
    InMux I__14724 (
            .O(N__65512),
            .I(N__65480));
    InMux I__14723 (
            .O(N__65511),
            .I(N__65477));
    InMux I__14722 (
            .O(N__65510),
            .I(N__65468));
    InMux I__14721 (
            .O(N__65509),
            .I(N__65468));
    InMux I__14720 (
            .O(N__65508),
            .I(N__65468));
    InMux I__14719 (
            .O(N__65507),
            .I(N__65468));
    Span4Mux_h I__14718 (
            .O(N__65504),
            .I(N__65464));
    Span4Mux_v I__14717 (
            .O(N__65499),
            .I(N__65459));
    LocalMux I__14716 (
            .O(N__65496),
            .I(N__65459));
    Span4Mux_h I__14715 (
            .O(N__65493),
            .I(N__65456));
    InMux I__14714 (
            .O(N__65492),
            .I(N__65453));
    Span4Mux_v I__14713 (
            .O(N__65483),
            .I(N__65448));
    LocalMux I__14712 (
            .O(N__65480),
            .I(N__65448));
    LocalMux I__14711 (
            .O(N__65477),
            .I(N__65445));
    LocalMux I__14710 (
            .O(N__65468),
            .I(N__65442));
    InMux I__14709 (
            .O(N__65467),
            .I(N__65439));
    Span4Mux_v I__14708 (
            .O(N__65464),
            .I(N__65432));
    Span4Mux_h I__14707 (
            .O(N__65459),
            .I(N__65432));
    Sp12to4 I__14706 (
            .O(N__65456),
            .I(N__65427));
    LocalMux I__14705 (
            .O(N__65453),
            .I(N__65427));
    Span4Mux_v I__14704 (
            .O(N__65448),
            .I(N__65418));
    Span4Mux_v I__14703 (
            .O(N__65445),
            .I(N__65418));
    Span4Mux_v I__14702 (
            .O(N__65442),
            .I(N__65418));
    LocalMux I__14701 (
            .O(N__65439),
            .I(N__65418));
    InMux I__14700 (
            .O(N__65438),
            .I(N__65413));
    InMux I__14699 (
            .O(N__65437),
            .I(N__65413));
    Odrv4 I__14698 (
            .O(N__65432),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ));
    Odrv12 I__14697 (
            .O(N__65427),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ));
    Odrv4 I__14696 (
            .O(N__65418),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ));
    LocalMux I__14695 (
            .O(N__65413),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ));
    CascadeMux I__14694 (
            .O(N__65404),
            .I(N__65401));
    InMux I__14693 (
            .O(N__65401),
            .I(N__65398));
    LocalMux I__14692 (
            .O(N__65398),
            .I(N__65395));
    Odrv4 I__14691 (
            .O(N__65395),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n660 ));
    InMux I__14690 (
            .O(N__65392),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18275 ));
    InMux I__14689 (
            .O(N__65389),
            .I(N__65381));
    InMux I__14688 (
            .O(N__65388),
            .I(N__65378));
    InMux I__14687 (
            .O(N__65387),
            .I(N__65375));
    CascadeMux I__14686 (
            .O(N__65386),
            .I(N__65371));
    InMux I__14685 (
            .O(N__65385),
            .I(N__65368));
    InMux I__14684 (
            .O(N__65384),
            .I(N__65365));
    LocalMux I__14683 (
            .O(N__65381),
            .I(N__65362));
    LocalMux I__14682 (
            .O(N__65378),
            .I(N__65356));
    LocalMux I__14681 (
            .O(N__65375),
            .I(N__65356));
    InMux I__14680 (
            .O(N__65374),
            .I(N__65353));
    InMux I__14679 (
            .O(N__65371),
            .I(N__65349));
    LocalMux I__14678 (
            .O(N__65368),
            .I(N__65343));
    LocalMux I__14677 (
            .O(N__65365),
            .I(N__65343));
    Span4Mux_v I__14676 (
            .O(N__65362),
            .I(N__65338));
    InMux I__14675 (
            .O(N__65361),
            .I(N__65335));
    Span4Mux_h I__14674 (
            .O(N__65356),
            .I(N__65330));
    LocalMux I__14673 (
            .O(N__65353),
            .I(N__65330));
    InMux I__14672 (
            .O(N__65352),
            .I(N__65327));
    LocalMux I__14671 (
            .O(N__65349),
            .I(N__65324));
    InMux I__14670 (
            .O(N__65348),
            .I(N__65321));
    Span4Mux_h I__14669 (
            .O(N__65343),
            .I(N__65317));
    InMux I__14668 (
            .O(N__65342),
            .I(N__65314));
    InMux I__14667 (
            .O(N__65341),
            .I(N__65310));
    Span4Mux_h I__14666 (
            .O(N__65338),
            .I(N__65301));
    LocalMux I__14665 (
            .O(N__65335),
            .I(N__65301));
    Span4Mux_h I__14664 (
            .O(N__65330),
            .I(N__65301));
    LocalMux I__14663 (
            .O(N__65327),
            .I(N__65301));
    Span4Mux_v I__14662 (
            .O(N__65324),
            .I(N__65296));
    LocalMux I__14661 (
            .O(N__65321),
            .I(N__65296));
    InMux I__14660 (
            .O(N__65320),
            .I(N__65293));
    Span4Mux_v I__14659 (
            .O(N__65317),
            .I(N__65288));
    LocalMux I__14658 (
            .O(N__65314),
            .I(N__65288));
    InMux I__14657 (
            .O(N__65313),
            .I(N__65285));
    LocalMux I__14656 (
            .O(N__65310),
            .I(N__65281));
    Span4Mux_v I__14655 (
            .O(N__65301),
            .I(N__65274));
    Span4Mux_v I__14654 (
            .O(N__65296),
            .I(N__65274));
    LocalMux I__14653 (
            .O(N__65293),
            .I(N__65274));
    Span4Mux_h I__14652 (
            .O(N__65288),
            .I(N__65271));
    LocalMux I__14651 (
            .O(N__65285),
            .I(N__65268));
    InMux I__14650 (
            .O(N__65284),
            .I(N__65265));
    Span4Mux_h I__14649 (
            .O(N__65281),
            .I(N__65261));
    Span4Mux_h I__14648 (
            .O(N__65274),
            .I(N__65258));
    Span4Mux_h I__14647 (
            .O(N__65271),
            .I(N__65251));
    Span4Mux_v I__14646 (
            .O(N__65268),
            .I(N__65251));
    LocalMux I__14645 (
            .O(N__65265),
            .I(N__65251));
    CascadeMux I__14644 (
            .O(N__65264),
            .I(N__65248));
    Sp12to4 I__14643 (
            .O(N__65261),
            .I(N__65245));
    Span4Mux_v I__14642 (
            .O(N__65258),
            .I(N__65242));
    Span4Mux_h I__14641 (
            .O(N__65251),
            .I(N__65239));
    InMux I__14640 (
            .O(N__65248),
            .I(N__65236));
    Odrv12 I__14639 (
            .O(N__65245),
            .I(n141_adj_2421));
    Odrv4 I__14638 (
            .O(N__65242),
            .I(n141_adj_2421));
    Odrv4 I__14637 (
            .O(N__65239),
            .I(n141_adj_2421));
    LocalMux I__14636 (
            .O(N__65236),
            .I(n141_adj_2421));
    CascadeMux I__14635 (
            .O(N__65227),
            .I(N__65224));
    InMux I__14634 (
            .O(N__65224),
            .I(N__65221));
    LocalMux I__14633 (
            .O(N__65221),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n663 ));
    CascadeMux I__14632 (
            .O(N__65218),
            .I(N__65215));
    InMux I__14631 (
            .O(N__65215),
            .I(N__65212));
    LocalMux I__14630 (
            .O(N__65212),
            .I(N__65209));
    Odrv12 I__14629 (
            .O(N__65209),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n709 ));
    InMux I__14628 (
            .O(N__65206),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18276 ));
    InMux I__14627 (
            .O(N__65203),
            .I(N__65198));
    InMux I__14626 (
            .O(N__65202),
            .I(N__65195));
    InMux I__14625 (
            .O(N__65201),
            .I(N__65189));
    LocalMux I__14624 (
            .O(N__65198),
            .I(N__65185));
    LocalMux I__14623 (
            .O(N__65195),
            .I(N__65182));
    InMux I__14622 (
            .O(N__65194),
            .I(N__65179));
    InMux I__14621 (
            .O(N__65193),
            .I(N__65175));
    InMux I__14620 (
            .O(N__65192),
            .I(N__65172));
    LocalMux I__14619 (
            .O(N__65189),
            .I(N__65166));
    CascadeMux I__14618 (
            .O(N__65188),
            .I(N__65163));
    Span4Mux_v I__14617 (
            .O(N__65185),
            .I(N__65156));
    Span4Mux_h I__14616 (
            .O(N__65182),
            .I(N__65156));
    LocalMux I__14615 (
            .O(N__65179),
            .I(N__65156));
    CascadeMux I__14614 (
            .O(N__65178),
            .I(N__65153));
    LocalMux I__14613 (
            .O(N__65175),
            .I(N__65149));
    LocalMux I__14612 (
            .O(N__65172),
            .I(N__65146));
    InMux I__14611 (
            .O(N__65171),
            .I(N__65143));
    InMux I__14610 (
            .O(N__65170),
            .I(N__65140));
    CascadeMux I__14609 (
            .O(N__65169),
            .I(N__65136));
    Span4Mux_v I__14608 (
            .O(N__65166),
            .I(N__65132));
    InMux I__14607 (
            .O(N__65163),
            .I(N__65129));
    Span4Mux_v I__14606 (
            .O(N__65156),
            .I(N__65126));
    InMux I__14605 (
            .O(N__65153),
            .I(N__65123));
    CascadeMux I__14604 (
            .O(N__65152),
            .I(N__65120));
    Span4Mux_h I__14603 (
            .O(N__65149),
            .I(N__65109));
    Span4Mux_v I__14602 (
            .O(N__65146),
            .I(N__65109));
    LocalMux I__14601 (
            .O(N__65143),
            .I(N__65109));
    LocalMux I__14600 (
            .O(N__65140),
            .I(N__65109));
    InMux I__14599 (
            .O(N__65139),
            .I(N__65106));
    InMux I__14598 (
            .O(N__65136),
            .I(N__65103));
    InMux I__14597 (
            .O(N__65135),
            .I(N__65100));
    Span4Mux_h I__14596 (
            .O(N__65132),
            .I(N__65095));
    LocalMux I__14595 (
            .O(N__65129),
            .I(N__65095));
    Span4Mux_h I__14594 (
            .O(N__65126),
            .I(N__65090));
    LocalMux I__14593 (
            .O(N__65123),
            .I(N__65090));
    InMux I__14592 (
            .O(N__65120),
            .I(N__65087));
    InMux I__14591 (
            .O(N__65119),
            .I(N__65082));
    InMux I__14590 (
            .O(N__65118),
            .I(N__65082));
    Span4Mux_v I__14589 (
            .O(N__65109),
            .I(N__65077));
    LocalMux I__14588 (
            .O(N__65106),
            .I(N__65077));
    LocalMux I__14587 (
            .O(N__65103),
            .I(N__65072));
    LocalMux I__14586 (
            .O(N__65100),
            .I(N__65072));
    Span4Mux_v I__14585 (
            .O(N__65095),
            .I(N__65065));
    Span4Mux_h I__14584 (
            .O(N__65090),
            .I(N__65065));
    LocalMux I__14583 (
            .O(N__65087),
            .I(N__65065));
    LocalMux I__14582 (
            .O(N__65082),
            .I(N__65062));
    Span4Mux_v I__14581 (
            .O(N__65077),
            .I(N__65058));
    Span12Mux_v I__14580 (
            .O(N__65072),
            .I(N__65055));
    Span4Mux_v I__14579 (
            .O(N__65065),
            .I(N__65050));
    Span4Mux_h I__14578 (
            .O(N__65062),
            .I(N__65050));
    InMux I__14577 (
            .O(N__65061),
            .I(N__65047));
    Odrv4 I__14576 (
            .O(N__65058),
            .I(n146_adj_2423));
    Odrv12 I__14575 (
            .O(N__65055),
            .I(n146_adj_2423));
    Odrv4 I__14574 (
            .O(N__65050),
            .I(n146_adj_2423));
    LocalMux I__14573 (
            .O(N__65047),
            .I(n146_adj_2423));
    CascadeMux I__14572 (
            .O(N__65038),
            .I(N__65035));
    InMux I__14571 (
            .O(N__65035),
            .I(N__65032));
    LocalMux I__14570 (
            .O(N__65032),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n712 ));
    InMux I__14569 (
            .O(N__65029),
            .I(N__65026));
    LocalMux I__14568 (
            .O(N__65026),
            .I(N__65023));
    Span12Mux_h I__14567 (
            .O(N__65023),
            .I(N__65020));
    Odrv12 I__14566 (
            .O(N__65020),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n766 ));
    CascadeMux I__14565 (
            .O(N__65017),
            .I(N__65001));
    CascadeMux I__14564 (
            .O(N__65016),
            .I(N__64998));
    CascadeMux I__14563 (
            .O(N__65015),
            .I(N__64995));
    CascadeMux I__14562 (
            .O(N__65014),
            .I(N__64992));
    CascadeMux I__14561 (
            .O(N__65013),
            .I(N__64989));
    CascadeMux I__14560 (
            .O(N__65012),
            .I(N__64986));
    CascadeMux I__14559 (
            .O(N__65011),
            .I(N__64983));
    CascadeMux I__14558 (
            .O(N__65010),
            .I(N__64980));
    CascadeMux I__14557 (
            .O(N__65009),
            .I(N__64977));
    CascadeMux I__14556 (
            .O(N__65008),
            .I(N__64974));
    CascadeMux I__14555 (
            .O(N__65007),
            .I(N__64971));
    CascadeMux I__14554 (
            .O(N__65006),
            .I(N__64968));
    CascadeMux I__14553 (
            .O(N__65005),
            .I(N__64965));
    CascadeMux I__14552 (
            .O(N__65004),
            .I(N__64961));
    InMux I__14551 (
            .O(N__65001),
            .I(N__64957));
    InMux I__14550 (
            .O(N__64998),
            .I(N__64948));
    InMux I__14549 (
            .O(N__64995),
            .I(N__64948));
    InMux I__14548 (
            .O(N__64992),
            .I(N__64948));
    InMux I__14547 (
            .O(N__64989),
            .I(N__64940));
    InMux I__14546 (
            .O(N__64986),
            .I(N__64940));
    InMux I__14545 (
            .O(N__64983),
            .I(N__64940));
    InMux I__14544 (
            .O(N__64980),
            .I(N__64933));
    InMux I__14543 (
            .O(N__64977),
            .I(N__64933));
    InMux I__14542 (
            .O(N__64974),
            .I(N__64933));
    InMux I__14541 (
            .O(N__64971),
            .I(N__64922));
    InMux I__14540 (
            .O(N__64968),
            .I(N__64922));
    InMux I__14539 (
            .O(N__64965),
            .I(N__64922));
    InMux I__14538 (
            .O(N__64964),
            .I(N__64922));
    InMux I__14537 (
            .O(N__64961),
            .I(N__64922));
    InMux I__14536 (
            .O(N__64960),
            .I(N__64918));
    LocalMux I__14535 (
            .O(N__64957),
            .I(N__64915));
    InMux I__14534 (
            .O(N__64956),
            .I(N__64911));
    CascadeMux I__14533 (
            .O(N__64955),
            .I(N__64907));
    LocalMux I__14532 (
            .O(N__64948),
            .I(N__64904));
    InMux I__14531 (
            .O(N__64947),
            .I(N__64901));
    LocalMux I__14530 (
            .O(N__64940),
            .I(N__64892));
    LocalMux I__14529 (
            .O(N__64933),
            .I(N__64892));
    LocalMux I__14528 (
            .O(N__64922),
            .I(N__64892));
    InMux I__14527 (
            .O(N__64921),
            .I(N__64889));
    LocalMux I__14526 (
            .O(N__64918),
            .I(N__64884));
    Span4Mux_v I__14525 (
            .O(N__64915),
            .I(N__64881));
    InMux I__14524 (
            .O(N__64914),
            .I(N__64878));
    LocalMux I__14523 (
            .O(N__64911),
            .I(N__64875));
    InMux I__14522 (
            .O(N__64910),
            .I(N__64872));
    InMux I__14521 (
            .O(N__64907),
            .I(N__64869));
    Span4Mux_v I__14520 (
            .O(N__64904),
            .I(N__64864));
    LocalMux I__14519 (
            .O(N__64901),
            .I(N__64864));
    CascadeMux I__14518 (
            .O(N__64900),
            .I(N__64859));
    InMux I__14517 (
            .O(N__64899),
            .I(N__64856));
    Span4Mux_v I__14516 (
            .O(N__64892),
            .I(N__64851));
    LocalMux I__14515 (
            .O(N__64889),
            .I(N__64851));
    InMux I__14514 (
            .O(N__64888),
            .I(N__64848));
    CascadeMux I__14513 (
            .O(N__64887),
            .I(N__64845));
    Span4Mux_v I__14512 (
            .O(N__64884),
            .I(N__64837));
    Span4Mux_h I__14511 (
            .O(N__64881),
            .I(N__64837));
    LocalMux I__14510 (
            .O(N__64878),
            .I(N__64837));
    Span4Mux_v I__14509 (
            .O(N__64875),
            .I(N__64832));
    LocalMux I__14508 (
            .O(N__64872),
            .I(N__64832));
    LocalMux I__14507 (
            .O(N__64869),
            .I(N__64829));
    Span4Mux_v I__14506 (
            .O(N__64864),
            .I(N__64826));
    InMux I__14505 (
            .O(N__64863),
            .I(N__64823));
    InMux I__14504 (
            .O(N__64862),
            .I(N__64820));
    InMux I__14503 (
            .O(N__64859),
            .I(N__64817));
    LocalMux I__14502 (
            .O(N__64856),
            .I(N__64810));
    Span4Mux_h I__14501 (
            .O(N__64851),
            .I(N__64810));
    LocalMux I__14500 (
            .O(N__64848),
            .I(N__64810));
    InMux I__14499 (
            .O(N__64845),
            .I(N__64807));
    CascadeMux I__14498 (
            .O(N__64844),
            .I(N__64804));
    Span4Mux_v I__14497 (
            .O(N__64837),
            .I(N__64801));
    Span4Mux_v I__14496 (
            .O(N__64832),
            .I(N__64798));
    Span4Mux_v I__14495 (
            .O(N__64829),
            .I(N__64787));
    Span4Mux_h I__14494 (
            .O(N__64826),
            .I(N__64787));
    LocalMux I__14493 (
            .O(N__64823),
            .I(N__64787));
    LocalMux I__14492 (
            .O(N__64820),
            .I(N__64787));
    LocalMux I__14491 (
            .O(N__64817),
            .I(N__64787));
    Span4Mux_v I__14490 (
            .O(N__64810),
            .I(N__64782));
    LocalMux I__14489 (
            .O(N__64807),
            .I(N__64782));
    InMux I__14488 (
            .O(N__64804),
            .I(N__64779));
    Span4Mux_v I__14487 (
            .O(N__64801),
            .I(N__64776));
    Span4Mux_h I__14486 (
            .O(N__64798),
            .I(N__64771));
    Span4Mux_v I__14485 (
            .O(N__64787),
            .I(N__64771));
    Span4Mux_v I__14484 (
            .O(N__64782),
            .I(N__64766));
    LocalMux I__14483 (
            .O(N__64779),
            .I(N__64766));
    Odrv4 I__14482 (
            .O(N__64776),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n102 ));
    Odrv4 I__14481 (
            .O(N__64771),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n102 ));
    Odrv4 I__14480 (
            .O(N__64766),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n102 ));
    CascadeMux I__14479 (
            .O(N__64759),
            .I(N__64755));
    CascadeMux I__14478 (
            .O(N__64758),
            .I(N__64750));
    InMux I__14477 (
            .O(N__64755),
            .I(N__64744));
    CascadeMux I__14476 (
            .O(N__64754),
            .I(N__64741));
    CascadeMux I__14475 (
            .O(N__64753),
            .I(N__64738));
    InMux I__14474 (
            .O(N__64750),
            .I(N__64735));
    CascadeMux I__14473 (
            .O(N__64749),
            .I(N__64731));
    CascadeMux I__14472 (
            .O(N__64748),
            .I(N__64728));
    InMux I__14471 (
            .O(N__64747),
            .I(N__64723));
    LocalMux I__14470 (
            .O(N__64744),
            .I(N__64720));
    InMux I__14469 (
            .O(N__64741),
            .I(N__64717));
    InMux I__14468 (
            .O(N__64738),
            .I(N__64714));
    LocalMux I__14467 (
            .O(N__64735),
            .I(N__64709));
    CascadeMux I__14466 (
            .O(N__64734),
            .I(N__64706));
    InMux I__14465 (
            .O(N__64731),
            .I(N__64703));
    InMux I__14464 (
            .O(N__64728),
            .I(N__64700));
    CascadeMux I__14463 (
            .O(N__64727),
            .I(N__64697));
    CascadeMux I__14462 (
            .O(N__64726),
            .I(N__64694));
    LocalMux I__14461 (
            .O(N__64723),
            .I(N__64690));
    Span4Mux_v I__14460 (
            .O(N__64720),
            .I(N__64683));
    LocalMux I__14459 (
            .O(N__64717),
            .I(N__64683));
    LocalMux I__14458 (
            .O(N__64714),
            .I(N__64683));
    InMux I__14457 (
            .O(N__64713),
            .I(N__64680));
    InMux I__14456 (
            .O(N__64712),
            .I(N__64677));
    Span4Mux_v I__14455 (
            .O(N__64709),
            .I(N__64674));
    InMux I__14454 (
            .O(N__64706),
            .I(N__64671));
    LocalMux I__14453 (
            .O(N__64703),
            .I(N__64666));
    LocalMux I__14452 (
            .O(N__64700),
            .I(N__64666));
    InMux I__14451 (
            .O(N__64697),
            .I(N__64663));
    InMux I__14450 (
            .O(N__64694),
            .I(N__64660));
    CascadeMux I__14449 (
            .O(N__64693),
            .I(N__64657));
    Span4Mux_v I__14448 (
            .O(N__64690),
            .I(N__64648));
    Span4Mux_h I__14447 (
            .O(N__64683),
            .I(N__64648));
    LocalMux I__14446 (
            .O(N__64680),
            .I(N__64648));
    LocalMux I__14445 (
            .O(N__64677),
            .I(N__64648));
    Span4Mux_h I__14444 (
            .O(N__64674),
            .I(N__64633));
    LocalMux I__14443 (
            .O(N__64671),
            .I(N__64633));
    Span4Mux_v I__14442 (
            .O(N__64666),
            .I(N__64625));
    LocalMux I__14441 (
            .O(N__64663),
            .I(N__64625));
    LocalMux I__14440 (
            .O(N__64660),
            .I(N__64625));
    InMux I__14439 (
            .O(N__64657),
            .I(N__64622));
    Span4Mux_v I__14438 (
            .O(N__64648),
            .I(N__64619));
    CascadeMux I__14437 (
            .O(N__64647),
            .I(N__64616));
    CascadeMux I__14436 (
            .O(N__64646),
            .I(N__64613));
    CascadeMux I__14435 (
            .O(N__64645),
            .I(N__64609));
    CascadeMux I__14434 (
            .O(N__64644),
            .I(N__64606));
    CascadeMux I__14433 (
            .O(N__64643),
            .I(N__64603));
    CascadeMux I__14432 (
            .O(N__64642),
            .I(N__64600));
    CascadeMux I__14431 (
            .O(N__64641),
            .I(N__64596));
    CascadeMux I__14430 (
            .O(N__64640),
            .I(N__64593));
    CascadeMux I__14429 (
            .O(N__64639),
            .I(N__64589));
    CascadeMux I__14428 (
            .O(N__64638),
            .I(N__64585));
    Span4Mux_v I__14427 (
            .O(N__64633),
            .I(N__64582));
    InMux I__14426 (
            .O(N__64632),
            .I(N__64579));
    Span4Mux_h I__14425 (
            .O(N__64625),
            .I(N__64576));
    LocalMux I__14424 (
            .O(N__64622),
            .I(N__64573));
    Span4Mux_h I__14423 (
            .O(N__64619),
            .I(N__64570));
    InMux I__14422 (
            .O(N__64616),
            .I(N__64565));
    InMux I__14421 (
            .O(N__64613),
            .I(N__64565));
    InMux I__14420 (
            .O(N__64612),
            .I(N__64556));
    InMux I__14419 (
            .O(N__64609),
            .I(N__64556));
    InMux I__14418 (
            .O(N__64606),
            .I(N__64556));
    InMux I__14417 (
            .O(N__64603),
            .I(N__64556));
    InMux I__14416 (
            .O(N__64600),
            .I(N__64549));
    InMux I__14415 (
            .O(N__64599),
            .I(N__64549));
    InMux I__14414 (
            .O(N__64596),
            .I(N__64549));
    InMux I__14413 (
            .O(N__64593),
            .I(N__64538));
    InMux I__14412 (
            .O(N__64592),
            .I(N__64538));
    InMux I__14411 (
            .O(N__64589),
            .I(N__64538));
    InMux I__14410 (
            .O(N__64588),
            .I(N__64538));
    InMux I__14409 (
            .O(N__64585),
            .I(N__64538));
    Sp12to4 I__14408 (
            .O(N__64582),
            .I(N__64533));
    LocalMux I__14407 (
            .O(N__64579),
            .I(N__64533));
    Span4Mux_v I__14406 (
            .O(N__64576),
            .I(N__64528));
    Span4Mux_h I__14405 (
            .O(N__64573),
            .I(N__64528));
    Sp12to4 I__14404 (
            .O(N__64570),
            .I(N__64519));
    LocalMux I__14403 (
            .O(N__64565),
            .I(N__64519));
    LocalMux I__14402 (
            .O(N__64556),
            .I(N__64519));
    LocalMux I__14401 (
            .O(N__64549),
            .I(N__64519));
    LocalMux I__14400 (
            .O(N__64538),
            .I(N__64516));
    Odrv12 I__14399 (
            .O(N__64533),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ));
    Odrv4 I__14398 (
            .O(N__64528),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ));
    Odrv12 I__14397 (
            .O(N__64519),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ));
    Odrv4 I__14396 (
            .O(N__64516),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ));
    InMux I__14395 (
            .O(N__64507),
            .I(N__64504));
    LocalMux I__14394 (
            .O(N__64504),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n75 ));
    CascadeMux I__14393 (
            .O(N__64501),
            .I(N__64498));
    InMux I__14392 (
            .O(N__64498),
            .I(N__64493));
    CascadeMux I__14391 (
            .O(N__64497),
            .I(N__64490));
    CascadeMux I__14390 (
            .O(N__64496),
            .I(N__64485));
    LocalMux I__14389 (
            .O(N__64493),
            .I(N__64482));
    InMux I__14388 (
            .O(N__64490),
            .I(N__64479));
    CascadeMux I__14387 (
            .O(N__64489),
            .I(N__64475));
    CascadeMux I__14386 (
            .O(N__64488),
            .I(N__64472));
    InMux I__14385 (
            .O(N__64485),
            .I(N__64467));
    Span4Mux_h I__14384 (
            .O(N__64482),
            .I(N__64461));
    LocalMux I__14383 (
            .O(N__64479),
            .I(N__64461));
    InMux I__14382 (
            .O(N__64478),
            .I(N__64458));
    InMux I__14381 (
            .O(N__64475),
            .I(N__64455));
    InMux I__14380 (
            .O(N__64472),
            .I(N__64447));
    InMux I__14379 (
            .O(N__64471),
            .I(N__64444));
    CascadeMux I__14378 (
            .O(N__64470),
            .I(N__64441));
    LocalMux I__14377 (
            .O(N__64467),
            .I(N__64434));
    CascadeMux I__14376 (
            .O(N__64466),
            .I(N__64431));
    Span4Mux_v I__14375 (
            .O(N__64461),
            .I(N__64426));
    LocalMux I__14374 (
            .O(N__64458),
            .I(N__64426));
    LocalMux I__14373 (
            .O(N__64455),
            .I(N__64423));
    InMux I__14372 (
            .O(N__64454),
            .I(N__64420));
    InMux I__14371 (
            .O(N__64453),
            .I(N__64417));
    CascadeMux I__14370 (
            .O(N__64452),
            .I(N__64414));
    CascadeMux I__14369 (
            .O(N__64451),
            .I(N__64411));
    CascadeMux I__14368 (
            .O(N__64450),
            .I(N__64408));
    LocalMux I__14367 (
            .O(N__64447),
            .I(N__64403));
    LocalMux I__14366 (
            .O(N__64444),
            .I(N__64403));
    InMux I__14365 (
            .O(N__64441),
            .I(N__64400));
    InMux I__14364 (
            .O(N__64440),
            .I(N__64397));
    CascadeMux I__14363 (
            .O(N__64439),
            .I(N__64393));
    CascadeMux I__14362 (
            .O(N__64438),
            .I(N__64389));
    CascadeMux I__14361 (
            .O(N__64437),
            .I(N__64385));
    Span4Mux_v I__14360 (
            .O(N__64434),
            .I(N__64378));
    InMux I__14359 (
            .O(N__64431),
            .I(N__64375));
    Span4Mux_v I__14358 (
            .O(N__64426),
            .I(N__64368));
    Span4Mux_v I__14357 (
            .O(N__64423),
            .I(N__64368));
    LocalMux I__14356 (
            .O(N__64420),
            .I(N__64368));
    LocalMux I__14355 (
            .O(N__64417),
            .I(N__64365));
    InMux I__14354 (
            .O(N__64414),
            .I(N__64362));
    InMux I__14353 (
            .O(N__64411),
            .I(N__64359));
    InMux I__14352 (
            .O(N__64408),
            .I(N__64356));
    Span4Mux_v I__14351 (
            .O(N__64403),
            .I(N__64349));
    LocalMux I__14350 (
            .O(N__64400),
            .I(N__64349));
    LocalMux I__14349 (
            .O(N__64397),
            .I(N__64349));
    InMux I__14348 (
            .O(N__64396),
            .I(N__64336));
    InMux I__14347 (
            .O(N__64393),
            .I(N__64336));
    InMux I__14346 (
            .O(N__64392),
            .I(N__64336));
    InMux I__14345 (
            .O(N__64389),
            .I(N__64336));
    InMux I__14344 (
            .O(N__64388),
            .I(N__64336));
    InMux I__14343 (
            .O(N__64385),
            .I(N__64336));
    CascadeMux I__14342 (
            .O(N__64384),
            .I(N__64332));
    CascadeMux I__14341 (
            .O(N__64383),
            .I(N__64328));
    CascadeMux I__14340 (
            .O(N__64382),
            .I(N__64324));
    CascadeMux I__14339 (
            .O(N__64381),
            .I(N__64320));
    Span4Mux_h I__14338 (
            .O(N__64378),
            .I(N__64315));
    LocalMux I__14337 (
            .O(N__64375),
            .I(N__64315));
    Span4Mux_h I__14336 (
            .O(N__64368),
            .I(N__64308));
    Span4Mux_h I__14335 (
            .O(N__64365),
            .I(N__64308));
    LocalMux I__14334 (
            .O(N__64362),
            .I(N__64308));
    LocalMux I__14333 (
            .O(N__64359),
            .I(N__64303));
    LocalMux I__14332 (
            .O(N__64356),
            .I(N__64303));
    Span4Mux_h I__14331 (
            .O(N__64349),
            .I(N__64298));
    LocalMux I__14330 (
            .O(N__64336),
            .I(N__64298));
    InMux I__14329 (
            .O(N__64335),
            .I(N__64281));
    InMux I__14328 (
            .O(N__64332),
            .I(N__64281));
    InMux I__14327 (
            .O(N__64331),
            .I(N__64281));
    InMux I__14326 (
            .O(N__64328),
            .I(N__64281));
    InMux I__14325 (
            .O(N__64327),
            .I(N__64281));
    InMux I__14324 (
            .O(N__64324),
            .I(N__64281));
    InMux I__14323 (
            .O(N__64323),
            .I(N__64281));
    InMux I__14322 (
            .O(N__64320),
            .I(N__64281));
    Span4Mux_v I__14321 (
            .O(N__64315),
            .I(N__64278));
    Span4Mux_v I__14320 (
            .O(N__64308),
            .I(N__64275));
    Span12Mux_h I__14319 (
            .O(N__64303),
            .I(N__64268));
    Sp12to4 I__14318 (
            .O(N__64298),
            .I(N__64268));
    LocalMux I__14317 (
            .O(N__64281),
            .I(N__64268));
    Odrv4 I__14316 (
            .O(N__64278),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n105 ));
    Odrv4 I__14315 (
            .O(N__64275),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n105 ));
    Odrv12 I__14314 (
            .O(N__64268),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n105 ));
    InMux I__14313 (
            .O(N__64261),
            .I(N__64258));
    LocalMux I__14312 (
            .O(N__64258),
            .I(N__64255));
    Odrv12 I__14311 (
            .O(N__64255),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n121 ));
    InMux I__14310 (
            .O(N__64252),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18264 ));
    InMux I__14309 (
            .O(N__64249),
            .I(N__64246));
    LocalMux I__14308 (
            .O(N__64246),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n124 ));
    CascadeMux I__14307 (
            .O(N__64243),
            .I(N__64227));
    CascadeMux I__14306 (
            .O(N__64242),
            .I(N__64224));
    CascadeMux I__14305 (
            .O(N__64241),
            .I(N__64221));
    CascadeMux I__14304 (
            .O(N__64240),
            .I(N__64216));
    CascadeMux I__14303 (
            .O(N__64239),
            .I(N__64212));
    CascadeMux I__14302 (
            .O(N__64238),
            .I(N__64208));
    CascadeMux I__14301 (
            .O(N__64237),
            .I(N__64204));
    CascadeMux I__14300 (
            .O(N__64236),
            .I(N__64201));
    CascadeMux I__14299 (
            .O(N__64235),
            .I(N__64197));
    CascadeMux I__14298 (
            .O(N__64234),
            .I(N__64193));
    CascadeMux I__14297 (
            .O(N__64233),
            .I(N__64189));
    CascadeMux I__14296 (
            .O(N__64232),
            .I(N__64186));
    CascadeMux I__14295 (
            .O(N__64231),
            .I(N__64183));
    CascadeMux I__14294 (
            .O(N__64230),
            .I(N__64179));
    InMux I__14293 (
            .O(N__64227),
            .I(N__64175));
    InMux I__14292 (
            .O(N__64224),
            .I(N__64172));
    InMux I__14291 (
            .O(N__64221),
            .I(N__64169));
    CascadeMux I__14290 (
            .O(N__64220),
            .I(N__64166));
    InMux I__14289 (
            .O(N__64219),
            .I(N__64149));
    InMux I__14288 (
            .O(N__64216),
            .I(N__64149));
    InMux I__14287 (
            .O(N__64215),
            .I(N__64149));
    InMux I__14286 (
            .O(N__64212),
            .I(N__64149));
    InMux I__14285 (
            .O(N__64211),
            .I(N__64149));
    InMux I__14284 (
            .O(N__64208),
            .I(N__64149));
    InMux I__14283 (
            .O(N__64207),
            .I(N__64149));
    InMux I__14282 (
            .O(N__64204),
            .I(N__64149));
    InMux I__14281 (
            .O(N__64201),
            .I(N__64146));
    InMux I__14280 (
            .O(N__64200),
            .I(N__64133));
    InMux I__14279 (
            .O(N__64197),
            .I(N__64133));
    InMux I__14278 (
            .O(N__64196),
            .I(N__64133));
    InMux I__14277 (
            .O(N__64193),
            .I(N__64133));
    InMux I__14276 (
            .O(N__64192),
            .I(N__64133));
    InMux I__14275 (
            .O(N__64189),
            .I(N__64133));
    InMux I__14274 (
            .O(N__64186),
            .I(N__64129));
    InMux I__14273 (
            .O(N__64183),
            .I(N__64126));
    InMux I__14272 (
            .O(N__64182),
            .I(N__64123));
    InMux I__14271 (
            .O(N__64179),
            .I(N__64120));
    CascadeMux I__14270 (
            .O(N__64178),
            .I(N__64117));
    LocalMux I__14269 (
            .O(N__64175),
            .I(N__64112));
    LocalMux I__14268 (
            .O(N__64172),
            .I(N__64112));
    LocalMux I__14267 (
            .O(N__64169),
            .I(N__64108));
    InMux I__14266 (
            .O(N__64166),
            .I(N__64105));
    LocalMux I__14265 (
            .O(N__64149),
            .I(N__64102));
    LocalMux I__14264 (
            .O(N__64146),
            .I(N__64098));
    LocalMux I__14263 (
            .O(N__64133),
            .I(N__64095));
    InMux I__14262 (
            .O(N__64132),
            .I(N__64092));
    LocalMux I__14261 (
            .O(N__64129),
            .I(N__64081));
    LocalMux I__14260 (
            .O(N__64126),
            .I(N__64081));
    LocalMux I__14259 (
            .O(N__64123),
            .I(N__64081));
    LocalMux I__14258 (
            .O(N__64120),
            .I(N__64081));
    InMux I__14257 (
            .O(N__64117),
            .I(N__64078));
    Span4Mux_v I__14256 (
            .O(N__64112),
            .I(N__64075));
    InMux I__14255 (
            .O(N__64111),
            .I(N__64072));
    Span4Mux_h I__14254 (
            .O(N__64108),
            .I(N__64067));
    LocalMux I__14253 (
            .O(N__64105),
            .I(N__64067));
    Span4Mux_v I__14252 (
            .O(N__64102),
            .I(N__64064));
    InMux I__14251 (
            .O(N__64101),
            .I(N__64061));
    Span4Mux_v I__14250 (
            .O(N__64098),
            .I(N__64054));
    Span4Mux_h I__14249 (
            .O(N__64095),
            .I(N__64054));
    LocalMux I__14248 (
            .O(N__64092),
            .I(N__64054));
    InMux I__14247 (
            .O(N__64091),
            .I(N__64051));
    CascadeMux I__14246 (
            .O(N__64090),
            .I(N__64048));
    Span4Mux_v I__14245 (
            .O(N__64081),
            .I(N__64043));
    LocalMux I__14244 (
            .O(N__64078),
            .I(N__64043));
    Span4Mux_h I__14243 (
            .O(N__64075),
            .I(N__64038));
    LocalMux I__14242 (
            .O(N__64072),
            .I(N__64038));
    Span4Mux_v I__14241 (
            .O(N__64067),
            .I(N__64031));
    Span4Mux_h I__14240 (
            .O(N__64064),
            .I(N__64031));
    LocalMux I__14239 (
            .O(N__64061),
            .I(N__64031));
    Span4Mux_h I__14238 (
            .O(N__64054),
            .I(N__64026));
    LocalMux I__14237 (
            .O(N__64051),
            .I(N__64026));
    InMux I__14236 (
            .O(N__64048),
            .I(N__64023));
    Span4Mux_v I__14235 (
            .O(N__64043),
            .I(N__64020));
    Span4Mux_v I__14234 (
            .O(N__64038),
            .I(N__64017));
    Span4Mux_h I__14233 (
            .O(N__64031),
            .I(N__64014));
    Sp12to4 I__14232 (
            .O(N__64026),
            .I(N__64009));
    LocalMux I__14231 (
            .O(N__64023),
            .I(N__64009));
    Odrv4 I__14230 (
            .O(N__64020),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ));
    Odrv4 I__14229 (
            .O(N__64017),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ));
    Odrv4 I__14228 (
            .O(N__64014),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ));
    Odrv12 I__14227 (
            .O(N__64009),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ));
    InMux I__14226 (
            .O(N__64000),
            .I(N__63997));
    LocalMux I__14225 (
            .O(N__63997),
            .I(N__63994));
    Odrv4 I__14224 (
            .O(N__63994),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n170 ));
    InMux I__14223 (
            .O(N__63991),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18265 ));
    InMux I__14222 (
            .O(N__63988),
            .I(N__63985));
    LocalMux I__14221 (
            .O(N__63985),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n173 ));
    CascadeMux I__14220 (
            .O(N__63982),
            .I(N__63976));
    CascadeMux I__14219 (
            .O(N__63981),
            .I(N__63971));
    CascadeMux I__14218 (
            .O(N__63980),
            .I(N__63968));
    CascadeMux I__14217 (
            .O(N__63979),
            .I(N__63964));
    InMux I__14216 (
            .O(N__63976),
            .I(N__63959));
    InMux I__14215 (
            .O(N__63975),
            .I(N__63956));
    CascadeMux I__14214 (
            .O(N__63974),
            .I(N__63952));
    InMux I__14213 (
            .O(N__63971),
            .I(N__63943));
    InMux I__14212 (
            .O(N__63968),
            .I(N__63940));
    CascadeMux I__14211 (
            .O(N__63967),
            .I(N__63937));
    InMux I__14210 (
            .O(N__63964),
            .I(N__63933));
    CascadeMux I__14209 (
            .O(N__63963),
            .I(N__63930));
    CascadeMux I__14208 (
            .O(N__63962),
            .I(N__63926));
    LocalMux I__14207 (
            .O(N__63959),
            .I(N__63921));
    LocalMux I__14206 (
            .O(N__63956),
            .I(N__63921));
    CascadeMux I__14205 (
            .O(N__63955),
            .I(N__63918));
    InMux I__14204 (
            .O(N__63952),
            .I(N__63915));
    CascadeMux I__14203 (
            .O(N__63951),
            .I(N__63912));
    CascadeMux I__14202 (
            .O(N__63950),
            .I(N__63909));
    CascadeMux I__14201 (
            .O(N__63949),
            .I(N__63906));
    CascadeMux I__14200 (
            .O(N__63948),
            .I(N__63903));
    CascadeMux I__14199 (
            .O(N__63947),
            .I(N__63900));
    CascadeMux I__14198 (
            .O(N__63946),
            .I(N__63897));
    LocalMux I__14197 (
            .O(N__63943),
            .I(N__63885));
    LocalMux I__14196 (
            .O(N__63940),
            .I(N__63882));
    InMux I__14195 (
            .O(N__63937),
            .I(N__63879));
    CascadeMux I__14194 (
            .O(N__63936),
            .I(N__63876));
    LocalMux I__14193 (
            .O(N__63933),
            .I(N__63872));
    InMux I__14192 (
            .O(N__63930),
            .I(N__63869));
    CascadeMux I__14191 (
            .O(N__63929),
            .I(N__63866));
    InMux I__14190 (
            .O(N__63926),
            .I(N__63863));
    Span4Mux_h I__14189 (
            .O(N__63921),
            .I(N__63859));
    InMux I__14188 (
            .O(N__63918),
            .I(N__63856));
    LocalMux I__14187 (
            .O(N__63915),
            .I(N__63853));
    InMux I__14186 (
            .O(N__63912),
            .I(N__63846));
    InMux I__14185 (
            .O(N__63909),
            .I(N__63846));
    InMux I__14184 (
            .O(N__63906),
            .I(N__63846));
    InMux I__14183 (
            .O(N__63903),
            .I(N__63839));
    InMux I__14182 (
            .O(N__63900),
            .I(N__63839));
    InMux I__14181 (
            .O(N__63897),
            .I(N__63839));
    CascadeMux I__14180 (
            .O(N__63896),
            .I(N__63836));
    CascadeMux I__14179 (
            .O(N__63895),
            .I(N__63833));
    CascadeMux I__14178 (
            .O(N__63894),
            .I(N__63830));
    CascadeMux I__14177 (
            .O(N__63893),
            .I(N__63827));
    CascadeMux I__14176 (
            .O(N__63892),
            .I(N__63824));
    CascadeMux I__14175 (
            .O(N__63891),
            .I(N__63821));
    CascadeMux I__14174 (
            .O(N__63890),
            .I(N__63818));
    CascadeMux I__14173 (
            .O(N__63889),
            .I(N__63815));
    CascadeMux I__14172 (
            .O(N__63888),
            .I(N__63812));
    Span4Mux_v I__14171 (
            .O(N__63885),
            .I(N__63805));
    Span4Mux_h I__14170 (
            .O(N__63882),
            .I(N__63805));
    LocalMux I__14169 (
            .O(N__63879),
            .I(N__63805));
    InMux I__14168 (
            .O(N__63876),
            .I(N__63802));
    InMux I__14167 (
            .O(N__63875),
            .I(N__63799));
    Span4Mux_v I__14166 (
            .O(N__63872),
            .I(N__63794));
    LocalMux I__14165 (
            .O(N__63869),
            .I(N__63794));
    InMux I__14164 (
            .O(N__63866),
            .I(N__63791));
    LocalMux I__14163 (
            .O(N__63863),
            .I(N__63788));
    InMux I__14162 (
            .O(N__63862),
            .I(N__63785));
    Span4Mux_v I__14161 (
            .O(N__63859),
            .I(N__63780));
    LocalMux I__14160 (
            .O(N__63856),
            .I(N__63780));
    Span4Mux_v I__14159 (
            .O(N__63853),
            .I(N__63777));
    LocalMux I__14158 (
            .O(N__63846),
            .I(N__63772));
    LocalMux I__14157 (
            .O(N__63839),
            .I(N__63772));
    InMux I__14156 (
            .O(N__63836),
            .I(N__63763));
    InMux I__14155 (
            .O(N__63833),
            .I(N__63763));
    InMux I__14154 (
            .O(N__63830),
            .I(N__63763));
    InMux I__14153 (
            .O(N__63827),
            .I(N__63763));
    InMux I__14152 (
            .O(N__63824),
            .I(N__63754));
    InMux I__14151 (
            .O(N__63821),
            .I(N__63754));
    InMux I__14150 (
            .O(N__63818),
            .I(N__63754));
    InMux I__14149 (
            .O(N__63815),
            .I(N__63754));
    InMux I__14148 (
            .O(N__63812),
            .I(N__63751));
    Span4Mux_v I__14147 (
            .O(N__63805),
            .I(N__63746));
    LocalMux I__14146 (
            .O(N__63802),
            .I(N__63746));
    LocalMux I__14145 (
            .O(N__63799),
            .I(N__63739));
    Span4Mux_h I__14144 (
            .O(N__63794),
            .I(N__63739));
    LocalMux I__14143 (
            .O(N__63791),
            .I(N__63739));
    Span4Mux_h I__14142 (
            .O(N__63788),
            .I(N__63734));
    LocalMux I__14141 (
            .O(N__63785),
            .I(N__63734));
    Span4Mux_h I__14140 (
            .O(N__63780),
            .I(N__63731));
    Sp12to4 I__14139 (
            .O(N__63777),
            .I(N__63720));
    Span12Mux_s9_v I__14138 (
            .O(N__63772),
            .I(N__63720));
    LocalMux I__14137 (
            .O(N__63763),
            .I(N__63720));
    LocalMux I__14136 (
            .O(N__63754),
            .I(N__63720));
    LocalMux I__14135 (
            .O(N__63751),
            .I(N__63720));
    Span4Mux_h I__14134 (
            .O(N__63746),
            .I(N__63715));
    Span4Mux_h I__14133 (
            .O(N__63739),
            .I(N__63715));
    Odrv4 I__14132 (
            .O(N__63734),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ));
    Odrv4 I__14131 (
            .O(N__63731),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ));
    Odrv12 I__14130 (
            .O(N__63720),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ));
    Odrv4 I__14129 (
            .O(N__63715),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ));
    InMux I__14128 (
            .O(N__63706),
            .I(N__63703));
    LocalMux I__14127 (
            .O(N__63703),
            .I(N__63700));
    Odrv12 I__14126 (
            .O(N__63700),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n219 ));
    InMux I__14125 (
            .O(N__63697),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18266 ));
    InMux I__14124 (
            .O(N__63694),
            .I(N__63691));
    LocalMux I__14123 (
            .O(N__63691),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n222 ));
    CascadeMux I__14122 (
            .O(N__63688),
            .I(N__63683));
    CascadeMux I__14121 (
            .O(N__63687),
            .I(N__63679));
    CascadeMux I__14120 (
            .O(N__63686),
            .I(N__63676));
    InMux I__14119 (
            .O(N__63683),
            .I(N__63673));
    CascadeMux I__14118 (
            .O(N__63682),
            .I(N__63670));
    InMux I__14117 (
            .O(N__63679),
            .I(N__63665));
    InMux I__14116 (
            .O(N__63676),
            .I(N__63662));
    LocalMux I__14115 (
            .O(N__63673),
            .I(N__63659));
    InMux I__14114 (
            .O(N__63670),
            .I(N__63656));
    CascadeMux I__14113 (
            .O(N__63669),
            .I(N__63652));
    CascadeMux I__14112 (
            .O(N__63668),
            .I(N__63649));
    LocalMux I__14111 (
            .O(N__63665),
            .I(N__63644));
    LocalMux I__14110 (
            .O(N__63662),
            .I(N__63641));
    Span4Mux_v I__14109 (
            .O(N__63659),
            .I(N__63636));
    LocalMux I__14108 (
            .O(N__63656),
            .I(N__63636));
    CascadeMux I__14107 (
            .O(N__63655),
            .I(N__63627));
    InMux I__14106 (
            .O(N__63652),
            .I(N__63619));
    InMux I__14105 (
            .O(N__63649),
            .I(N__63616));
    CascadeMux I__14104 (
            .O(N__63648),
            .I(N__63613));
    CascadeMux I__14103 (
            .O(N__63647),
            .I(N__63610));
    Span4Mux_v I__14102 (
            .O(N__63644),
            .I(N__63600));
    Span4Mux_v I__14101 (
            .O(N__63641),
            .I(N__63600));
    Span4Mux_v I__14100 (
            .O(N__63636),
            .I(N__63600));
    CascadeMux I__14099 (
            .O(N__63635),
            .I(N__63596));
    CascadeMux I__14098 (
            .O(N__63634),
            .I(N__63592));
    CascadeMux I__14097 (
            .O(N__63633),
            .I(N__63588));
    CascadeMux I__14096 (
            .O(N__63632),
            .I(N__63584));
    CascadeMux I__14095 (
            .O(N__63631),
            .I(N__63581));
    InMux I__14094 (
            .O(N__63630),
            .I(N__63578));
    InMux I__14093 (
            .O(N__63627),
            .I(N__63575));
    CascadeMux I__14092 (
            .O(N__63626),
            .I(N__63572));
    CascadeMux I__14091 (
            .O(N__63625),
            .I(N__63569));
    CascadeMux I__14090 (
            .O(N__63624),
            .I(N__63566));
    CascadeMux I__14089 (
            .O(N__63623),
            .I(N__63562));
    CascadeMux I__14088 (
            .O(N__63622),
            .I(N__63558));
    LocalMux I__14087 (
            .O(N__63619),
            .I(N__63553));
    LocalMux I__14086 (
            .O(N__63616),
            .I(N__63553));
    InMux I__14085 (
            .O(N__63613),
            .I(N__63550));
    InMux I__14084 (
            .O(N__63610),
            .I(N__63547));
    CascadeMux I__14083 (
            .O(N__63609),
            .I(N__63544));
    CascadeMux I__14082 (
            .O(N__63608),
            .I(N__63541));
    InMux I__14081 (
            .O(N__63607),
            .I(N__63538));
    Span4Mux_h I__14080 (
            .O(N__63600),
            .I(N__63535));
    InMux I__14079 (
            .O(N__63599),
            .I(N__63518));
    InMux I__14078 (
            .O(N__63596),
            .I(N__63518));
    InMux I__14077 (
            .O(N__63595),
            .I(N__63518));
    InMux I__14076 (
            .O(N__63592),
            .I(N__63518));
    InMux I__14075 (
            .O(N__63591),
            .I(N__63518));
    InMux I__14074 (
            .O(N__63588),
            .I(N__63518));
    InMux I__14073 (
            .O(N__63587),
            .I(N__63518));
    InMux I__14072 (
            .O(N__63584),
            .I(N__63518));
    InMux I__14071 (
            .O(N__63581),
            .I(N__63515));
    LocalMux I__14070 (
            .O(N__63578),
            .I(N__63510));
    LocalMux I__14069 (
            .O(N__63575),
            .I(N__63510));
    InMux I__14068 (
            .O(N__63572),
            .I(N__63507));
    InMux I__14067 (
            .O(N__63569),
            .I(N__63504));
    InMux I__14066 (
            .O(N__63566),
            .I(N__63493));
    InMux I__14065 (
            .O(N__63565),
            .I(N__63493));
    InMux I__14064 (
            .O(N__63562),
            .I(N__63493));
    InMux I__14063 (
            .O(N__63561),
            .I(N__63493));
    InMux I__14062 (
            .O(N__63558),
            .I(N__63493));
    Span4Mux_v I__14061 (
            .O(N__63553),
            .I(N__63488));
    LocalMux I__14060 (
            .O(N__63550),
            .I(N__63488));
    LocalMux I__14059 (
            .O(N__63547),
            .I(N__63485));
    InMux I__14058 (
            .O(N__63544),
            .I(N__63482));
    InMux I__14057 (
            .O(N__63541),
            .I(N__63479));
    LocalMux I__14056 (
            .O(N__63538),
            .I(N__63472));
    Sp12to4 I__14055 (
            .O(N__63535),
            .I(N__63472));
    LocalMux I__14054 (
            .O(N__63518),
            .I(N__63472));
    LocalMux I__14053 (
            .O(N__63515),
            .I(N__63469));
    Span4Mux_h I__14052 (
            .O(N__63510),
            .I(N__63464));
    LocalMux I__14051 (
            .O(N__63507),
            .I(N__63464));
    LocalMux I__14050 (
            .O(N__63504),
            .I(N__63457));
    LocalMux I__14049 (
            .O(N__63493),
            .I(N__63457));
    Span4Mux_h I__14048 (
            .O(N__63488),
            .I(N__63457));
    Span4Mux_h I__14047 (
            .O(N__63485),
            .I(N__63454));
    LocalMux I__14046 (
            .O(N__63482),
            .I(N__63451));
    LocalMux I__14045 (
            .O(N__63479),
            .I(N__63448));
    Span12Mux_h I__14044 (
            .O(N__63472),
            .I(N__63443));
    Span12Mux_h I__14043 (
            .O(N__63469),
            .I(N__63443));
    Span4Mux_v I__14042 (
            .O(N__63464),
            .I(N__63438));
    Span4Mux_h I__14041 (
            .O(N__63457),
            .I(N__63438));
    Span4Mux_v I__14040 (
            .O(N__63454),
            .I(N__63433));
    Span4Mux_h I__14039 (
            .O(N__63451),
            .I(N__63433));
    Odrv12 I__14038 (
            .O(N__63448),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ));
    Odrv12 I__14037 (
            .O(N__63443),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ));
    Odrv4 I__14036 (
            .O(N__63438),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ));
    Odrv4 I__14035 (
            .O(N__63433),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ));
    InMux I__14034 (
            .O(N__63424),
            .I(N__63421));
    LocalMux I__14033 (
            .O(N__63421),
            .I(N__63418));
    Odrv4 I__14032 (
            .O(N__63418),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n268 ));
    InMux I__14031 (
            .O(N__63415),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18267 ));
    InMux I__14030 (
            .O(N__63412),
            .I(N__63409));
    LocalMux I__14029 (
            .O(N__63409),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n271 ));
    CascadeMux I__14028 (
            .O(N__63406),
            .I(N__63402));
    CascadeMux I__14027 (
            .O(N__63405),
            .I(N__63396));
    InMux I__14026 (
            .O(N__63402),
            .I(N__63393));
    CascadeMux I__14025 (
            .O(N__63401),
            .I(N__63390));
    CascadeMux I__14024 (
            .O(N__63400),
            .I(N__63386));
    CascadeMux I__14023 (
            .O(N__63399),
            .I(N__63379));
    InMux I__14022 (
            .O(N__63396),
            .I(N__63374));
    LocalMux I__14021 (
            .O(N__63393),
            .I(N__63371));
    InMux I__14020 (
            .O(N__63390),
            .I(N__63368));
    CascadeMux I__14019 (
            .O(N__63389),
            .I(N__63365));
    InMux I__14018 (
            .O(N__63386),
            .I(N__63362));
    CascadeMux I__14017 (
            .O(N__63385),
            .I(N__63355));
    CascadeMux I__14016 (
            .O(N__63384),
            .I(N__63352));
    CascadeMux I__14015 (
            .O(N__63383),
            .I(N__63349));
    CascadeMux I__14014 (
            .O(N__63382),
            .I(N__63346));
    InMux I__14013 (
            .O(N__63379),
            .I(N__63343));
    CascadeMux I__14012 (
            .O(N__63378),
            .I(N__63340));
    CascadeMux I__14011 (
            .O(N__63377),
            .I(N__63337));
    LocalMux I__14010 (
            .O(N__63374),
            .I(N__63329));
    Span4Mux_v I__14009 (
            .O(N__63371),
            .I(N__63329));
    LocalMux I__14008 (
            .O(N__63368),
            .I(N__63329));
    InMux I__14007 (
            .O(N__63365),
            .I(N__63326));
    LocalMux I__14006 (
            .O(N__63362),
            .I(N__63323));
    CascadeMux I__14005 (
            .O(N__63361),
            .I(N__63320));
    CascadeMux I__14004 (
            .O(N__63360),
            .I(N__63316));
    CascadeMux I__14003 (
            .O(N__63359),
            .I(N__63312));
    CascadeMux I__14002 (
            .O(N__63358),
            .I(N__63308));
    InMux I__14001 (
            .O(N__63355),
            .I(N__63305));
    InMux I__14000 (
            .O(N__63352),
            .I(N__63302));
    InMux I__13999 (
            .O(N__63349),
            .I(N__63299));
    InMux I__13998 (
            .O(N__63346),
            .I(N__63296));
    LocalMux I__13997 (
            .O(N__63343),
            .I(N__63293));
    InMux I__13996 (
            .O(N__63340),
            .I(N__63290));
    InMux I__13995 (
            .O(N__63337),
            .I(N__63287));
    CascadeMux I__13994 (
            .O(N__63336),
            .I(N__63281));
    Span4Mux_h I__13993 (
            .O(N__63329),
            .I(N__63274));
    LocalMux I__13992 (
            .O(N__63326),
            .I(N__63274));
    Span4Mux_h I__13991 (
            .O(N__63323),
            .I(N__63271));
    InMux I__13990 (
            .O(N__63320),
            .I(N__63268));
    InMux I__13989 (
            .O(N__63319),
            .I(N__63255));
    InMux I__13988 (
            .O(N__63316),
            .I(N__63255));
    InMux I__13987 (
            .O(N__63315),
            .I(N__63255));
    InMux I__13986 (
            .O(N__63312),
            .I(N__63255));
    InMux I__13985 (
            .O(N__63311),
            .I(N__63255));
    InMux I__13984 (
            .O(N__63308),
            .I(N__63255));
    LocalMux I__13983 (
            .O(N__63305),
            .I(N__63252));
    LocalMux I__13982 (
            .O(N__63302),
            .I(N__63247));
    LocalMux I__13981 (
            .O(N__63299),
            .I(N__63247));
    LocalMux I__13980 (
            .O(N__63296),
            .I(N__63238));
    Span4Mux_h I__13979 (
            .O(N__63293),
            .I(N__63238));
    LocalMux I__13978 (
            .O(N__63290),
            .I(N__63238));
    LocalMux I__13977 (
            .O(N__63287),
            .I(N__63238));
    CascadeMux I__13976 (
            .O(N__63286),
            .I(N__63234));
    CascadeMux I__13975 (
            .O(N__63285),
            .I(N__63230));
    CascadeMux I__13974 (
            .O(N__63284),
            .I(N__63226));
    InMux I__13973 (
            .O(N__63281),
            .I(N__63221));
    InMux I__13972 (
            .O(N__63280),
            .I(N__63221));
    CascadeMux I__13971 (
            .O(N__63279),
            .I(N__63218));
    Span4Mux_h I__13970 (
            .O(N__63274),
            .I(N__63215));
    Span4Mux_v I__13969 (
            .O(N__63271),
            .I(N__63210));
    LocalMux I__13968 (
            .O(N__63268),
            .I(N__63210));
    LocalMux I__13967 (
            .O(N__63255),
            .I(N__63207));
    Span4Mux_v I__13966 (
            .O(N__63252),
            .I(N__63200));
    Span4Mux_h I__13965 (
            .O(N__63247),
            .I(N__63200));
    Span4Mux_v I__13964 (
            .O(N__63238),
            .I(N__63200));
    InMux I__13963 (
            .O(N__63237),
            .I(N__63187));
    InMux I__13962 (
            .O(N__63234),
            .I(N__63187));
    InMux I__13961 (
            .O(N__63233),
            .I(N__63187));
    InMux I__13960 (
            .O(N__63230),
            .I(N__63187));
    InMux I__13959 (
            .O(N__63229),
            .I(N__63187));
    InMux I__13958 (
            .O(N__63226),
            .I(N__63187));
    LocalMux I__13957 (
            .O(N__63221),
            .I(N__63184));
    InMux I__13956 (
            .O(N__63218),
            .I(N__63181));
    Span4Mux_v I__13955 (
            .O(N__63215),
            .I(N__63177));
    Span4Mux_v I__13954 (
            .O(N__63210),
            .I(N__63174));
    Span4Mux_v I__13953 (
            .O(N__63207),
            .I(N__63167));
    Span4Mux_h I__13952 (
            .O(N__63200),
            .I(N__63167));
    LocalMux I__13951 (
            .O(N__63187),
            .I(N__63167));
    Span4Mux_h I__13950 (
            .O(N__63184),
            .I(N__63162));
    LocalMux I__13949 (
            .O(N__63181),
            .I(N__63162));
    InMux I__13948 (
            .O(N__63180),
            .I(N__63159));
    Odrv4 I__13947 (
            .O(N__63177),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ));
    Odrv4 I__13946 (
            .O(N__63174),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ));
    Odrv4 I__13945 (
            .O(N__63167),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ));
    Odrv4 I__13944 (
            .O(N__63162),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ));
    LocalMux I__13943 (
            .O(N__63159),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ));
    InMux I__13942 (
            .O(N__63148),
            .I(N__63145));
    LocalMux I__13941 (
            .O(N__63145),
            .I(N__63142));
    Odrv4 I__13940 (
            .O(N__63142),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n317 ));
    InMux I__13939 (
            .O(N__63139),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18268 ));
    CascadeMux I__13938 (
            .O(N__63136),
            .I(N__63128));
    CascadeMux I__13937 (
            .O(N__63135),
            .I(N__63124));
    CascadeMux I__13936 (
            .O(N__63134),
            .I(N__63121));
    CascadeMux I__13935 (
            .O(N__63133),
            .I(N__63118));
    CascadeMux I__13934 (
            .O(N__63132),
            .I(N__63115));
    CascadeMux I__13933 (
            .O(N__63131),
            .I(N__63106));
    InMux I__13932 (
            .O(N__63128),
            .I(N__63103));
    CascadeMux I__13931 (
            .O(N__63127),
            .I(N__63100));
    InMux I__13930 (
            .O(N__63124),
            .I(N__63084));
    InMux I__13929 (
            .O(N__63121),
            .I(N__63084));
    InMux I__13928 (
            .O(N__63118),
            .I(N__63084));
    InMux I__13927 (
            .O(N__63115),
            .I(N__63084));
    CascadeMux I__13926 (
            .O(N__63114),
            .I(N__63081));
    CascadeMux I__13925 (
            .O(N__63113),
            .I(N__63078));
    CascadeMux I__13924 (
            .O(N__63112),
            .I(N__63075));
    CascadeMux I__13923 (
            .O(N__63111),
            .I(N__63072));
    InMux I__13922 (
            .O(N__63110),
            .I(N__63069));
    CascadeMux I__13921 (
            .O(N__63109),
            .I(N__63066));
    InMux I__13920 (
            .O(N__63106),
            .I(N__63062));
    LocalMux I__13919 (
            .O(N__63103),
            .I(N__63059));
    InMux I__13918 (
            .O(N__63100),
            .I(N__63056));
    CascadeMux I__13917 (
            .O(N__63099),
            .I(N__63053));
    CascadeMux I__13916 (
            .O(N__63098),
            .I(N__63049));
    CascadeMux I__13915 (
            .O(N__63097),
            .I(N__63045));
    CascadeMux I__13914 (
            .O(N__63096),
            .I(N__63041));
    CascadeMux I__13913 (
            .O(N__63095),
            .I(N__63038));
    InMux I__13912 (
            .O(N__63094),
            .I(N__63035));
    InMux I__13911 (
            .O(N__63093),
            .I(N__63032));
    LocalMux I__13910 (
            .O(N__63084),
            .I(N__63028));
    InMux I__13909 (
            .O(N__63081),
            .I(N__63019));
    InMux I__13908 (
            .O(N__63078),
            .I(N__63019));
    InMux I__13907 (
            .O(N__63075),
            .I(N__63019));
    InMux I__13906 (
            .O(N__63072),
            .I(N__63019));
    LocalMux I__13905 (
            .O(N__63069),
            .I(N__63016));
    InMux I__13904 (
            .O(N__63066),
            .I(N__63013));
    CascadeMux I__13903 (
            .O(N__63065),
            .I(N__63010));
    LocalMux I__13902 (
            .O(N__63062),
            .I(N__63003));
    Span4Mux_v I__13901 (
            .O(N__63059),
            .I(N__63003));
    LocalMux I__13900 (
            .O(N__63056),
            .I(N__63003));
    InMux I__13899 (
            .O(N__63053),
            .I(N__63000));
    InMux I__13898 (
            .O(N__63052),
            .I(N__62986));
    InMux I__13897 (
            .O(N__63049),
            .I(N__62986));
    InMux I__13896 (
            .O(N__63048),
            .I(N__62986));
    InMux I__13895 (
            .O(N__63045),
            .I(N__62986));
    InMux I__13894 (
            .O(N__63044),
            .I(N__62986));
    InMux I__13893 (
            .O(N__63041),
            .I(N__62986));
    InMux I__13892 (
            .O(N__63038),
            .I(N__62983));
    LocalMux I__13891 (
            .O(N__63035),
            .I(N__62978));
    LocalMux I__13890 (
            .O(N__63032),
            .I(N__62978));
    CascadeMux I__13889 (
            .O(N__63031),
            .I(N__62975));
    Span4Mux_v I__13888 (
            .O(N__63028),
            .I(N__62971));
    LocalMux I__13887 (
            .O(N__63019),
            .I(N__62968));
    Span4Mux_h I__13886 (
            .O(N__63016),
            .I(N__62963));
    LocalMux I__13885 (
            .O(N__63013),
            .I(N__62963));
    InMux I__13884 (
            .O(N__63010),
            .I(N__62960));
    Span4Mux_h I__13883 (
            .O(N__63003),
            .I(N__62954));
    LocalMux I__13882 (
            .O(N__63000),
            .I(N__62954));
    InMux I__13881 (
            .O(N__62999),
            .I(N__62951));
    LocalMux I__13880 (
            .O(N__62986),
            .I(N__62948));
    LocalMux I__13879 (
            .O(N__62983),
            .I(N__62945));
    Span4Mux_v I__13878 (
            .O(N__62978),
            .I(N__62942));
    InMux I__13877 (
            .O(N__62975),
            .I(N__62939));
    CascadeMux I__13876 (
            .O(N__62974),
            .I(N__62935));
    Span4Mux_h I__13875 (
            .O(N__62971),
            .I(N__62930));
    Span4Mux_v I__13874 (
            .O(N__62968),
            .I(N__62930));
    Span4Mux_v I__13873 (
            .O(N__62963),
            .I(N__62925));
    LocalMux I__13872 (
            .O(N__62960),
            .I(N__62925));
    CascadeMux I__13871 (
            .O(N__62959),
            .I(N__62922));
    Span4Mux_v I__13870 (
            .O(N__62954),
            .I(N__62919));
    LocalMux I__13869 (
            .O(N__62951),
            .I(N__62916));
    Span4Mux_v I__13868 (
            .O(N__62948),
            .I(N__62913));
    Span4Mux_v I__13867 (
            .O(N__62945),
            .I(N__62906));
    Span4Mux_h I__13866 (
            .O(N__62942),
            .I(N__62906));
    LocalMux I__13865 (
            .O(N__62939),
            .I(N__62906));
    InMux I__13864 (
            .O(N__62938),
            .I(N__62903));
    InMux I__13863 (
            .O(N__62935),
            .I(N__62900));
    Span4Mux_h I__13862 (
            .O(N__62930),
            .I(N__62895));
    Span4Mux_v I__13861 (
            .O(N__62925),
            .I(N__62895));
    InMux I__13860 (
            .O(N__62922),
            .I(N__62892));
    Span4Mux_h I__13859 (
            .O(N__62919),
            .I(N__62887));
    Span4Mux_v I__13858 (
            .O(N__62916),
            .I(N__62887));
    Span4Mux_h I__13857 (
            .O(N__62913),
            .I(N__62882));
    Span4Mux_h I__13856 (
            .O(N__62906),
            .I(N__62882));
    LocalMux I__13855 (
            .O(N__62903),
            .I(N__62879));
    LocalMux I__13854 (
            .O(N__62900),
            .I(N__62872));
    Span4Mux_h I__13853 (
            .O(N__62895),
            .I(N__62872));
    LocalMux I__13852 (
            .O(N__62892),
            .I(N__62872));
    Span4Mux_v I__13851 (
            .O(N__62887),
            .I(N__62869));
    Span4Mux_v I__13850 (
            .O(N__62882),
            .I(N__62866));
    Span4Mux_h I__13849 (
            .O(N__62879),
            .I(N__62861));
    Span4Mux_v I__13848 (
            .O(N__62872),
            .I(N__62861));
    Odrv4 I__13847 (
            .O(N__62869),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n120 ));
    Odrv4 I__13846 (
            .O(N__62866),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n120 ));
    Odrv4 I__13845 (
            .O(N__62861),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n120 ));
    CascadeMux I__13844 (
            .O(N__62854),
            .I(N__62851));
    InMux I__13843 (
            .O(N__62851),
            .I(N__62848));
    LocalMux I__13842 (
            .O(N__62848),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n320 ));
    InMux I__13841 (
            .O(N__62845),
            .I(N__62842));
    LocalMux I__13840 (
            .O(N__62842),
            .I(N__62839));
    Odrv4 I__13839 (
            .O(N__62839),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n366 ));
    InMux I__13838 (
            .O(N__62836),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18269 ));
    InMux I__13837 (
            .O(N__62833),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18255 ));
    InMux I__13836 (
            .O(N__62830),
            .I(N__62827));
    LocalMux I__13835 (
            .O(N__62827),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n461 ));
    InMux I__13834 (
            .O(N__62824),
            .I(bfn_23_26_0_));
    InMux I__13833 (
            .O(N__62821),
            .I(N__62818));
    LocalMux I__13832 (
            .O(N__62818),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n510 ));
    InMux I__13831 (
            .O(N__62815),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18257 ));
    InMux I__13830 (
            .O(N__62812),
            .I(N__62809));
    LocalMux I__13829 (
            .O(N__62809),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n559 ));
    InMux I__13828 (
            .O(N__62806),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18258 ));
    InMux I__13827 (
            .O(N__62803),
            .I(N__62800));
    LocalMux I__13826 (
            .O(N__62800),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n608 ));
    InMux I__13825 (
            .O(N__62797),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18259 ));
    CascadeMux I__13824 (
            .O(N__62794),
            .I(N__62791));
    InMux I__13823 (
            .O(N__62791),
            .I(N__62788));
    LocalMux I__13822 (
            .O(N__62788),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n657 ));
    InMux I__13821 (
            .O(N__62785),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18260 ));
    CascadeMux I__13820 (
            .O(N__62782),
            .I(N__62779));
    InMux I__13819 (
            .O(N__62779),
            .I(N__62776));
    LocalMux I__13818 (
            .O(N__62776),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n706 ));
    InMux I__13817 (
            .O(N__62773),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18261 ));
    InMux I__13816 (
            .O(N__62770),
            .I(N__62767));
    LocalMux I__13815 (
            .O(N__62767),
            .I(N__62764));
    Span4Mux_v I__13814 (
            .O(N__62764),
            .I(N__62761));
    Span4Mux_h I__13813 (
            .O(N__62761),
            .I(N__62758));
    Odrv4 I__13812 (
            .O(N__62758),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n762 ));
    InMux I__13811 (
            .O(N__62755),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18262 ));
    InMux I__13810 (
            .O(N__62752),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763 ));
    CascadeMux I__13809 (
            .O(N__62749),
            .I(N__62746));
    InMux I__13808 (
            .O(N__62746),
            .I(N__62743));
    LocalMux I__13807 (
            .O(N__62743),
            .I(N__62740));
    Span4Mux_h I__13806 (
            .O(N__62740),
            .I(N__62737));
    Span4Mux_v I__13805 (
            .O(N__62737),
            .I(N__62734));
    Odrv4 I__13804 (
            .O(N__62734),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO ));
    InMux I__13803 (
            .O(N__62731),
            .I(N__62728));
    LocalMux I__13802 (
            .O(N__62728),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19755 ));
    InMux I__13801 (
            .O(N__62725),
            .I(N__62722));
    LocalMux I__13800 (
            .O(N__62722),
            .I(N__62718));
    InMux I__13799 (
            .O(N__62721),
            .I(N__62715));
    Span4Mux_h I__13798 (
            .O(N__62718),
            .I(N__62711));
    LocalMux I__13797 (
            .O(N__62715),
            .I(N__62708));
    InMux I__13796 (
            .O(N__62714),
            .I(N__62705));
    Odrv4 I__13795 (
            .O(N__62711),
            .I(Add_add_temp_11_adj_2409));
    Odrv4 I__13794 (
            .O(N__62708),
            .I(Add_add_temp_11_adj_2409));
    LocalMux I__13793 (
            .O(N__62705),
            .I(Add_add_temp_11_adj_2409));
    CascadeMux I__13792 (
            .O(N__62698),
            .I(N__62694));
    InMux I__13791 (
            .O(N__62697),
            .I(N__62691));
    InMux I__13790 (
            .O(N__62694),
            .I(N__62688));
    LocalMux I__13789 (
            .O(N__62691),
            .I(N__62684));
    LocalMux I__13788 (
            .O(N__62688),
            .I(N__62681));
    InMux I__13787 (
            .O(N__62687),
            .I(N__62678));
    Odrv12 I__13786 (
            .O(N__62684),
            .I(Add_add_temp_9_adj_2411));
    Odrv4 I__13785 (
            .O(N__62681),
            .I(Add_add_temp_9_adj_2411));
    LocalMux I__13784 (
            .O(N__62678),
            .I(Add_add_temp_9_adj_2411));
    InMux I__13783 (
            .O(N__62671),
            .I(N__62668));
    LocalMux I__13782 (
            .O(N__62668),
            .I(N__62664));
    InMux I__13781 (
            .O(N__62667),
            .I(N__62661));
    Span4Mux_v I__13780 (
            .O(N__62664),
            .I(N__62655));
    LocalMux I__13779 (
            .O(N__62661),
            .I(N__62655));
    InMux I__13778 (
            .O(N__62660),
            .I(N__62652));
    Odrv4 I__13777 (
            .O(N__62655),
            .I(Add_add_temp_10_adj_2410));
    LocalMux I__13776 (
            .O(N__62652),
            .I(Add_add_temp_10_adj_2410));
    InMux I__13775 (
            .O(N__62647),
            .I(N__62644));
    LocalMux I__13774 (
            .O(N__62644),
            .I(N__62641));
    Span4Mux_h I__13773 (
            .O(N__62641),
            .I(N__62638));
    Odrv4 I__13772 (
            .O(N__62638),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20718 ));
    InMux I__13771 (
            .O(N__62635),
            .I(N__62632));
    LocalMux I__13770 (
            .O(N__62632),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n72 ));
    InMux I__13769 (
            .O(N__62629),
            .I(N__62626));
    LocalMux I__13768 (
            .O(N__62626),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n118 ));
    InMux I__13767 (
            .O(N__62623),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18249 ));
    InMux I__13766 (
            .O(N__62620),
            .I(N__62617));
    LocalMux I__13765 (
            .O(N__62617),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n167 ));
    InMux I__13764 (
            .O(N__62614),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18250 ));
    InMux I__13763 (
            .O(N__62611),
            .I(N__62608));
    LocalMux I__13762 (
            .O(N__62608),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n216 ));
    InMux I__13761 (
            .O(N__62605),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18251 ));
    InMux I__13760 (
            .O(N__62602),
            .I(N__62599));
    LocalMux I__13759 (
            .O(N__62599),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n265 ));
    InMux I__13758 (
            .O(N__62596),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18252 ));
    InMux I__13757 (
            .O(N__62593),
            .I(N__62590));
    LocalMux I__13756 (
            .O(N__62590),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n314 ));
    InMux I__13755 (
            .O(N__62587),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18253 ));
    InMux I__13754 (
            .O(N__62584),
            .I(N__62581));
    LocalMux I__13753 (
            .O(N__62581),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n363 ));
    InMux I__13752 (
            .O(N__62578),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18254 ));
    InMux I__13751 (
            .O(N__62575),
            .I(N__62572));
    LocalMux I__13750 (
            .O(N__62572),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n412 ));
    InMux I__13749 (
            .O(N__62569),
            .I(N__62566));
    LocalMux I__13748 (
            .O(N__62566),
            .I(N__62561));
    InMux I__13747 (
            .O(N__62565),
            .I(N__62556));
    InMux I__13746 (
            .O(N__62564),
            .I(N__62556));
    Odrv12 I__13745 (
            .O(N__62561),
            .I(Add_add_temp_5));
    LocalMux I__13744 (
            .O(N__62556),
            .I(Add_add_temp_5));
    InMux I__13743 (
            .O(N__62551),
            .I(N__62548));
    LocalMux I__13742 (
            .O(N__62548),
            .I(N__62544));
    InMux I__13741 (
            .O(N__62547),
            .I(N__62541));
    Odrv4 I__13740 (
            .O(N__62544),
            .I(Add_add_temp_4));
    LocalMux I__13739 (
            .O(N__62541),
            .I(Add_add_temp_4));
    InMux I__13738 (
            .O(N__62536),
            .I(N__62531));
    InMux I__13737 (
            .O(N__62535),
            .I(N__62528));
    InMux I__13736 (
            .O(N__62534),
            .I(N__62525));
    LocalMux I__13735 (
            .O(N__62531),
            .I(Add_add_temp_8));
    LocalMux I__13734 (
            .O(N__62528),
            .I(Add_add_temp_8));
    LocalMux I__13733 (
            .O(N__62525),
            .I(Add_add_temp_8));
    InMux I__13732 (
            .O(N__62518),
            .I(N__62513));
    CascadeMux I__13731 (
            .O(N__62517),
            .I(N__62510));
    InMux I__13730 (
            .O(N__62516),
            .I(N__62507));
    LocalMux I__13729 (
            .O(N__62513),
            .I(N__62504));
    InMux I__13728 (
            .O(N__62510),
            .I(N__62501));
    LocalMux I__13727 (
            .O(N__62507),
            .I(Add_add_temp_7));
    Odrv4 I__13726 (
            .O(N__62504),
            .I(Add_add_temp_7));
    LocalMux I__13725 (
            .O(N__62501),
            .I(Add_add_temp_7));
    CascadeMux I__13724 (
            .O(N__62494),
            .I(N__62491));
    InMux I__13723 (
            .O(N__62491),
            .I(N__62487));
    InMux I__13722 (
            .O(N__62490),
            .I(N__62484));
    LocalMux I__13721 (
            .O(N__62487),
            .I(N__62480));
    LocalMux I__13720 (
            .O(N__62484),
            .I(N__62477));
    InMux I__13719 (
            .O(N__62483),
            .I(N__62474));
    Odrv4 I__13718 (
            .O(N__62480),
            .I(Add_add_temp_6));
    Odrv12 I__13717 (
            .O(N__62477),
            .I(Add_add_temp_6));
    LocalMux I__13716 (
            .O(N__62474),
            .I(Add_add_temp_6));
    InMux I__13715 (
            .O(N__62467),
            .I(N__62464));
    LocalMux I__13714 (
            .O(N__62464),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20712 ));
    InMux I__13713 (
            .O(N__62461),
            .I(N__62456));
    InMux I__13712 (
            .O(N__62460),
            .I(N__62453));
    InMux I__13711 (
            .O(N__62459),
            .I(N__62450));
    LocalMux I__13710 (
            .O(N__62456),
            .I(Add_add_temp_9));
    LocalMux I__13709 (
            .O(N__62453),
            .I(Add_add_temp_9));
    LocalMux I__13708 (
            .O(N__62450),
            .I(Add_add_temp_9));
    InMux I__13707 (
            .O(N__62443),
            .I(N__62440));
    LocalMux I__13706 (
            .O(N__62440),
            .I(N__62437));
    Span4Mux_v I__13705 (
            .O(N__62437),
            .I(N__62432));
    InMux I__13704 (
            .O(N__62436),
            .I(N__62429));
    InMux I__13703 (
            .O(N__62435),
            .I(N__62426));
    Odrv4 I__13702 (
            .O(N__62432),
            .I(Add_add_temp_11));
    LocalMux I__13701 (
            .O(N__62429),
            .I(Add_add_temp_11));
    LocalMux I__13700 (
            .O(N__62426),
            .I(Add_add_temp_11));
    CascadeMux I__13699 (
            .O(N__62419),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_ ));
    InMux I__13698 (
            .O(N__62416),
            .I(N__62412));
    InMux I__13697 (
            .O(N__62415),
            .I(N__62408));
    LocalMux I__13696 (
            .O(N__62412),
            .I(N__62405));
    InMux I__13695 (
            .O(N__62411),
            .I(N__62402));
    LocalMux I__13694 (
            .O(N__62408),
            .I(Add_add_temp_10));
    Odrv4 I__13693 (
            .O(N__62405),
            .I(Add_add_temp_10));
    LocalMux I__13692 (
            .O(N__62402),
            .I(Add_add_temp_10));
    InMux I__13691 (
            .O(N__62395),
            .I(N__62392));
    LocalMux I__13690 (
            .O(N__62392),
            .I(N__62389));
    Span4Mux_h I__13689 (
            .O(N__62389),
            .I(N__62384));
    InMux I__13688 (
            .O(N__62388),
            .I(N__62381));
    InMux I__13687 (
            .O(N__62387),
            .I(N__62378));
    Odrv4 I__13686 (
            .O(N__62384),
            .I(Add_add_temp_14));
    LocalMux I__13685 (
            .O(N__62381),
            .I(Add_add_temp_14));
    LocalMux I__13684 (
            .O(N__62378),
            .I(Add_add_temp_14));
    InMux I__13683 (
            .O(N__62371),
            .I(N__62368));
    LocalMux I__13682 (
            .O(N__62368),
            .I(N__62363));
    InMux I__13681 (
            .O(N__62367),
            .I(N__62360));
    InMux I__13680 (
            .O(N__62366),
            .I(N__62357));
    Odrv4 I__13679 (
            .O(N__62363),
            .I(Add_add_temp_13));
    LocalMux I__13678 (
            .O(N__62360),
            .I(Add_add_temp_13));
    LocalMux I__13677 (
            .O(N__62357),
            .I(Add_add_temp_13));
    CascadeMux I__13676 (
            .O(N__62350),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_ ));
    InMux I__13675 (
            .O(N__62347),
            .I(N__62344));
    LocalMux I__13674 (
            .O(N__62344),
            .I(N__62341));
    Span4Mux_v I__13673 (
            .O(N__62341),
            .I(N__62336));
    InMux I__13672 (
            .O(N__62340),
            .I(N__62333));
    InMux I__13671 (
            .O(N__62339),
            .I(N__62330));
    Odrv4 I__13670 (
            .O(N__62336),
            .I(Add_add_temp_12));
    LocalMux I__13669 (
            .O(N__62333),
            .I(Add_add_temp_12));
    LocalMux I__13668 (
            .O(N__62330),
            .I(Add_add_temp_12));
    InMux I__13667 (
            .O(N__62323),
            .I(N__62320));
    LocalMux I__13666 (
            .O(N__62320),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15205 ));
    InMux I__13665 (
            .O(N__62317),
            .I(N__62314));
    LocalMux I__13664 (
            .O(N__62314),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20670 ));
    InMux I__13663 (
            .O(N__62311),
            .I(N__62308));
    LocalMux I__13662 (
            .O(N__62308),
            .I(N__62304));
    InMux I__13661 (
            .O(N__62307),
            .I(N__62301));
    Span4Mux_h I__13660 (
            .O(N__62304),
            .I(N__62297));
    LocalMux I__13659 (
            .O(N__62301),
            .I(N__62294));
    InMux I__13658 (
            .O(N__62300),
            .I(N__62291));
    Odrv4 I__13657 (
            .O(N__62297),
            .I(Add_add_temp_20));
    Odrv12 I__13656 (
            .O(N__62294),
            .I(Add_add_temp_20));
    LocalMux I__13655 (
            .O(N__62291),
            .I(Add_add_temp_20));
    CascadeMux I__13654 (
            .O(N__62284),
            .I(N__62280));
    InMux I__13653 (
            .O(N__62283),
            .I(N__62276));
    InMux I__13652 (
            .O(N__62280),
            .I(N__62273));
    CascadeMux I__13651 (
            .O(N__62279),
            .I(N__62270));
    LocalMux I__13650 (
            .O(N__62276),
            .I(N__62267));
    LocalMux I__13649 (
            .O(N__62273),
            .I(N__62264));
    InMux I__13648 (
            .O(N__62270),
            .I(N__62261));
    Odrv4 I__13647 (
            .O(N__62267),
            .I(Add_add_temp_18));
    Odrv4 I__13646 (
            .O(N__62264),
            .I(Add_add_temp_18));
    LocalMux I__13645 (
            .O(N__62261),
            .I(Add_add_temp_18));
    InMux I__13644 (
            .O(N__62254),
            .I(N__62251));
    LocalMux I__13643 (
            .O(N__62251),
            .I(N__62247));
    InMux I__13642 (
            .O(N__62250),
            .I(N__62244));
    Span4Mux_h I__13641 (
            .O(N__62247),
            .I(N__62238));
    LocalMux I__13640 (
            .O(N__62244),
            .I(N__62238));
    InMux I__13639 (
            .O(N__62243),
            .I(N__62235));
    Odrv4 I__13638 (
            .O(N__62238),
            .I(Add_add_temp_19));
    LocalMux I__13637 (
            .O(N__62235),
            .I(Add_add_temp_19));
    InMux I__13636 (
            .O(N__62230),
            .I(N__62227));
    LocalMux I__13635 (
            .O(N__62227),
            .I(N__62223));
    InMux I__13634 (
            .O(N__62226),
            .I(N__62220));
    Span4Mux_v I__13633 (
            .O(N__62223),
            .I(N__62215));
    LocalMux I__13632 (
            .O(N__62220),
            .I(N__62215));
    Span4Mux_h I__13631 (
            .O(N__62215),
            .I(N__62211));
    InMux I__13630 (
            .O(N__62214),
            .I(N__62208));
    Odrv4 I__13629 (
            .O(N__62211),
            .I(Add_add_temp_21));
    LocalMux I__13628 (
            .O(N__62208),
            .I(Add_add_temp_21));
    InMux I__13627 (
            .O(N__62203),
            .I(N__62199));
    InMux I__13626 (
            .O(N__62202),
            .I(N__62196));
    LocalMux I__13625 (
            .O(N__62199),
            .I(N__62191));
    LocalMux I__13624 (
            .O(N__62196),
            .I(N__62191));
    Span4Mux_h I__13623 (
            .O(N__62191),
            .I(N__62187));
    InMux I__13622 (
            .O(N__62190),
            .I(N__62184));
    Odrv4 I__13621 (
            .O(N__62187),
            .I(Add_add_temp_23));
    LocalMux I__13620 (
            .O(N__62184),
            .I(Add_add_temp_23));
    CascadeMux I__13619 (
            .O(N__62179),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_ ));
    InMux I__13618 (
            .O(N__62176),
            .I(N__62172));
    InMux I__13617 (
            .O(N__62175),
            .I(N__62169));
    LocalMux I__13616 (
            .O(N__62172),
            .I(N__62166));
    LocalMux I__13615 (
            .O(N__62169),
            .I(N__62160));
    Sp12to4 I__13614 (
            .O(N__62166),
            .I(N__62160));
    InMux I__13613 (
            .O(N__62165),
            .I(N__62157));
    Odrv12 I__13612 (
            .O(N__62160),
            .I(Add_add_temp_22));
    LocalMux I__13611 (
            .O(N__62157),
            .I(Add_add_temp_22));
    InMux I__13610 (
            .O(N__62152),
            .I(N__62149));
    LocalMux I__13609 (
            .O(N__62149),
            .I(N__62146));
    Odrv4 I__13608 (
            .O(N__62146),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20656 ));
    InMux I__13607 (
            .O(N__62143),
            .I(N__62139));
    InMux I__13606 (
            .O(N__62142),
            .I(N__62136));
    LocalMux I__13605 (
            .O(N__62139),
            .I(N__62131));
    LocalMux I__13604 (
            .O(N__62136),
            .I(N__62131));
    Span4Mux_v I__13603 (
            .O(N__62131),
            .I(N__62127));
    InMux I__13602 (
            .O(N__62130),
            .I(N__62124));
    Odrv4 I__13601 (
            .O(N__62127),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31 ));
    LocalMux I__13600 (
            .O(N__62124),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31 ));
    ClkMux I__13599 (
            .O(N__62119),
            .I(N__62071));
    ClkMux I__13598 (
            .O(N__62118),
            .I(N__62071));
    ClkMux I__13597 (
            .O(N__62117),
            .I(N__62071));
    ClkMux I__13596 (
            .O(N__62116),
            .I(N__62071));
    ClkMux I__13595 (
            .O(N__62115),
            .I(N__62071));
    ClkMux I__13594 (
            .O(N__62114),
            .I(N__62071));
    ClkMux I__13593 (
            .O(N__62113),
            .I(N__62071));
    ClkMux I__13592 (
            .O(N__62112),
            .I(N__62071));
    ClkMux I__13591 (
            .O(N__62111),
            .I(N__62071));
    ClkMux I__13590 (
            .O(N__62110),
            .I(N__62071));
    ClkMux I__13589 (
            .O(N__62109),
            .I(N__62071));
    ClkMux I__13588 (
            .O(N__62108),
            .I(N__62071));
    ClkMux I__13587 (
            .O(N__62107),
            .I(N__62071));
    ClkMux I__13586 (
            .O(N__62106),
            .I(N__62071));
    ClkMux I__13585 (
            .O(N__62105),
            .I(N__62071));
    ClkMux I__13584 (
            .O(N__62104),
            .I(N__62071));
    GlobalMux I__13583 (
            .O(N__62071),
            .I(N__62068));
    gio2CtrlBuf I__13582 (
            .O(N__62068),
            .I(pin3_clk_16mhz_N));
    InMux I__13581 (
            .O(N__62065),
            .I(N__62061));
    CascadeMux I__13580 (
            .O(N__62064),
            .I(N__62057));
    LocalMux I__13579 (
            .O(N__62061),
            .I(N__62054));
    InMux I__13578 (
            .O(N__62060),
            .I(N__62051));
    InMux I__13577 (
            .O(N__62057),
            .I(N__62048));
    Span4Mux_v I__13576 (
            .O(N__62054),
            .I(N__62045));
    LocalMux I__13575 (
            .O(N__62051),
            .I(N__62040));
    LocalMux I__13574 (
            .O(N__62048),
            .I(N__62040));
    Odrv4 I__13573 (
            .O(N__62045),
            .I(Add_add_temp_25));
    Odrv12 I__13572 (
            .O(N__62040),
            .I(Add_add_temp_25));
    InMux I__13571 (
            .O(N__62035),
            .I(N__62032));
    LocalMux I__13570 (
            .O(N__62032),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5 ));
    InMux I__13569 (
            .O(N__62029),
            .I(N__61998));
    InMux I__13568 (
            .O(N__62028),
            .I(N__61998));
    InMux I__13567 (
            .O(N__62027),
            .I(N__61998));
    InMux I__13566 (
            .O(N__62026),
            .I(N__61998));
    InMux I__13565 (
            .O(N__62025),
            .I(N__61998));
    InMux I__13564 (
            .O(N__62024),
            .I(N__61998));
    InMux I__13563 (
            .O(N__62023),
            .I(N__61998));
    InMux I__13562 (
            .O(N__62022),
            .I(N__61998));
    InMux I__13561 (
            .O(N__62021),
            .I(N__61987));
    InMux I__13560 (
            .O(N__62020),
            .I(N__61987));
    InMux I__13559 (
            .O(N__62019),
            .I(N__61987));
    InMux I__13558 (
            .O(N__62018),
            .I(N__61987));
    InMux I__13557 (
            .O(N__62017),
            .I(N__61987));
    CascadeMux I__13556 (
            .O(N__62016),
            .I(N__61982));
    CascadeMux I__13555 (
            .O(N__62015),
            .I(N__61978));
    LocalMux I__13554 (
            .O(N__61998),
            .I(N__61961));
    LocalMux I__13553 (
            .O(N__61987),
            .I(N__61961));
    InMux I__13552 (
            .O(N__61986),
            .I(N__61956));
    InMux I__13551 (
            .O(N__61985),
            .I(N__61956));
    InMux I__13550 (
            .O(N__61982),
            .I(N__61943));
    InMux I__13549 (
            .O(N__61981),
            .I(N__61943));
    InMux I__13548 (
            .O(N__61978),
            .I(N__61943));
    InMux I__13547 (
            .O(N__61977),
            .I(N__61943));
    InMux I__13546 (
            .O(N__61976),
            .I(N__61943));
    InMux I__13545 (
            .O(N__61975),
            .I(N__61943));
    InMux I__13544 (
            .O(N__61974),
            .I(N__61934));
    InMux I__13543 (
            .O(N__61973),
            .I(N__61934));
    InMux I__13542 (
            .O(N__61972),
            .I(N__61934));
    InMux I__13541 (
            .O(N__61971),
            .I(N__61934));
    InMux I__13540 (
            .O(N__61970),
            .I(N__61923));
    InMux I__13539 (
            .O(N__61969),
            .I(N__61923));
    InMux I__13538 (
            .O(N__61968),
            .I(N__61923));
    InMux I__13537 (
            .O(N__61967),
            .I(N__61923));
    InMux I__13536 (
            .O(N__61966),
            .I(N__61923));
    Odrv4 I__13535 (
            .O(N__61961),
            .I(Saturate_out1_31__N_267));
    LocalMux I__13534 (
            .O(N__61956),
            .I(Saturate_out1_31__N_267));
    LocalMux I__13533 (
            .O(N__61943),
            .I(Saturate_out1_31__N_267));
    LocalMux I__13532 (
            .O(N__61934),
            .I(Saturate_out1_31__N_267));
    LocalMux I__13531 (
            .O(N__61923),
            .I(Saturate_out1_31__N_267));
    InMux I__13530 (
            .O(N__61912),
            .I(N__61878));
    InMux I__13529 (
            .O(N__61911),
            .I(N__61878));
    InMux I__13528 (
            .O(N__61910),
            .I(N__61869));
    InMux I__13527 (
            .O(N__61909),
            .I(N__61869));
    InMux I__13526 (
            .O(N__61908),
            .I(N__61869));
    InMux I__13525 (
            .O(N__61907),
            .I(N__61869));
    InMux I__13524 (
            .O(N__61906),
            .I(N__61856));
    InMux I__13523 (
            .O(N__61905),
            .I(N__61856));
    InMux I__13522 (
            .O(N__61904),
            .I(N__61856));
    InMux I__13521 (
            .O(N__61903),
            .I(N__61856));
    InMux I__13520 (
            .O(N__61902),
            .I(N__61856));
    InMux I__13519 (
            .O(N__61901),
            .I(N__61856));
    InMux I__13518 (
            .O(N__61900),
            .I(N__61839));
    InMux I__13517 (
            .O(N__61899),
            .I(N__61839));
    InMux I__13516 (
            .O(N__61898),
            .I(N__61839));
    InMux I__13515 (
            .O(N__61897),
            .I(N__61839));
    InMux I__13514 (
            .O(N__61896),
            .I(N__61839));
    InMux I__13513 (
            .O(N__61895),
            .I(N__61839));
    InMux I__13512 (
            .O(N__61894),
            .I(N__61839));
    InMux I__13511 (
            .O(N__61893),
            .I(N__61839));
    InMux I__13510 (
            .O(N__61892),
            .I(N__61834));
    InMux I__13509 (
            .O(N__61891),
            .I(N__61834));
    InMux I__13508 (
            .O(N__61890),
            .I(N__61827));
    InMux I__13507 (
            .O(N__61889),
            .I(N__61827));
    InMux I__13506 (
            .O(N__61888),
            .I(N__61827));
    InMux I__13505 (
            .O(N__61887),
            .I(N__61822));
    InMux I__13504 (
            .O(N__61886),
            .I(N__61822));
    InMux I__13503 (
            .O(N__61885),
            .I(N__61815));
    InMux I__13502 (
            .O(N__61884),
            .I(N__61815));
    InMux I__13501 (
            .O(N__61883),
            .I(N__61815));
    LocalMux I__13500 (
            .O(N__61878),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13499 (
            .O(N__61869),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13498 (
            .O(N__61856),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13497 (
            .O(N__61839),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13496 (
            .O(N__61834),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13495 (
            .O(N__61827),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13494 (
            .O(N__61822),
            .I(Saturate_out1_31__N_266));
    LocalMux I__13493 (
            .O(N__61815),
            .I(Saturate_out1_31__N_266));
    CascadeMux I__13492 (
            .O(N__61798),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_ ));
    CascadeMux I__13491 (
            .O(N__61795),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_ ));
    CascadeMux I__13490 (
            .O(N__61792),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_ ));
    InMux I__13489 (
            .O(N__61789),
            .I(N__61786));
    LocalMux I__13488 (
            .O(N__61786),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20688 ));
    InMux I__13487 (
            .O(N__61783),
            .I(N__61780));
    LocalMux I__13486 (
            .O(N__61780),
            .I(N__61777));
    Span4Mux_h I__13485 (
            .O(N__61777),
            .I(N__61772));
    InMux I__13484 (
            .O(N__61776),
            .I(N__61767));
    InMux I__13483 (
            .O(N__61775),
            .I(N__61767));
    Odrv4 I__13482 (
            .O(N__61772),
            .I(Add_add_temp_17));
    LocalMux I__13481 (
            .O(N__61767),
            .I(Add_add_temp_17));
    InMux I__13480 (
            .O(N__61762),
            .I(N__61759));
    LocalMux I__13479 (
            .O(N__61759),
            .I(N__61755));
    CascadeMux I__13478 (
            .O(N__61758),
            .I(N__61751));
    Span4Mux_v I__13477 (
            .O(N__61755),
            .I(N__61748));
    InMux I__13476 (
            .O(N__61754),
            .I(N__61743));
    InMux I__13475 (
            .O(N__61751),
            .I(N__61743));
    Odrv4 I__13474 (
            .O(N__61748),
            .I(Add_add_temp_16));
    LocalMux I__13473 (
            .O(N__61743),
            .I(Add_add_temp_16));
    InMux I__13472 (
            .O(N__61738),
            .I(N__61735));
    LocalMux I__13471 (
            .O(N__61735),
            .I(N__61732));
    Span4Mux_h I__13470 (
            .O(N__61732),
            .I(N__61727));
    InMux I__13469 (
            .O(N__61731),
            .I(N__61722));
    InMux I__13468 (
            .O(N__61730),
            .I(N__61722));
    Odrv4 I__13467 (
            .O(N__61727),
            .I(Add_add_temp_15));
    LocalMux I__13466 (
            .O(N__61722),
            .I(Add_add_temp_15));
    InMux I__13465 (
            .O(N__61717),
            .I(N__61713));
    CascadeMux I__13464 (
            .O(N__61716),
            .I(N__61709));
    LocalMux I__13463 (
            .O(N__61713),
            .I(N__61706));
    InMux I__13462 (
            .O(N__61712),
            .I(N__61703));
    InMux I__13461 (
            .O(N__61709),
            .I(N__61700));
    Span4Mux_v I__13460 (
            .O(N__61706),
            .I(N__61697));
    LocalMux I__13459 (
            .O(N__61703),
            .I(N__61692));
    LocalMux I__13458 (
            .O(N__61700),
            .I(N__61692));
    Odrv4 I__13457 (
            .O(N__61697),
            .I(Add_add_temp_31));
    Odrv12 I__13456 (
            .O(N__61692),
            .I(Add_add_temp_31));
    InMux I__13455 (
            .O(N__61687),
            .I(N__61680));
    InMux I__13454 (
            .O(N__61686),
            .I(N__61680));
    InMux I__13453 (
            .O(N__61685),
            .I(N__61677));
    LocalMux I__13452 (
            .O(N__61680),
            .I(N__61674));
    LocalMux I__13451 (
            .O(N__61677),
            .I(N__61671));
    Span4Mux_v I__13450 (
            .O(N__61674),
            .I(N__61668));
    Span4Mux_v I__13449 (
            .O(N__61671),
            .I(N__61665));
    Odrv4 I__13448 (
            .O(N__61668),
            .I(Add_add_temp_32));
    Odrv4 I__13447 (
            .O(N__61665),
            .I(Add_add_temp_32));
    CascadeMux I__13446 (
            .O(N__61660),
            .I(N__61657));
    InMux I__13445 (
            .O(N__61657),
            .I(N__61650));
    InMux I__13444 (
            .O(N__61656),
            .I(N__61650));
    InMux I__13443 (
            .O(N__61655),
            .I(N__61647));
    LocalMux I__13442 (
            .O(N__61650),
            .I(N__61642));
    LocalMux I__13441 (
            .O(N__61647),
            .I(N__61642));
    Span4Mux_v I__13440 (
            .O(N__61642),
            .I(N__61639));
    Odrv4 I__13439 (
            .O(N__61639),
            .I(Add_add_temp_30));
    InMux I__13438 (
            .O(N__61636),
            .I(N__61633));
    LocalMux I__13437 (
            .O(N__61633),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20644 ));
    InMux I__13436 (
            .O(N__61630),
            .I(N__61626));
    InMux I__13435 (
            .O(N__61629),
            .I(N__61623));
    LocalMux I__13434 (
            .O(N__61626),
            .I(N__61619));
    LocalMux I__13433 (
            .O(N__61623),
            .I(N__61616));
    InMux I__13432 (
            .O(N__61622),
            .I(N__61613));
    Span4Mux_v I__13431 (
            .O(N__61619),
            .I(N__61610));
    Span12Mux_s10_h I__13430 (
            .O(N__61616),
            .I(N__61605));
    LocalMux I__13429 (
            .O(N__61613),
            .I(N__61605));
    Odrv4 I__13428 (
            .O(N__61610),
            .I(Add_add_temp_34));
    Odrv12 I__13427 (
            .O(N__61605),
            .I(Add_add_temp_34));
    CascadeMux I__13426 (
            .O(N__61600),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_ ));
    InMux I__13425 (
            .O(N__61597),
            .I(N__61593));
    InMux I__13424 (
            .O(N__61596),
            .I(N__61589));
    LocalMux I__13423 (
            .O(N__61593),
            .I(N__61586));
    InMux I__13422 (
            .O(N__61592),
            .I(N__61583));
    LocalMux I__13421 (
            .O(N__61589),
            .I(N__61580));
    Span4Mux_v I__13420 (
            .O(N__61586),
            .I(N__61575));
    LocalMux I__13419 (
            .O(N__61583),
            .I(N__61575));
    Span4Mux_h I__13418 (
            .O(N__61580),
            .I(N__61570));
    Span4Mux_h I__13417 (
            .O(N__61575),
            .I(N__61570));
    Span4Mux_v I__13416 (
            .O(N__61570),
            .I(N__61567));
    Odrv4 I__13415 (
            .O(N__61567),
            .I(Add_add_temp_33));
    CascadeMux I__13414 (
            .O(N__61564),
            .I(Saturate_out1_31__N_266_cascade_));
    InMux I__13413 (
            .O(N__61561),
            .I(N__61558));
    LocalMux I__13412 (
            .O(N__61558),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4 ));
    InMux I__13411 (
            .O(N__61555),
            .I(N__61552));
    LocalMux I__13410 (
            .O(N__61552),
            .I(N__61547));
    InMux I__13409 (
            .O(N__61551),
            .I(N__61542));
    InMux I__13408 (
            .O(N__61550),
            .I(N__61542));
    Span4Mux_v I__13407 (
            .O(N__61547),
            .I(N__61539));
    LocalMux I__13406 (
            .O(N__61542),
            .I(N__61536));
    Odrv4 I__13405 (
            .O(N__61539),
            .I(Add_add_temp_26));
    Odrv12 I__13404 (
            .O(N__61536),
            .I(Add_add_temp_26));
    InMux I__13403 (
            .O(N__61531),
            .I(N__61526));
    InMux I__13402 (
            .O(N__61530),
            .I(N__61521));
    InMux I__13401 (
            .O(N__61529),
            .I(N__61521));
    LocalMux I__13400 (
            .O(N__61526),
            .I(N__61516));
    LocalMux I__13399 (
            .O(N__61521),
            .I(N__61516));
    Span4Mux_v I__13398 (
            .O(N__61516),
            .I(N__61513));
    Odrv4 I__13397 (
            .O(N__61513),
            .I(Add_add_temp_27));
    CascadeMux I__13396 (
            .O(N__61510),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_ ));
    CascadeMux I__13395 (
            .O(N__61507),
            .I(\foc.dVoltage_13_cascade_ ));
    CascadeMux I__13394 (
            .O(N__61504),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_ ));
    InMux I__13393 (
            .O(N__61501),
            .I(N__61498));
    LocalMux I__13392 (
            .O(N__61498),
            .I(N__61495));
    Odrv4 I__13391 (
            .O(N__61495),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20576 ));
    InMux I__13390 (
            .O(N__61492),
            .I(N__61489));
    LocalMux I__13389 (
            .O(N__61489),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n14 ));
    InMux I__13388 (
            .O(N__61486),
            .I(N__61483));
    LocalMux I__13387 (
            .O(N__61483),
            .I(\foc.dVoltage_6 ));
    CascadeMux I__13386 (
            .O(N__61480),
            .I(N__61472));
    CascadeMux I__13385 (
            .O(N__61479),
            .I(N__61466));
    CascadeMux I__13384 (
            .O(N__61478),
            .I(N__61463));
    InMux I__13383 (
            .O(N__61477),
            .I(N__61455));
    CascadeMux I__13382 (
            .O(N__61476),
            .I(N__61451));
    CascadeMux I__13381 (
            .O(N__61475),
            .I(N__61446));
    InMux I__13380 (
            .O(N__61472),
            .I(N__61437));
    InMux I__13379 (
            .O(N__61471),
            .I(N__61437));
    InMux I__13378 (
            .O(N__61470),
            .I(N__61437));
    InMux I__13377 (
            .O(N__61469),
            .I(N__61437));
    InMux I__13376 (
            .O(N__61466),
            .I(N__61426));
    InMux I__13375 (
            .O(N__61463),
            .I(N__61426));
    InMux I__13374 (
            .O(N__61462),
            .I(N__61426));
    InMux I__13373 (
            .O(N__61461),
            .I(N__61426));
    InMux I__13372 (
            .O(N__61460),
            .I(N__61426));
    InMux I__13371 (
            .O(N__61459),
            .I(N__61421));
    InMux I__13370 (
            .O(N__61458),
            .I(N__61421));
    LocalMux I__13369 (
            .O(N__61455),
            .I(N__61418));
    InMux I__13368 (
            .O(N__61454),
            .I(N__61415));
    InMux I__13367 (
            .O(N__61451),
            .I(N__61412));
    InMux I__13366 (
            .O(N__61450),
            .I(N__61405));
    InMux I__13365 (
            .O(N__61449),
            .I(N__61405));
    InMux I__13364 (
            .O(N__61446),
            .I(N__61405));
    LocalMux I__13363 (
            .O(N__61437),
            .I(\foc.Out_31__N_332_adj_2312 ));
    LocalMux I__13362 (
            .O(N__61426),
            .I(\foc.Out_31__N_332_adj_2312 ));
    LocalMux I__13361 (
            .O(N__61421),
            .I(\foc.Out_31__N_332_adj_2312 ));
    Odrv12 I__13360 (
            .O(N__61418),
            .I(\foc.Out_31__N_332_adj_2312 ));
    LocalMux I__13359 (
            .O(N__61415),
            .I(\foc.Out_31__N_332_adj_2312 ));
    LocalMux I__13358 (
            .O(N__61412),
            .I(\foc.Out_31__N_332_adj_2312 ));
    LocalMux I__13357 (
            .O(N__61405),
            .I(\foc.Out_31__N_332_adj_2312 ));
    CascadeMux I__13356 (
            .O(N__61390),
            .I(N__61383));
    InMux I__13355 (
            .O(N__61389),
            .I(N__61368));
    InMux I__13354 (
            .O(N__61388),
            .I(N__61365));
    InMux I__13353 (
            .O(N__61387),
            .I(N__61356));
    InMux I__13352 (
            .O(N__61386),
            .I(N__61356));
    InMux I__13351 (
            .O(N__61383),
            .I(N__61356));
    InMux I__13350 (
            .O(N__61382),
            .I(N__61356));
    InMux I__13349 (
            .O(N__61381),
            .I(N__61347));
    InMux I__13348 (
            .O(N__61380),
            .I(N__61347));
    InMux I__13347 (
            .O(N__61379),
            .I(N__61347));
    InMux I__13346 (
            .O(N__61378),
            .I(N__61347));
    InMux I__13345 (
            .O(N__61377),
            .I(N__61336));
    InMux I__13344 (
            .O(N__61376),
            .I(N__61336));
    InMux I__13343 (
            .O(N__61375),
            .I(N__61336));
    InMux I__13342 (
            .O(N__61374),
            .I(N__61336));
    InMux I__13341 (
            .O(N__61373),
            .I(N__61336));
    InMux I__13340 (
            .O(N__61372),
            .I(N__61331));
    InMux I__13339 (
            .O(N__61371),
            .I(N__61331));
    LocalMux I__13338 (
            .O(N__61368),
            .I(\foc.Out_31__N_333_adj_2310 ));
    LocalMux I__13337 (
            .O(N__61365),
            .I(\foc.Out_31__N_333_adj_2310 ));
    LocalMux I__13336 (
            .O(N__61356),
            .I(\foc.Out_31__N_333_adj_2310 ));
    LocalMux I__13335 (
            .O(N__61347),
            .I(\foc.Out_31__N_333_adj_2310 ));
    LocalMux I__13334 (
            .O(N__61336),
            .I(\foc.Out_31__N_333_adj_2310 ));
    LocalMux I__13333 (
            .O(N__61331),
            .I(\foc.Out_31__N_333_adj_2310 ));
    InMux I__13332 (
            .O(N__61318),
            .I(N__61315));
    LocalMux I__13331 (
            .O(N__61315),
            .I(\foc.dVoltage_7 ));
    InMux I__13330 (
            .O(N__61312),
            .I(N__61309));
    LocalMux I__13329 (
            .O(N__61309),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747 ));
    InMux I__13328 (
            .O(N__61306),
            .I(N__61303));
    LocalMux I__13327 (
            .O(N__61303),
            .I(N__61300));
    Span4Mux_v I__13326 (
            .O(N__61300),
            .I(N__61297));
    Odrv4 I__13325 (
            .O(N__61297),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19858 ));
    InMux I__13324 (
            .O(N__61294),
            .I(N__61291));
    LocalMux I__13323 (
            .O(N__61291),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904 ));
    InMux I__13322 (
            .O(N__61288),
            .I(N__61285));
    LocalMux I__13321 (
            .O(N__61285),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n446 ));
    InMux I__13320 (
            .O(N__61282),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17529 ));
    InMux I__13319 (
            .O(N__61279),
            .I(N__61276));
    LocalMux I__13318 (
            .O(N__61276),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n495 ));
    InMux I__13317 (
            .O(N__61273),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17530 ));
    InMux I__13316 (
            .O(N__61270),
            .I(N__61267));
    LocalMux I__13315 (
            .O(N__61267),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n544 ));
    InMux I__13314 (
            .O(N__61264),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17531 ));
    InMux I__13313 (
            .O(N__61261),
            .I(N__61258));
    LocalMux I__13312 (
            .O(N__61258),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n593 ));
    InMux I__13311 (
            .O(N__61255),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17532 ));
    InMux I__13310 (
            .O(N__61252),
            .I(N__61249));
    LocalMux I__13309 (
            .O(N__61249),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n642 ));
    InMux I__13308 (
            .O(N__61246),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17533 ));
    InMux I__13307 (
            .O(N__61243),
            .I(N__61240));
    LocalMux I__13306 (
            .O(N__61240),
            .I(N__61237));
    Span4Mux_v I__13305 (
            .O(N__61237),
            .I(N__61233));
    InMux I__13304 (
            .O(N__61236),
            .I(N__61230));
    Span4Mux_h I__13303 (
            .O(N__61233),
            .I(N__61227));
    LocalMux I__13302 (
            .O(N__61230),
            .I(N__61224));
    Span4Mux_v I__13301 (
            .O(N__61227),
            .I(N__61221));
    Span4Mux_v I__13300 (
            .O(N__61224),
            .I(N__61218));
    Odrv4 I__13299 (
            .O(N__61221),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n737 ));
    Odrv4 I__13298 (
            .O(N__61218),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n737 ));
    CascadeMux I__13297 (
            .O(N__61213),
            .I(N__61210));
    InMux I__13296 (
            .O(N__61210),
            .I(N__61207));
    LocalMux I__13295 (
            .O(N__61207),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440 ));
    CascadeMux I__13294 (
            .O(N__61204),
            .I(N__61201));
    InMux I__13293 (
            .O(N__61201),
            .I(N__61197));
    InMux I__13292 (
            .O(N__61200),
            .I(N__61194));
    LocalMux I__13291 (
            .O(N__61197),
            .I(N__61189));
    LocalMux I__13290 (
            .O(N__61194),
            .I(N__61189));
    Span4Mux_h I__13289 (
            .O(N__61189),
            .I(N__61186));
    Odrv4 I__13288 (
            .O(N__61186),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n738 ));
    InMux I__13287 (
            .O(N__61183),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17534 ));
    InMux I__13286 (
            .O(N__61180),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n739 ));
    CascadeMux I__13285 (
            .O(N__61177),
            .I(N__61174));
    InMux I__13284 (
            .O(N__61174),
            .I(N__61171));
    LocalMux I__13283 (
            .O(N__61171),
            .I(N__61168));
    Span4Mux_v I__13282 (
            .O(N__61168),
            .I(N__61165));
    Odrv4 I__13281 (
            .O(N__61165),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO ));
    InMux I__13280 (
            .O(N__61162),
            .I(N__61159));
    LocalMux I__13279 (
            .O(N__61159),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932 ));
    InMux I__13278 (
            .O(N__61156),
            .I(N__61153));
    LocalMux I__13277 (
            .O(N__61153),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20546 ));
    CascadeMux I__13276 (
            .O(N__61150),
            .I(N__61147));
    InMux I__13275 (
            .O(N__61147),
            .I(N__61144));
    LocalMux I__13274 (
            .O(N__61144),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n54 ));
    InMux I__13273 (
            .O(N__61141),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17521 ));
    InMux I__13272 (
            .O(N__61138),
            .I(N__61135));
    LocalMux I__13271 (
            .O(N__61135),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n103 ));
    InMux I__13270 (
            .O(N__61132),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17522 ));
    CascadeMux I__13269 (
            .O(N__61129),
            .I(N__61126));
    InMux I__13268 (
            .O(N__61126),
            .I(N__61123));
    LocalMux I__13267 (
            .O(N__61123),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n152 ));
    InMux I__13266 (
            .O(N__61120),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17523 ));
    InMux I__13265 (
            .O(N__61117),
            .I(N__61114));
    LocalMux I__13264 (
            .O(N__61114),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n201 ));
    InMux I__13263 (
            .O(N__61111),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17524 ));
    CascadeMux I__13262 (
            .O(N__61108),
            .I(N__61105));
    InMux I__13261 (
            .O(N__61105),
            .I(N__61102));
    LocalMux I__13260 (
            .O(N__61102),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n250 ));
    InMux I__13259 (
            .O(N__61099),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17525 ));
    InMux I__13258 (
            .O(N__61096),
            .I(N__61093));
    LocalMux I__13257 (
            .O(N__61093),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n299 ));
    InMux I__13256 (
            .O(N__61090),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17526 ));
    CascadeMux I__13255 (
            .O(N__61087),
            .I(N__61084));
    InMux I__13254 (
            .O(N__61084),
            .I(N__61081));
    LocalMux I__13253 (
            .O(N__61081),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n348 ));
    InMux I__13252 (
            .O(N__61078),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17527 ));
    CascadeMux I__13251 (
            .O(N__61075),
            .I(N__61072));
    InMux I__13250 (
            .O(N__61072),
            .I(N__61069));
    LocalMux I__13249 (
            .O(N__61069),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n397 ));
    InMux I__13248 (
            .O(N__61066),
            .I(bfn_23_12_0_));
    InMux I__13247 (
            .O(N__61063),
            .I(N__61060));
    LocalMux I__13246 (
            .O(N__61060),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594 ));
    InMux I__13245 (
            .O(N__61057),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18287 ));
    InMux I__13244 (
            .O(N__61054),
            .I(N__61051));
    LocalMux I__13243 (
            .O(N__61051),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593 ));
    InMux I__13242 (
            .O(N__61048),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18288 ));
    InMux I__13241 (
            .O(N__61045),
            .I(N__61042));
    LocalMux I__13240 (
            .O(N__61042),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592 ));
    InMux I__13239 (
            .O(N__61039),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18289 ));
    InMux I__13238 (
            .O(N__61036),
            .I(N__61033));
    LocalMux I__13237 (
            .O(N__61033),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591 ));
    InMux I__13236 (
            .O(N__61030),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18290 ));
    CascadeMux I__13235 (
            .O(N__61027),
            .I(N__61024));
    InMux I__13234 (
            .O(N__61024),
            .I(N__61021));
    LocalMux I__13233 (
            .O(N__61021),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n666 ));
    InMux I__13232 (
            .O(N__61018),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18291 ));
    CascadeMux I__13231 (
            .O(N__61015),
            .I(N__61012));
    InMux I__13230 (
            .O(N__61012),
            .I(N__61009));
    LocalMux I__13229 (
            .O(N__61009),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n715 ));
    InMux I__13228 (
            .O(N__61006),
            .I(N__61003));
    LocalMux I__13227 (
            .O(N__61003),
            .I(N__61000));
    Span4Mux_h I__13226 (
            .O(N__61000),
            .I(N__60997));
    Span4Mux_v I__13225 (
            .O(N__60997),
            .I(N__60994));
    Odrv4 I__13224 (
            .O(N__60994),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n770 ));
    InMux I__13223 (
            .O(N__60991),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18292 ));
    InMux I__13222 (
            .O(N__60988),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771 ));
    CascadeMux I__13221 (
            .O(N__60985),
            .I(N__60982));
    InMux I__13220 (
            .O(N__60982),
            .I(N__60979));
    LocalMux I__13219 (
            .O(N__60979),
            .I(N__60976));
    Span4Mux_h I__13218 (
            .O(N__60976),
            .I(N__60973));
    Span4Mux_v I__13217 (
            .O(N__60973),
            .I(N__60970));
    Odrv4 I__13216 (
            .O(N__60970),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO ));
    InMux I__13215 (
            .O(N__60967),
            .I(N__60963));
    InMux I__13214 (
            .O(N__60966),
            .I(N__60960));
    LocalMux I__13213 (
            .O(N__60963),
            .I(N__60946));
    LocalMux I__13212 (
            .O(N__60960),
            .I(N__60946));
    InMux I__13211 (
            .O(N__60959),
            .I(N__60943));
    InMux I__13210 (
            .O(N__60958),
            .I(N__60940));
    CascadeMux I__13209 (
            .O(N__60957),
            .I(N__60935));
    CascadeMux I__13208 (
            .O(N__60956),
            .I(N__60931));
    CascadeMux I__13207 (
            .O(N__60955),
            .I(N__60927));
    CascadeMux I__13206 (
            .O(N__60954),
            .I(N__60923));
    CascadeMux I__13205 (
            .O(N__60953),
            .I(N__60919));
    CascadeMux I__13204 (
            .O(N__60952),
            .I(N__60915));
    CascadeMux I__13203 (
            .O(N__60951),
            .I(N__60911));
    Span4Mux_v I__13202 (
            .O(N__60946),
            .I(N__60904));
    LocalMux I__13201 (
            .O(N__60943),
            .I(N__60904));
    LocalMux I__13200 (
            .O(N__60940),
            .I(N__60904));
    InMux I__13199 (
            .O(N__60939),
            .I(N__60899));
    InMux I__13198 (
            .O(N__60938),
            .I(N__60886));
    InMux I__13197 (
            .O(N__60935),
            .I(N__60886));
    InMux I__13196 (
            .O(N__60934),
            .I(N__60886));
    InMux I__13195 (
            .O(N__60931),
            .I(N__60886));
    InMux I__13194 (
            .O(N__60930),
            .I(N__60886));
    InMux I__13193 (
            .O(N__60927),
            .I(N__60886));
    InMux I__13192 (
            .O(N__60926),
            .I(N__60869));
    InMux I__13191 (
            .O(N__60923),
            .I(N__60869));
    InMux I__13190 (
            .O(N__60922),
            .I(N__60869));
    InMux I__13189 (
            .O(N__60919),
            .I(N__60869));
    InMux I__13188 (
            .O(N__60918),
            .I(N__60869));
    InMux I__13187 (
            .O(N__60915),
            .I(N__60869));
    InMux I__13186 (
            .O(N__60914),
            .I(N__60869));
    InMux I__13185 (
            .O(N__60911),
            .I(N__60869));
    Span4Mux_v I__13184 (
            .O(N__60904),
            .I(N__60866));
    InMux I__13183 (
            .O(N__60903),
            .I(N__60863));
    InMux I__13182 (
            .O(N__60902),
            .I(N__60859));
    LocalMux I__13181 (
            .O(N__60899),
            .I(N__60853));
    LocalMux I__13180 (
            .O(N__60886),
            .I(N__60848));
    LocalMux I__13179 (
            .O(N__60869),
            .I(N__60848));
    Span4Mux_h I__13178 (
            .O(N__60866),
            .I(N__60843));
    LocalMux I__13177 (
            .O(N__60863),
            .I(N__60843));
    CascadeMux I__13176 (
            .O(N__60862),
            .I(N__60840));
    LocalMux I__13175 (
            .O(N__60859),
            .I(N__60836));
    InMux I__13174 (
            .O(N__60858),
            .I(N__60833));
    InMux I__13173 (
            .O(N__60857),
            .I(N__60830));
    InMux I__13172 (
            .O(N__60856),
            .I(N__60825));
    Span4Mux_v I__13171 (
            .O(N__60853),
            .I(N__60822));
    Span4Mux_v I__13170 (
            .O(N__60848),
            .I(N__60817));
    Span4Mux_v I__13169 (
            .O(N__60843),
            .I(N__60817));
    InMux I__13168 (
            .O(N__60840),
            .I(N__60814));
    InMux I__13167 (
            .O(N__60839),
            .I(N__60811));
    Span4Mux_h I__13166 (
            .O(N__60836),
            .I(N__60806));
    LocalMux I__13165 (
            .O(N__60833),
            .I(N__60806));
    LocalMux I__13164 (
            .O(N__60830),
            .I(N__60803));
    InMux I__13163 (
            .O(N__60829),
            .I(N__60800));
    InMux I__13162 (
            .O(N__60828),
            .I(N__60797));
    LocalMux I__13161 (
            .O(N__60825),
            .I(N__60793));
    Sp12to4 I__13160 (
            .O(N__60822),
            .I(N__60786));
    Sp12to4 I__13159 (
            .O(N__60817),
            .I(N__60786));
    LocalMux I__13158 (
            .O(N__60814),
            .I(N__60786));
    LocalMux I__13157 (
            .O(N__60811),
            .I(N__60783));
    Span4Mux_v I__13156 (
            .O(N__60806),
            .I(N__60774));
    Span4Mux_h I__13155 (
            .O(N__60803),
            .I(N__60774));
    LocalMux I__13154 (
            .O(N__60800),
            .I(N__60774));
    LocalMux I__13153 (
            .O(N__60797),
            .I(N__60774));
    InMux I__13152 (
            .O(N__60796),
            .I(N__60771));
    Span4Mux_v I__13151 (
            .O(N__60793),
            .I(N__60768));
    Span12Mux_h I__13150 (
            .O(N__60786),
            .I(N__60765));
    Span4Mux_h I__13149 (
            .O(N__60783),
            .I(N__60762));
    Span4Mux_v I__13148 (
            .O(N__60774),
            .I(N__60757));
    LocalMux I__13147 (
            .O(N__60771),
            .I(N__60757));
    Odrv4 I__13146 (
            .O(N__60768),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n102 ));
    Odrv12 I__13145 (
            .O(N__60765),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n102 ));
    Odrv4 I__13144 (
            .O(N__60762),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n102 ));
    Odrv4 I__13143 (
            .O(N__60757),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n102 ));
    InMux I__13142 (
            .O(N__60748),
            .I(N__60745));
    LocalMux I__13141 (
            .O(N__60745),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n78 ));
    InMux I__13140 (
            .O(N__60742),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18279 ));
    InMux I__13139 (
            .O(N__60739),
            .I(N__60736));
    LocalMux I__13138 (
            .O(N__60736),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n127 ));
    InMux I__13137 (
            .O(N__60733),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18280 ));
    InMux I__13136 (
            .O(N__60730),
            .I(N__60727));
    LocalMux I__13135 (
            .O(N__60727),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n176 ));
    InMux I__13134 (
            .O(N__60724),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18281 ));
    InMux I__13133 (
            .O(N__60721),
            .I(N__60718));
    LocalMux I__13132 (
            .O(N__60718),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n225 ));
    InMux I__13131 (
            .O(N__60715),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18282 ));
    InMux I__13130 (
            .O(N__60712),
            .I(N__60709));
    LocalMux I__13129 (
            .O(N__60709),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n274 ));
    InMux I__13128 (
            .O(N__60706),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18283 ));
    InMux I__13127 (
            .O(N__60703),
            .I(N__60700));
    LocalMux I__13126 (
            .O(N__60700),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n323 ));
    InMux I__13125 (
            .O(N__60697),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18284 ));
    CascadeMux I__13124 (
            .O(N__60694),
            .I(N__60691));
    InMux I__13123 (
            .O(N__60691),
            .I(N__60688));
    LocalMux I__13122 (
            .O(N__60688),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596 ));
    InMux I__13121 (
            .O(N__60685),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18285 ));
    InMux I__13120 (
            .O(N__60682),
            .I(N__60679));
    LocalMux I__13119 (
            .O(N__60679),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595 ));
    InMux I__13118 (
            .O(N__60676),
            .I(bfn_22_29_0_));
    InMux I__13117 (
            .O(N__60673),
            .I(N__60670));
    LocalMux I__13116 (
            .O(N__60670),
            .I(N__60667));
    Odrv12 I__13115 (
            .O(N__60667),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n458 ));
    InMux I__13114 (
            .O(N__60664),
            .I(bfn_22_26_0_));
    InMux I__13113 (
            .O(N__60661),
            .I(N__60658));
    LocalMux I__13112 (
            .O(N__60658),
            .I(N__60655));
    Odrv12 I__13111 (
            .O(N__60655),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n507 ));
    InMux I__13110 (
            .O(N__60652),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18242 ));
    InMux I__13109 (
            .O(N__60649),
            .I(N__60646));
    LocalMux I__13108 (
            .O(N__60646),
            .I(N__60643));
    Odrv12 I__13107 (
            .O(N__60643),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n556 ));
    InMux I__13106 (
            .O(N__60640),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18243 ));
    InMux I__13105 (
            .O(N__60637),
            .I(N__60634));
    LocalMux I__13104 (
            .O(N__60634),
            .I(N__60631));
    Odrv12 I__13103 (
            .O(N__60631),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n605 ));
    InMux I__13102 (
            .O(N__60628),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18244 ));
    CascadeMux I__13101 (
            .O(N__60625),
            .I(N__60622));
    InMux I__13100 (
            .O(N__60622),
            .I(N__60619));
    LocalMux I__13099 (
            .O(N__60619),
            .I(N__60616));
    Odrv12 I__13098 (
            .O(N__60616),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n654 ));
    InMux I__13097 (
            .O(N__60613),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18245 ));
    CascadeMux I__13096 (
            .O(N__60610),
            .I(N__60607));
    InMux I__13095 (
            .O(N__60607),
            .I(N__60604));
    LocalMux I__13094 (
            .O(N__60604),
            .I(N__60601));
    Odrv4 I__13093 (
            .O(N__60601),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n703 ));
    InMux I__13092 (
            .O(N__60598),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18246 ));
    InMux I__13091 (
            .O(N__60595),
            .I(N__60592));
    LocalMux I__13090 (
            .O(N__60592),
            .I(N__60589));
    Span4Mux_v I__13089 (
            .O(N__60589),
            .I(N__60586));
    Span4Mux_v I__13088 (
            .O(N__60586),
            .I(N__60583));
    Odrv4 I__13087 (
            .O(N__60583),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n758 ));
    InMux I__13086 (
            .O(N__60580),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18247 ));
    InMux I__13085 (
            .O(N__60577),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759 ));
    CascadeMux I__13084 (
            .O(N__60574),
            .I(N__60571));
    InMux I__13083 (
            .O(N__60571),
            .I(N__60568));
    LocalMux I__13082 (
            .O(N__60568),
            .I(N__60565));
    Span12Mux_h I__13081 (
            .O(N__60565),
            .I(N__60562));
    Odrv12 I__13080 (
            .O(N__60562),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO ));
    CascadeMux I__13079 (
            .O(N__60559),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_ ));
    InMux I__13078 (
            .O(N__60556),
            .I(N__60553));
    LocalMux I__13077 (
            .O(N__60553),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20704 ));
    InMux I__13076 (
            .O(N__60550),
            .I(N__60547));
    LocalMux I__13075 (
            .O(N__60547),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n69 ));
    InMux I__13074 (
            .O(N__60544),
            .I(N__60541));
    LocalMux I__13073 (
            .O(N__60541),
            .I(N__60538));
    Odrv12 I__13072 (
            .O(N__60538),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n115 ));
    InMux I__13071 (
            .O(N__60535),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18234 ));
    InMux I__13070 (
            .O(N__60532),
            .I(N__60529));
    LocalMux I__13069 (
            .O(N__60529),
            .I(N__60526));
    Odrv12 I__13068 (
            .O(N__60526),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n164 ));
    InMux I__13067 (
            .O(N__60523),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18235 ));
    InMux I__13066 (
            .O(N__60520),
            .I(N__60517));
    LocalMux I__13065 (
            .O(N__60517),
            .I(N__60514));
    Odrv12 I__13064 (
            .O(N__60514),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n213 ));
    InMux I__13063 (
            .O(N__60511),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18236 ));
    InMux I__13062 (
            .O(N__60508),
            .I(N__60505));
    LocalMux I__13061 (
            .O(N__60505),
            .I(N__60502));
    Odrv12 I__13060 (
            .O(N__60502),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n262 ));
    InMux I__13059 (
            .O(N__60499),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18237 ));
    CascadeMux I__13058 (
            .O(N__60496),
            .I(N__60493));
    InMux I__13057 (
            .O(N__60493),
            .I(N__60490));
    LocalMux I__13056 (
            .O(N__60490),
            .I(N__60487));
    Odrv4 I__13055 (
            .O(N__60487),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n311 ));
    InMux I__13054 (
            .O(N__60484),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18238 ));
    CascadeMux I__13053 (
            .O(N__60481),
            .I(N__60478));
    InMux I__13052 (
            .O(N__60478),
            .I(N__60475));
    LocalMux I__13051 (
            .O(N__60475),
            .I(N__60472));
    Odrv12 I__13050 (
            .O(N__60472),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n360 ));
    InMux I__13049 (
            .O(N__60469),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18239 ));
    InMux I__13048 (
            .O(N__60466),
            .I(N__60463));
    LocalMux I__13047 (
            .O(N__60463),
            .I(N__60460));
    Span4Mux_v I__13046 (
            .O(N__60460),
            .I(N__60457));
    Odrv4 I__13045 (
            .O(N__60457),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n409 ));
    InMux I__13044 (
            .O(N__60454),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18240 ));
    InMux I__13043 (
            .O(N__60451),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n16002 ));
    CascadeMux I__13042 (
            .O(N__60448),
            .I(N__60444));
    CascadeMux I__13041 (
            .O(N__60447),
            .I(N__60438));
    InMux I__13040 (
            .O(N__60444),
            .I(N__60433));
    InMux I__13039 (
            .O(N__60443),
            .I(N__60433));
    InMux I__13038 (
            .O(N__60442),
            .I(N__60426));
    InMux I__13037 (
            .O(N__60441),
            .I(N__60426));
    InMux I__13036 (
            .O(N__60438),
            .I(N__60426));
    LocalMux I__13035 (
            .O(N__60433),
            .I(N__60421));
    LocalMux I__13034 (
            .O(N__60426),
            .I(N__60421));
    Span4Mux_v I__13033 (
            .O(N__60421),
            .I(N__60418));
    Odrv4 I__13032 (
            .O(N__60418),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31 ));
    InMux I__13031 (
            .O(N__60415),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n16003 ));
    InMux I__13030 (
            .O(N__60412),
            .I(N__60408));
    InMux I__13029 (
            .O(N__60411),
            .I(N__60405));
    LocalMux I__13028 (
            .O(N__60408),
            .I(N__60402));
    LocalMux I__13027 (
            .O(N__60405),
            .I(N__60399));
    Span4Mux_h I__13026 (
            .O(N__60402),
            .I(N__60395));
    Span12Mux_h I__13025 (
            .O(N__60399),
            .I(N__60392));
    InMux I__13024 (
            .O(N__60398),
            .I(N__60389));
    Odrv4 I__13023 (
            .O(N__60395),
            .I(Add_add_temp_14_adj_2406));
    Odrv12 I__13022 (
            .O(N__60392),
            .I(Add_add_temp_14_adj_2406));
    LocalMux I__13021 (
            .O(N__60389),
            .I(Add_add_temp_14_adj_2406));
    InMux I__13020 (
            .O(N__60382),
            .I(N__60376));
    InMux I__13019 (
            .O(N__60381),
            .I(N__60376));
    LocalMux I__13018 (
            .O(N__60376),
            .I(N__60372));
    CascadeMux I__13017 (
            .O(N__60375),
            .I(N__60369));
    Span4Mux_v I__13016 (
            .O(N__60372),
            .I(N__60366));
    InMux I__13015 (
            .O(N__60369),
            .I(N__60363));
    Odrv4 I__13014 (
            .O(N__60366),
            .I(Add_add_temp_12_adj_2408));
    LocalMux I__13013 (
            .O(N__60363),
            .I(Add_add_temp_12_adj_2408));
    InMux I__13012 (
            .O(N__60358),
            .I(N__60355));
    LocalMux I__13011 (
            .O(N__60355),
            .I(N__60351));
    CascadeMux I__13010 (
            .O(N__60354),
            .I(N__60348));
    Span4Mux_h I__13009 (
            .O(N__60351),
            .I(N__60345));
    InMux I__13008 (
            .O(N__60348),
            .I(N__60342));
    Span4Mux_h I__13007 (
            .O(N__60345),
            .I(N__60336));
    LocalMux I__13006 (
            .O(N__60342),
            .I(N__60336));
    InMux I__13005 (
            .O(N__60341),
            .I(N__60333));
    Odrv4 I__13004 (
            .O(N__60336),
            .I(Add_add_temp_13_adj_2407));
    LocalMux I__13003 (
            .O(N__60333),
            .I(Add_add_temp_13_adj_2407));
    InMux I__13002 (
            .O(N__60328),
            .I(N__60322));
    InMux I__13001 (
            .O(N__60327),
            .I(N__60322));
    LocalMux I__13000 (
            .O(N__60322),
            .I(N__60318));
    InMux I__12999 (
            .O(N__60321),
            .I(N__60315));
    Odrv4 I__12998 (
            .O(N__60318),
            .I(Add_add_temp_16_adj_2404));
    LocalMux I__12997 (
            .O(N__60315),
            .I(Add_add_temp_16_adj_2404));
    InMux I__12996 (
            .O(N__60310),
            .I(N__60304));
    InMux I__12995 (
            .O(N__60309),
            .I(N__60304));
    LocalMux I__12994 (
            .O(N__60304),
            .I(N__60300));
    InMux I__12993 (
            .O(N__60303),
            .I(N__60297));
    Odrv4 I__12992 (
            .O(N__60300),
            .I(Add_add_temp_17_adj_2403));
    LocalMux I__12991 (
            .O(N__60297),
            .I(Add_add_temp_17_adj_2403));
    CascadeMux I__12990 (
            .O(N__60292),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_ ));
    InMux I__12989 (
            .O(N__60289),
            .I(N__60286));
    LocalMux I__12988 (
            .O(N__60286),
            .I(N__60282));
    InMux I__12987 (
            .O(N__60285),
            .I(N__60279));
    Span4Mux_v I__12986 (
            .O(N__60282),
            .I(N__60274));
    LocalMux I__12985 (
            .O(N__60279),
            .I(N__60274));
    Span4Mux_v I__12984 (
            .O(N__60274),
            .I(N__60271));
    Sp12to4 I__12983 (
            .O(N__60271),
            .I(N__60267));
    InMux I__12982 (
            .O(N__60270),
            .I(N__60264));
    Odrv12 I__12981 (
            .O(N__60267),
            .I(Add_add_temp_15_adj_2405));
    LocalMux I__12980 (
            .O(N__60264),
            .I(Add_add_temp_15_adj_2405));
    InMux I__12979 (
            .O(N__60259),
            .I(N__60255));
    InMux I__12978 (
            .O(N__60258),
            .I(N__60252));
    LocalMux I__12977 (
            .O(N__60255),
            .I(N__60248));
    LocalMux I__12976 (
            .O(N__60252),
            .I(N__60245));
    InMux I__12975 (
            .O(N__60251),
            .I(N__60242));
    Span4Mux_h I__12974 (
            .O(N__60248),
            .I(N__60239));
    Span4Mux_h I__12973 (
            .O(N__60245),
            .I(N__60234));
    LocalMux I__12972 (
            .O(N__60242),
            .I(N__60234));
    Odrv4 I__12971 (
            .O(N__60239),
            .I(Add_add_temp_20_adj_2400));
    Odrv4 I__12970 (
            .O(N__60234),
            .I(Add_add_temp_20_adj_2400));
    InMux I__12969 (
            .O(N__60229),
            .I(N__60226));
    LocalMux I__12968 (
            .O(N__60226),
            .I(N__60223));
    Span4Mux_h I__12967 (
            .O(N__60223),
            .I(N__60219));
    InMux I__12966 (
            .O(N__60222),
            .I(N__60216));
    Span4Mux_v I__12965 (
            .O(N__60219),
            .I(N__60212));
    LocalMux I__12964 (
            .O(N__60216),
            .I(N__60209));
    InMux I__12963 (
            .O(N__60215),
            .I(N__60206));
    Odrv4 I__12962 (
            .O(N__60212),
            .I(Add_add_temp_19_adj_2401));
    Odrv4 I__12961 (
            .O(N__60209),
            .I(Add_add_temp_19_adj_2401));
    LocalMux I__12960 (
            .O(N__60206),
            .I(Add_add_temp_19_adj_2401));
    CascadeMux I__12959 (
            .O(N__60199),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_ ));
    InMux I__12958 (
            .O(N__60196),
            .I(N__60193));
    LocalMux I__12957 (
            .O(N__60193),
            .I(N__60190));
    Span4Mux_h I__12956 (
            .O(N__60190),
            .I(N__60186));
    InMux I__12955 (
            .O(N__60189),
            .I(N__60183));
    Span4Mux_v I__12954 (
            .O(N__60186),
            .I(N__60178));
    LocalMux I__12953 (
            .O(N__60183),
            .I(N__60178));
    Span4Mux_v I__12952 (
            .O(N__60178),
            .I(N__60175));
    Span4Mux_h I__12951 (
            .O(N__60175),
            .I(N__60171));
    InMux I__12950 (
            .O(N__60174),
            .I(N__60168));
    Odrv4 I__12949 (
            .O(N__60171),
            .I(Add_add_temp_18_adj_2402));
    LocalMux I__12948 (
            .O(N__60168),
            .I(Add_add_temp_18_adj_2402));
    InMux I__12947 (
            .O(N__60163),
            .I(N__60160));
    LocalMux I__12946 (
            .O(N__60160),
            .I(N__60157));
    Span4Mux_h I__12945 (
            .O(N__60157),
            .I(N__60154));
    Odrv4 I__12944 (
            .O(N__60154),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19733 ));
    InMux I__12943 (
            .O(N__60151),
            .I(N__60148));
    LocalMux I__12942 (
            .O(N__60148),
            .I(N__60144));
    CascadeMux I__12941 (
            .O(N__60147),
            .I(N__60141));
    Span4Mux_h I__12940 (
            .O(N__60144),
            .I(N__60137));
    InMux I__12939 (
            .O(N__60141),
            .I(N__60132));
    InMux I__12938 (
            .O(N__60140),
            .I(N__60132));
    Odrv4 I__12937 (
            .O(N__60137),
            .I(Add_add_temp_5_adj_2415));
    LocalMux I__12936 (
            .O(N__60132),
            .I(Add_add_temp_5_adj_2415));
    InMux I__12935 (
            .O(N__60127),
            .I(N__60124));
    LocalMux I__12934 (
            .O(N__60124),
            .I(N__60120));
    InMux I__12933 (
            .O(N__60123),
            .I(N__60117));
    Odrv4 I__12932 (
            .O(N__60120),
            .I(Add_add_temp_4_adj_2416));
    LocalMux I__12931 (
            .O(N__60117),
            .I(Add_add_temp_4_adj_2416));
    InMux I__12930 (
            .O(N__60112),
            .I(N__60107));
    InMux I__12929 (
            .O(N__60111),
            .I(N__60102));
    InMux I__12928 (
            .O(N__60110),
            .I(N__60102));
    LocalMux I__12927 (
            .O(N__60107),
            .I(Add_add_temp_8_adj_2412));
    LocalMux I__12926 (
            .O(N__60102),
            .I(Add_add_temp_8_adj_2412));
    InMux I__12925 (
            .O(N__60097),
            .I(N__60094));
    LocalMux I__12924 (
            .O(N__60094),
            .I(N__60089));
    InMux I__12923 (
            .O(N__60093),
            .I(N__60084));
    InMux I__12922 (
            .O(N__60092),
            .I(N__60084));
    Odrv12 I__12921 (
            .O(N__60089),
            .I(Add_add_temp_7_adj_2413));
    LocalMux I__12920 (
            .O(N__60084),
            .I(Add_add_temp_7_adj_2413));
    CascadeMux I__12919 (
            .O(N__60079),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_ ));
    InMux I__12918 (
            .O(N__60076),
            .I(N__60073));
    LocalMux I__12917 (
            .O(N__60073),
            .I(N__60070));
    Span4Mux_v I__12916 (
            .O(N__60070),
            .I(N__60065));
    InMux I__12915 (
            .O(N__60069),
            .I(N__60060));
    InMux I__12914 (
            .O(N__60068),
            .I(N__60060));
    Odrv4 I__12913 (
            .O(N__60065),
            .I(Add_add_temp_6_adj_2414));
    LocalMux I__12912 (
            .O(N__60060),
            .I(Add_add_temp_6_adj_2414));
    InMux I__12911 (
            .O(N__60055),
            .I(N__60052));
    LocalMux I__12910 (
            .O(N__60052),
            .I(N__60049));
    Span4Mux_h I__12909 (
            .O(N__60049),
            .I(N__60046));
    Odrv4 I__12908 (
            .O(N__60046),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26 ));
    InMux I__12907 (
            .O(N__60043),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15994 ));
    CascadeMux I__12906 (
            .O(N__60040),
            .I(N__60037));
    InMux I__12905 (
            .O(N__60037),
            .I(N__60034));
    LocalMux I__12904 (
            .O(N__60034),
            .I(N__60031));
    Span4Mux_h I__12903 (
            .O(N__60031),
            .I(N__60028));
    Odrv4 I__12902 (
            .O(N__60028),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27 ));
    InMux I__12901 (
            .O(N__60025),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15995 ));
    CascadeMux I__12900 (
            .O(N__60022),
            .I(N__60019));
    InMux I__12899 (
            .O(N__60019),
            .I(N__60016));
    LocalMux I__12898 (
            .O(N__60016),
            .I(N__60013));
    Span4Mux_v I__12897 (
            .O(N__60013),
            .I(N__60010));
    Odrv4 I__12896 (
            .O(N__60010),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28 ));
    InMux I__12895 (
            .O(N__60007),
            .I(N__59998));
    InMux I__12894 (
            .O(N__60006),
            .I(N__59998));
    InMux I__12893 (
            .O(N__60005),
            .I(N__59998));
    LocalMux I__12892 (
            .O(N__59998),
            .I(N__59995));
    Odrv12 I__12891 (
            .O(N__59995),
            .I(Add_add_temp_28));
    InMux I__12890 (
            .O(N__59992),
            .I(bfn_22_22_0_));
    CascadeMux I__12889 (
            .O(N__59989),
            .I(N__59986));
    InMux I__12888 (
            .O(N__59986),
            .I(N__59983));
    LocalMux I__12887 (
            .O(N__59983),
            .I(N__59980));
    Span4Mux_v I__12886 (
            .O(N__59980),
            .I(N__59977));
    Odrv4 I__12885 (
            .O(N__59977),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29 ));
    InMux I__12884 (
            .O(N__59974),
            .I(N__59965));
    InMux I__12883 (
            .O(N__59973),
            .I(N__59965));
    InMux I__12882 (
            .O(N__59972),
            .I(N__59965));
    LocalMux I__12881 (
            .O(N__59965),
            .I(N__59962));
    Span4Mux_v I__12880 (
            .O(N__59962),
            .I(N__59959));
    Odrv4 I__12879 (
            .O(N__59959),
            .I(Add_add_temp_29));
    InMux I__12878 (
            .O(N__59956),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15997 ));
    CascadeMux I__12877 (
            .O(N__59953),
            .I(N__59950));
    InMux I__12876 (
            .O(N__59950),
            .I(N__59947));
    LocalMux I__12875 (
            .O(N__59947),
            .I(N__59944));
    Span4Mux_v I__12874 (
            .O(N__59944),
            .I(N__59941));
    Span4Mux_h I__12873 (
            .O(N__59941),
            .I(N__59938));
    Odrv4 I__12872 (
            .O(N__59938),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30 ));
    InMux I__12871 (
            .O(N__59935),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15998 ));
    InMux I__12870 (
            .O(N__59932),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15999 ));
    InMux I__12869 (
            .O(N__59929),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n16000 ));
    InMux I__12868 (
            .O(N__59926),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n16001 ));
    CascadeMux I__12867 (
            .O(N__59923),
            .I(N__59920));
    InMux I__12866 (
            .O(N__59920),
            .I(N__59917));
    LocalMux I__12865 (
            .O(N__59917),
            .I(N__59914));
    Span4Mux_h I__12864 (
            .O(N__59914),
            .I(N__59911));
    Odrv4 I__12863 (
            .O(N__59911),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17 ));
    InMux I__12862 (
            .O(N__59908),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15985 ));
    CascadeMux I__12861 (
            .O(N__59905),
            .I(N__59902));
    InMux I__12860 (
            .O(N__59902),
            .I(N__59899));
    LocalMux I__12859 (
            .O(N__59899),
            .I(N__59896));
    Span4Mux_h I__12858 (
            .O(N__59896),
            .I(N__59893));
    Odrv4 I__12857 (
            .O(N__59893),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18 ));
    InMux I__12856 (
            .O(N__59890),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15986 ));
    InMux I__12855 (
            .O(N__59887),
            .I(N__59884));
    LocalMux I__12854 (
            .O(N__59884),
            .I(N__59881));
    Span4Mux_h I__12853 (
            .O(N__59881),
            .I(N__59878));
    Odrv4 I__12852 (
            .O(N__59878),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19 ));
    InMux I__12851 (
            .O(N__59875),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15987 ));
    CascadeMux I__12850 (
            .O(N__59872),
            .I(N__59869));
    InMux I__12849 (
            .O(N__59869),
            .I(N__59866));
    LocalMux I__12848 (
            .O(N__59866),
            .I(N__59863));
    Span4Mux_v I__12847 (
            .O(N__59863),
            .I(N__59860));
    Odrv4 I__12846 (
            .O(N__59860),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20 ));
    InMux I__12845 (
            .O(N__59857),
            .I(bfn_22_21_0_));
    CascadeMux I__12844 (
            .O(N__59854),
            .I(N__59851));
    InMux I__12843 (
            .O(N__59851),
            .I(N__59848));
    LocalMux I__12842 (
            .O(N__59848),
            .I(N__59845));
    Span4Mux_v I__12841 (
            .O(N__59845),
            .I(N__59842));
    Odrv4 I__12840 (
            .O(N__59842),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21 ));
    InMux I__12839 (
            .O(N__59839),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15989 ));
    CascadeMux I__12838 (
            .O(N__59836),
            .I(N__59833));
    InMux I__12837 (
            .O(N__59833),
            .I(N__59830));
    LocalMux I__12836 (
            .O(N__59830),
            .I(N__59827));
    Span4Mux_v I__12835 (
            .O(N__59827),
            .I(N__59824));
    Odrv4 I__12834 (
            .O(N__59824),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22 ));
    InMux I__12833 (
            .O(N__59821),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15990 ));
    InMux I__12832 (
            .O(N__59818),
            .I(N__59815));
    LocalMux I__12831 (
            .O(N__59815),
            .I(N__59812));
    Span4Mux_v I__12830 (
            .O(N__59812),
            .I(N__59809));
    Odrv4 I__12829 (
            .O(N__59809),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23 ));
    InMux I__12828 (
            .O(N__59806),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15991 ));
    InMux I__12827 (
            .O(N__59803),
            .I(N__59800));
    LocalMux I__12826 (
            .O(N__59800),
            .I(N__59797));
    Span4Mux_v I__12825 (
            .O(N__59797),
            .I(N__59794));
    Odrv4 I__12824 (
            .O(N__59794),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24 ));
    InMux I__12823 (
            .O(N__59791),
            .I(N__59788));
    LocalMux I__12822 (
            .O(N__59788),
            .I(N__59783));
    InMux I__12821 (
            .O(N__59787),
            .I(N__59778));
    InMux I__12820 (
            .O(N__59786),
            .I(N__59778));
    Span4Mux_h I__12819 (
            .O(N__59783),
            .I(N__59773));
    LocalMux I__12818 (
            .O(N__59778),
            .I(N__59773));
    Odrv4 I__12817 (
            .O(N__59773),
            .I(Add_add_temp_24));
    InMux I__12816 (
            .O(N__59770),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15992 ));
    CascadeMux I__12815 (
            .O(N__59767),
            .I(N__59764));
    InMux I__12814 (
            .O(N__59764),
            .I(N__59761));
    LocalMux I__12813 (
            .O(N__59761),
            .I(N__59758));
    Span4Mux_h I__12812 (
            .O(N__59758),
            .I(N__59755));
    Odrv4 I__12811 (
            .O(N__59755),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25 ));
    InMux I__12810 (
            .O(N__59752),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15993 ));
    CascadeMux I__12809 (
            .O(N__59749),
            .I(N__59746));
    InMux I__12808 (
            .O(N__59746),
            .I(N__59743));
    LocalMux I__12807 (
            .O(N__59743),
            .I(N__59740));
    Odrv4 I__12806 (
            .O(N__59740),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9 ));
    InMux I__12805 (
            .O(N__59737),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15977 ));
    InMux I__12804 (
            .O(N__59734),
            .I(N__59731));
    LocalMux I__12803 (
            .O(N__59731),
            .I(N__59728));
    Odrv12 I__12802 (
            .O(N__59728),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6 ));
    CascadeMux I__12801 (
            .O(N__59725),
            .I(N__59722));
    InMux I__12800 (
            .O(N__59722),
            .I(N__59719));
    LocalMux I__12799 (
            .O(N__59719),
            .I(N__59716));
    Span4Mux_h I__12798 (
            .O(N__59716),
            .I(N__59713));
    Odrv4 I__12797 (
            .O(N__59713),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10 ));
    InMux I__12796 (
            .O(N__59710),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15978 ));
    InMux I__12795 (
            .O(N__59707),
            .I(N__59704));
    LocalMux I__12794 (
            .O(N__59704),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11 ));
    InMux I__12793 (
            .O(N__59701),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15979 ));
    CascadeMux I__12792 (
            .O(N__59698),
            .I(N__59695));
    InMux I__12791 (
            .O(N__59695),
            .I(N__59692));
    LocalMux I__12790 (
            .O(N__59692),
            .I(N__59689));
    Odrv4 I__12789 (
            .O(N__59689),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12 ));
    InMux I__12788 (
            .O(N__59686),
            .I(bfn_22_20_0_));
    CascadeMux I__12787 (
            .O(N__59683),
            .I(N__59680));
    InMux I__12786 (
            .O(N__59680),
            .I(N__59677));
    LocalMux I__12785 (
            .O(N__59677),
            .I(N__59674));
    Odrv4 I__12784 (
            .O(N__59674),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13 ));
    InMux I__12783 (
            .O(N__59671),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15981 ));
    CascadeMux I__12782 (
            .O(N__59668),
            .I(N__59665));
    InMux I__12781 (
            .O(N__59665),
            .I(N__59662));
    LocalMux I__12780 (
            .O(N__59662),
            .I(N__59659));
    Odrv4 I__12779 (
            .O(N__59659),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14 ));
    InMux I__12778 (
            .O(N__59656),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15982 ));
    InMux I__12777 (
            .O(N__59653),
            .I(N__59650));
    LocalMux I__12776 (
            .O(N__59650),
            .I(N__59647));
    Odrv4 I__12775 (
            .O(N__59647),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15 ));
    InMux I__12774 (
            .O(N__59644),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15983 ));
    CascadeMux I__12773 (
            .O(N__59641),
            .I(N__59638));
    InMux I__12772 (
            .O(N__59638),
            .I(N__59635));
    LocalMux I__12771 (
            .O(N__59635),
            .I(N__59632));
    Span4Mux_v I__12770 (
            .O(N__59632),
            .I(N__59629));
    Span4Mux_h I__12769 (
            .O(N__59629),
            .I(N__59626));
    Odrv4 I__12768 (
            .O(N__59626),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16 ));
    InMux I__12767 (
            .O(N__59623),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15984 ));
    CascadeMux I__12766 (
            .O(N__59620),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_ ));
    CascadeMux I__12765 (
            .O(N__59617),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_ ));
    InMux I__12764 (
            .O(N__59614),
            .I(N__59611));
    LocalMux I__12763 (
            .O(N__59611),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20634 ));
    InMux I__12762 (
            .O(N__59608),
            .I(N__59605));
    LocalMux I__12761 (
            .O(N__59605),
            .I(N__59602));
    Odrv4 I__12760 (
            .O(N__59602),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0 ));
    CascadeMux I__12759 (
            .O(N__59599),
            .I(N__59596));
    InMux I__12758 (
            .O(N__59596),
            .I(N__59593));
    LocalMux I__12757 (
            .O(N__59593),
            .I(N__59590));
    Odrv4 I__12756 (
            .O(N__59590),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4 ));
    InMux I__12755 (
            .O(N__59587),
            .I(N__59584));
    LocalMux I__12754 (
            .O(N__59584),
            .I(N__59581));
    Odrv4 I__12753 (
            .O(N__59581),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1 ));
    CascadeMux I__12752 (
            .O(N__59578),
            .I(N__59575));
    InMux I__12751 (
            .O(N__59575),
            .I(N__59572));
    LocalMux I__12750 (
            .O(N__59572),
            .I(N__59569));
    Span4Mux_v I__12749 (
            .O(N__59569),
            .I(N__59566));
    Odrv4 I__12748 (
            .O(N__59566),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5 ));
    InMux I__12747 (
            .O(N__59563),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15973 ));
    InMux I__12746 (
            .O(N__59560),
            .I(N__59557));
    LocalMux I__12745 (
            .O(N__59557),
            .I(N__59554));
    Odrv4 I__12744 (
            .O(N__59554),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2 ));
    CascadeMux I__12743 (
            .O(N__59551),
            .I(N__59548));
    InMux I__12742 (
            .O(N__59548),
            .I(N__59545));
    LocalMux I__12741 (
            .O(N__59545),
            .I(N__59542));
    Odrv4 I__12740 (
            .O(N__59542),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6 ));
    InMux I__12739 (
            .O(N__59539),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15974 ));
    InMux I__12738 (
            .O(N__59536),
            .I(N__59533));
    LocalMux I__12737 (
            .O(N__59533),
            .I(N__59530));
    Odrv4 I__12736 (
            .O(N__59530),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3 ));
    CascadeMux I__12735 (
            .O(N__59527),
            .I(N__59524));
    InMux I__12734 (
            .O(N__59524),
            .I(N__59521));
    LocalMux I__12733 (
            .O(N__59521),
            .I(N__59518));
    Span4Mux_v I__12732 (
            .O(N__59518),
            .I(N__59515));
    Odrv4 I__12731 (
            .O(N__59515),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7 ));
    InMux I__12730 (
            .O(N__59512),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15975 ));
    CascadeMux I__12729 (
            .O(N__59509),
            .I(N__59506));
    InMux I__12728 (
            .O(N__59506),
            .I(N__59503));
    LocalMux I__12727 (
            .O(N__59503),
            .I(N__59500));
    Span4Mux_v I__12726 (
            .O(N__59500),
            .I(N__59497));
    Odrv4 I__12725 (
            .O(N__59497),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8 ));
    InMux I__12724 (
            .O(N__59494),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15976 ));
    CascadeMux I__12723 (
            .O(N__59491),
            .I(Saturate_out1_31__N_267_cascade_));
    CascadeMux I__12722 (
            .O(N__59488),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_ ));
    CascadeMux I__12721 (
            .O(N__59485),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_ ));
    InMux I__12720 (
            .O(N__59482),
            .I(N__59476));
    InMux I__12719 (
            .O(N__59481),
            .I(N__59476));
    LocalMux I__12718 (
            .O(N__59476),
            .I(N__59473));
    Span4Mux_h I__12717 (
            .O(N__59473),
            .I(N__59470));
    Span4Mux_v I__12716 (
            .O(N__59470),
            .I(N__59467));
    Span4Mux_v I__12715 (
            .O(N__59467),
            .I(N__59462));
    InMux I__12714 (
            .O(N__59466),
            .I(N__59459));
    InMux I__12713 (
            .O(N__59465),
            .I(N__59456));
    Odrv4 I__12712 (
            .O(N__59462),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15 ));
    LocalMux I__12711 (
            .O(N__59459),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15 ));
    LocalMux I__12710 (
            .O(N__59456),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15 ));
    InMux I__12709 (
            .O(N__59449),
            .I(N__59446));
    LocalMux I__12708 (
            .O(N__59446),
            .I(\foc.qVoltage_6 ));
    InMux I__12707 (
            .O(N__59443),
            .I(N__59437));
    InMux I__12706 (
            .O(N__59442),
            .I(N__59434));
    CascadeMux I__12705 (
            .O(N__59441),
            .I(N__59430));
    CascadeMux I__12704 (
            .O(N__59440),
            .I(N__59420));
    LocalMux I__12703 (
            .O(N__59437),
            .I(N__59412));
    LocalMux I__12702 (
            .O(N__59434),
            .I(N__59409));
    InMux I__12701 (
            .O(N__59433),
            .I(N__59402));
    InMux I__12700 (
            .O(N__59430),
            .I(N__59402));
    InMux I__12699 (
            .O(N__59429),
            .I(N__59402));
    InMux I__12698 (
            .O(N__59428),
            .I(N__59391));
    InMux I__12697 (
            .O(N__59427),
            .I(N__59391));
    InMux I__12696 (
            .O(N__59426),
            .I(N__59391));
    InMux I__12695 (
            .O(N__59425),
            .I(N__59391));
    InMux I__12694 (
            .O(N__59424),
            .I(N__59391));
    InMux I__12693 (
            .O(N__59423),
            .I(N__59388));
    InMux I__12692 (
            .O(N__59420),
            .I(N__59381));
    InMux I__12691 (
            .O(N__59419),
            .I(N__59381));
    InMux I__12690 (
            .O(N__59418),
            .I(N__59381));
    InMux I__12689 (
            .O(N__59417),
            .I(N__59374));
    InMux I__12688 (
            .O(N__59416),
            .I(N__59374));
    InMux I__12687 (
            .O(N__59415),
            .I(N__59374));
    Odrv4 I__12686 (
            .O(N__59412),
            .I(\foc.Out_31__N_332 ));
    Odrv4 I__12685 (
            .O(N__59409),
            .I(\foc.Out_31__N_332 ));
    LocalMux I__12684 (
            .O(N__59402),
            .I(\foc.Out_31__N_332 ));
    LocalMux I__12683 (
            .O(N__59391),
            .I(\foc.Out_31__N_332 ));
    LocalMux I__12682 (
            .O(N__59388),
            .I(\foc.Out_31__N_332 ));
    LocalMux I__12681 (
            .O(N__59381),
            .I(\foc.Out_31__N_332 ));
    LocalMux I__12680 (
            .O(N__59374),
            .I(\foc.Out_31__N_332 ));
    InMux I__12679 (
            .O(N__59359),
            .I(N__59355));
    InMux I__12678 (
            .O(N__59358),
            .I(N__59352));
    LocalMux I__12677 (
            .O(N__59355),
            .I(N__59345));
    LocalMux I__12676 (
            .O(N__59352),
            .I(N__59345));
    InMux I__12675 (
            .O(N__59351),
            .I(N__59342));
    InMux I__12674 (
            .O(N__59350),
            .I(N__59339));
    Span12Mux_v I__12673 (
            .O(N__59345),
            .I(N__59336));
    LocalMux I__12672 (
            .O(N__59342),
            .I(N__59331));
    LocalMux I__12671 (
            .O(N__59339),
            .I(N__59331));
    Odrv12 I__12670 (
            .O(N__59336),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21 ));
    Odrv12 I__12669 (
            .O(N__59331),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21 ));
    CascadeMux I__12668 (
            .O(N__59326),
            .I(N__59322));
    InMux I__12667 (
            .O(N__59325),
            .I(N__59319));
    InMux I__12666 (
            .O(N__59322),
            .I(N__59316));
    LocalMux I__12665 (
            .O(N__59319),
            .I(N__59312));
    LocalMux I__12664 (
            .O(N__59316),
            .I(N__59309));
    CascadeMux I__12663 (
            .O(N__59315),
            .I(N__59301));
    Span12Mux_s11_h I__12662 (
            .O(N__59312),
            .I(N__59287));
    Sp12to4 I__12661 (
            .O(N__59309),
            .I(N__59287));
    InMux I__12660 (
            .O(N__59308),
            .I(N__59280));
    InMux I__12659 (
            .O(N__59307),
            .I(N__59280));
    InMux I__12658 (
            .O(N__59306),
            .I(N__59280));
    InMux I__12657 (
            .O(N__59305),
            .I(N__59269));
    InMux I__12656 (
            .O(N__59304),
            .I(N__59269));
    InMux I__12655 (
            .O(N__59301),
            .I(N__59269));
    InMux I__12654 (
            .O(N__59300),
            .I(N__59269));
    InMux I__12653 (
            .O(N__59299),
            .I(N__59269));
    InMux I__12652 (
            .O(N__59298),
            .I(N__59266));
    InMux I__12651 (
            .O(N__59297),
            .I(N__59259));
    InMux I__12650 (
            .O(N__59296),
            .I(N__59259));
    InMux I__12649 (
            .O(N__59295),
            .I(N__59259));
    InMux I__12648 (
            .O(N__59294),
            .I(N__59252));
    InMux I__12647 (
            .O(N__59293),
            .I(N__59252));
    InMux I__12646 (
            .O(N__59292),
            .I(N__59252));
    Odrv12 I__12645 (
            .O(N__59287),
            .I(\foc.Out_31__N_333 ));
    LocalMux I__12644 (
            .O(N__59280),
            .I(\foc.Out_31__N_333 ));
    LocalMux I__12643 (
            .O(N__59269),
            .I(\foc.Out_31__N_333 ));
    LocalMux I__12642 (
            .O(N__59266),
            .I(\foc.Out_31__N_333 ));
    LocalMux I__12641 (
            .O(N__59259),
            .I(\foc.Out_31__N_333 ));
    LocalMux I__12640 (
            .O(N__59252),
            .I(\foc.Out_31__N_333 ));
    InMux I__12639 (
            .O(N__59239),
            .I(N__59236));
    LocalMux I__12638 (
            .O(N__59236),
            .I(\foc.qVoltage_12 ));
    CascadeMux I__12637 (
            .O(N__59233),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_ ));
    CascadeMux I__12636 (
            .O(N__59230),
            .I(\foc.Out_31__N_333_adj_2310_cascade_ ));
    InMux I__12635 (
            .O(N__59227),
            .I(N__59224));
    LocalMux I__12634 (
            .O(N__59224),
            .I(\foc.dVoltage_14 ));
    CascadeMux I__12633 (
            .O(N__59221),
            .I(\foc.dVoltage_3_cascade_ ));
    InMux I__12632 (
            .O(N__59218),
            .I(N__59215));
    LocalMux I__12631 (
            .O(N__59215),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20572 ));
    CascadeMux I__12630 (
            .O(N__59212),
            .I(\foc.dVoltage_11_cascade_ ));
    InMux I__12629 (
            .O(N__59209),
            .I(N__59206));
    LocalMux I__12628 (
            .O(N__59206),
            .I(\foc.dVoltage_9 ));
    InMux I__12627 (
            .O(N__59203),
            .I(N__59200));
    LocalMux I__12626 (
            .O(N__59200),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20566 ));
    InMux I__12625 (
            .O(N__59197),
            .I(N__59191));
    InMux I__12624 (
            .O(N__59196),
            .I(N__59191));
    LocalMux I__12623 (
            .O(N__59191),
            .I(N__59188));
    Span4Mux_h I__12622 (
            .O(N__59188),
            .I(N__59185));
    Span4Mux_v I__12621 (
            .O(N__59185),
            .I(N__59182));
    Span4Mux_v I__12620 (
            .O(N__59182),
            .I(N__59177));
    InMux I__12619 (
            .O(N__59181),
            .I(N__59174));
    InMux I__12618 (
            .O(N__59180),
            .I(N__59171));
    Odrv4 I__12617 (
            .O(N__59177),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11 ));
    LocalMux I__12616 (
            .O(N__59174),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11 ));
    LocalMux I__12615 (
            .O(N__59171),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11 ));
    CascadeMux I__12614 (
            .O(N__59164),
            .I(\foc.qVoltage_2_cascade_ ));
    InMux I__12613 (
            .O(N__59161),
            .I(N__59158));
    LocalMux I__12612 (
            .O(N__59158),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20594 ));
    InMux I__12611 (
            .O(N__59155),
            .I(N__59152));
    LocalMux I__12610 (
            .O(N__59152),
            .I(N__59147));
    InMux I__12609 (
            .O(N__59151),
            .I(N__59144));
    InMux I__12608 (
            .O(N__59150),
            .I(N__59141));
    Span12Mux_h I__12607 (
            .O(N__59147),
            .I(N__59134));
    LocalMux I__12606 (
            .O(N__59144),
            .I(N__59134));
    LocalMux I__12605 (
            .O(N__59141),
            .I(N__59134));
    Odrv12 I__12604 (
            .O(N__59134),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20 ));
    CascadeMux I__12603 (
            .O(N__59131),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_ ));
    InMux I__12602 (
            .O(N__59128),
            .I(N__59125));
    LocalMux I__12601 (
            .O(N__59125),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20612 ));
    InMux I__12600 (
            .O(N__59122),
            .I(N__59119));
    LocalMux I__12599 (
            .O(N__59119),
            .I(N__59116));
    Span4Mux_h I__12598 (
            .O(N__59116),
            .I(N__59113));
    Span4Mux_v I__12597 (
            .O(N__59113),
            .I(N__59110));
    Odrv4 I__12596 (
            .O(N__59110),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20618 ));
    CascadeMux I__12595 (
            .O(N__59107),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_ ));
    InMux I__12594 (
            .O(N__59104),
            .I(N__59101));
    LocalMux I__12593 (
            .O(N__59101),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20556 ));
    CascadeMux I__12592 (
            .O(N__59098),
            .I(\foc.dVoltage_5_cascade_ ));
    InMux I__12591 (
            .O(N__59095),
            .I(N__59092));
    LocalMux I__12590 (
            .O(N__59092),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20554 ));
    CascadeMux I__12589 (
            .O(N__59089),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_ ));
    InMux I__12588 (
            .O(N__59086),
            .I(N__59083));
    LocalMux I__12587 (
            .O(N__59083),
            .I(\foc.dVoltage_12 ));
    InMux I__12586 (
            .O(N__59080),
            .I(N__59077));
    LocalMux I__12585 (
            .O(N__59077),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20560 ));
    CascadeMux I__12584 (
            .O(N__59074),
            .I(\foc.Out_31__N_332_adj_2312_cascade_ ));
    InMux I__12583 (
            .O(N__59071),
            .I(N__59068));
    LocalMux I__12582 (
            .O(N__59068),
            .I(\foc.dVoltage_8 ));
    InMux I__12581 (
            .O(N__59065),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17542 ));
    InMux I__12580 (
            .O(N__59062),
            .I(N__59059));
    LocalMux I__12579 (
            .O(N__59059),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n400 ));
    InMux I__12578 (
            .O(N__59056),
            .I(bfn_22_12_0_));
    CascadeMux I__12577 (
            .O(N__59053),
            .I(N__59050));
    InMux I__12576 (
            .O(N__59050),
            .I(N__59047));
    LocalMux I__12575 (
            .O(N__59047),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n449 ));
    InMux I__12574 (
            .O(N__59044),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17544 ));
    InMux I__12573 (
            .O(N__59041),
            .I(N__59038));
    LocalMux I__12572 (
            .O(N__59038),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n498 ));
    InMux I__12571 (
            .O(N__59035),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17545 ));
    CascadeMux I__12570 (
            .O(N__59032),
            .I(N__59029));
    InMux I__12569 (
            .O(N__59029),
            .I(N__59026));
    LocalMux I__12568 (
            .O(N__59026),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n547 ));
    InMux I__12567 (
            .O(N__59023),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17546 ));
    InMux I__12566 (
            .O(N__59020),
            .I(N__59017));
    LocalMux I__12565 (
            .O(N__59017),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n596 ));
    InMux I__12564 (
            .O(N__59014),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17547 ));
    CascadeMux I__12563 (
            .O(N__59011),
            .I(N__59008));
    InMux I__12562 (
            .O(N__59008),
            .I(N__59005));
    LocalMux I__12561 (
            .O(N__59005),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n645 ));
    InMux I__12560 (
            .O(N__59002),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17548 ));
    InMux I__12559 (
            .O(N__58999),
            .I(N__58996));
    LocalMux I__12558 (
            .O(N__58996),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n694 ));
    CascadeMux I__12557 (
            .O(N__58993),
            .I(N__58990));
    InMux I__12556 (
            .O(N__58990),
            .I(N__58987));
    LocalMux I__12555 (
            .O(N__58987),
            .I(N__58984));
    Span4Mux_h I__12554 (
            .O(N__58984),
            .I(N__58980));
    InMux I__12553 (
            .O(N__58983),
            .I(N__58977));
    Span4Mux_v I__12552 (
            .O(N__58980),
            .I(N__58972));
    LocalMux I__12551 (
            .O(N__58977),
            .I(N__58972));
    Span4Mux_h I__12550 (
            .O(N__58972),
            .I(N__58969));
    Odrv4 I__12549 (
            .O(N__58969),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n741 ));
    InMux I__12548 (
            .O(N__58966),
            .I(N__58963));
    LocalMux I__12547 (
            .O(N__58963),
            .I(N__58960));
    Span12Mux_v I__12546 (
            .O(N__58960),
            .I(N__58957));
    Odrv12 I__12545 (
            .O(N__58957),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411 ));
    InMux I__12544 (
            .O(N__58954),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17549 ));
    InMux I__12543 (
            .O(N__58951),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410 ));
    InMux I__12542 (
            .O(N__58948),
            .I(N__58945));
    LocalMux I__12541 (
            .O(N__58945),
            .I(N__58942));
    Span4Mux_v I__12540 (
            .O(N__58942),
            .I(N__58939));
    Odrv4 I__12539 (
            .O(N__58939),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO ));
    InMux I__12538 (
            .O(N__58936),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590 ));
    CascadeMux I__12537 (
            .O(N__58933),
            .I(N__58930));
    InMux I__12536 (
            .O(N__58930),
            .I(N__58927));
    LocalMux I__12535 (
            .O(N__58927),
            .I(N__58924));
    Span4Mux_v I__12534 (
            .O(N__58924),
            .I(N__58921));
    Span4Mux_v I__12533 (
            .O(N__58921),
            .I(N__58918));
    Odrv4 I__12532 (
            .O(N__58918),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO ));
    CascadeMux I__12531 (
            .O(N__58915),
            .I(N__58912));
    InMux I__12530 (
            .O(N__58912),
            .I(N__58896));
    CascadeMux I__12529 (
            .O(N__58911),
            .I(N__58892));
    CascadeMux I__12528 (
            .O(N__58910),
            .I(N__58888));
    CascadeMux I__12527 (
            .O(N__58909),
            .I(N__58884));
    CascadeMux I__12526 (
            .O(N__58908),
            .I(N__58881));
    CascadeMux I__12525 (
            .O(N__58907),
            .I(N__58878));
    CascadeMux I__12524 (
            .O(N__58906),
            .I(N__58875));
    CascadeMux I__12523 (
            .O(N__58905),
            .I(N__58871));
    CascadeMux I__12522 (
            .O(N__58904),
            .I(N__58867));
    CascadeMux I__12521 (
            .O(N__58903),
            .I(N__58861));
    CascadeMux I__12520 (
            .O(N__58902),
            .I(N__58857));
    CascadeMux I__12519 (
            .O(N__58901),
            .I(N__58853));
    CascadeMux I__12518 (
            .O(N__58900),
            .I(N__58849));
    CascadeMux I__12517 (
            .O(N__58899),
            .I(N__58846));
    LocalMux I__12516 (
            .O(N__58896),
            .I(N__58842));
    InMux I__12515 (
            .O(N__58895),
            .I(N__58829));
    InMux I__12514 (
            .O(N__58892),
            .I(N__58829));
    InMux I__12513 (
            .O(N__58891),
            .I(N__58829));
    InMux I__12512 (
            .O(N__58888),
            .I(N__58829));
    InMux I__12511 (
            .O(N__58887),
            .I(N__58829));
    InMux I__12510 (
            .O(N__58884),
            .I(N__58829));
    InMux I__12509 (
            .O(N__58881),
            .I(N__58826));
    InMux I__12508 (
            .O(N__58878),
            .I(N__58823));
    InMux I__12507 (
            .O(N__58875),
            .I(N__58820));
    CascadeMux I__12506 (
            .O(N__58874),
            .I(N__58817));
    InMux I__12505 (
            .O(N__58871),
            .I(N__58814));
    CascadeMux I__12504 (
            .O(N__58870),
            .I(N__58811));
    InMux I__12503 (
            .O(N__58867),
            .I(N__58807));
    InMux I__12502 (
            .O(N__58866),
            .I(N__58804));
    InMux I__12501 (
            .O(N__58865),
            .I(N__58801));
    InMux I__12500 (
            .O(N__58864),
            .I(N__58784));
    InMux I__12499 (
            .O(N__58861),
            .I(N__58784));
    InMux I__12498 (
            .O(N__58860),
            .I(N__58784));
    InMux I__12497 (
            .O(N__58857),
            .I(N__58784));
    InMux I__12496 (
            .O(N__58856),
            .I(N__58784));
    InMux I__12495 (
            .O(N__58853),
            .I(N__58784));
    InMux I__12494 (
            .O(N__58852),
            .I(N__58784));
    InMux I__12493 (
            .O(N__58849),
            .I(N__58784));
    InMux I__12492 (
            .O(N__58846),
            .I(N__58781));
    CascadeMux I__12491 (
            .O(N__58845),
            .I(N__58777));
    Span4Mux_v I__12490 (
            .O(N__58842),
            .I(N__58772));
    LocalMux I__12489 (
            .O(N__58829),
            .I(N__58772));
    LocalMux I__12488 (
            .O(N__58826),
            .I(N__58765));
    LocalMux I__12487 (
            .O(N__58823),
            .I(N__58765));
    LocalMux I__12486 (
            .O(N__58820),
            .I(N__58765));
    InMux I__12485 (
            .O(N__58817),
            .I(N__58762));
    LocalMux I__12484 (
            .O(N__58814),
            .I(N__58759));
    InMux I__12483 (
            .O(N__58811),
            .I(N__58756));
    CascadeMux I__12482 (
            .O(N__58810),
            .I(N__58752));
    LocalMux I__12481 (
            .O(N__58807),
            .I(N__58747));
    LocalMux I__12480 (
            .O(N__58804),
            .I(N__58747));
    LocalMux I__12479 (
            .O(N__58801),
            .I(N__58740));
    LocalMux I__12478 (
            .O(N__58784),
            .I(N__58740));
    LocalMux I__12477 (
            .O(N__58781),
            .I(N__58740));
    InMux I__12476 (
            .O(N__58780),
            .I(N__58737));
    InMux I__12475 (
            .O(N__58777),
            .I(N__58734));
    Span4Mux_v I__12474 (
            .O(N__58772),
            .I(N__58731));
    Span4Mux_v I__12473 (
            .O(N__58765),
            .I(N__58722));
    LocalMux I__12472 (
            .O(N__58762),
            .I(N__58722));
    Span4Mux_h I__12471 (
            .O(N__58759),
            .I(N__58722));
    LocalMux I__12470 (
            .O(N__58756),
            .I(N__58722));
    InMux I__12469 (
            .O(N__58755),
            .I(N__58719));
    InMux I__12468 (
            .O(N__58752),
            .I(N__58716));
    Span4Mux_v I__12467 (
            .O(N__58747),
            .I(N__58707));
    Span4Mux_h I__12466 (
            .O(N__58740),
            .I(N__58707));
    LocalMux I__12465 (
            .O(N__58737),
            .I(N__58707));
    LocalMux I__12464 (
            .O(N__58734),
            .I(N__58707));
    Span4Mux_h I__12463 (
            .O(N__58731),
            .I(N__58698));
    Span4Mux_v I__12462 (
            .O(N__58722),
            .I(N__58698));
    LocalMux I__12461 (
            .O(N__58719),
            .I(N__58698));
    LocalMux I__12460 (
            .O(N__58716),
            .I(N__58698));
    Span4Mux_v I__12459 (
            .O(N__58707),
            .I(N__58695));
    Span4Mux_v I__12458 (
            .O(N__58698),
            .I(N__58692));
    Odrv4 I__12457 (
            .O(N__58695),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n105 ));
    Odrv4 I__12456 (
            .O(N__58692),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n105 ));
    CascadeMux I__12455 (
            .O(N__58687),
            .I(N__58684));
    InMux I__12454 (
            .O(N__58684),
            .I(N__58681));
    LocalMux I__12453 (
            .O(N__58681),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491 ));
    InMux I__12452 (
            .O(N__58678),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17536 ));
    InMux I__12451 (
            .O(N__58675),
            .I(N__58672));
    LocalMux I__12450 (
            .O(N__58672),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509 ));
    InMux I__12449 (
            .O(N__58669),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17537 ));
    CascadeMux I__12448 (
            .O(N__58666),
            .I(N__58663));
    InMux I__12447 (
            .O(N__58663),
            .I(N__58660));
    LocalMux I__12446 (
            .O(N__58660),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n155 ));
    InMux I__12445 (
            .O(N__58657),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17538 ));
    InMux I__12444 (
            .O(N__58654),
            .I(N__58651));
    LocalMux I__12443 (
            .O(N__58651),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n204 ));
    InMux I__12442 (
            .O(N__58648),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17539 ));
    CascadeMux I__12441 (
            .O(N__58645),
            .I(N__58642));
    InMux I__12440 (
            .O(N__58642),
            .I(N__58639));
    LocalMux I__12439 (
            .O(N__58639),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464 ));
    InMux I__12438 (
            .O(N__58636),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17540 ));
    InMux I__12437 (
            .O(N__58633),
            .I(N__58630));
    LocalMux I__12436 (
            .O(N__58630),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n302 ));
    InMux I__12435 (
            .O(N__58627),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17541 ));
    CascadeMux I__12434 (
            .O(N__58624),
            .I(N__58621));
    InMux I__12433 (
            .O(N__58621),
            .I(N__58618));
    LocalMux I__12432 (
            .O(N__58618),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396 ));
    CascadeMux I__12431 (
            .O(N__58615),
            .I(N__58612));
    InMux I__12430 (
            .O(N__58612),
            .I(N__58609));
    LocalMux I__12429 (
            .O(N__58609),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587 ));
    InMux I__12428 (
            .O(N__58606),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18300 ));
    CascadeMux I__12427 (
            .O(N__58603),
            .I(N__58600));
    InMux I__12426 (
            .O(N__58600),
            .I(N__58597));
    LocalMux I__12425 (
            .O(N__58597),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586 ));
    InMux I__12424 (
            .O(N__58594),
            .I(bfn_21_29_0_));
    InMux I__12423 (
            .O(N__58591),
            .I(N__58588));
    LocalMux I__12422 (
            .O(N__58588),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585 ));
    InMux I__12421 (
            .O(N__58585),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18302 ));
    InMux I__12420 (
            .O(N__58582),
            .I(N__58579));
    LocalMux I__12419 (
            .O(N__58579),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584 ));
    InMux I__12418 (
            .O(N__58576),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18303 ));
    InMux I__12417 (
            .O(N__58573),
            .I(N__58570));
    LocalMux I__12416 (
            .O(N__58570),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n571 ));
    InMux I__12415 (
            .O(N__58567),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18304 ));
    InMux I__12414 (
            .O(N__58564),
            .I(N__58561));
    LocalMux I__12413 (
            .O(N__58561),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n620 ));
    InMux I__12412 (
            .O(N__58558),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18305 ));
    CascadeMux I__12411 (
            .O(N__58555),
            .I(N__58552));
    InMux I__12410 (
            .O(N__58552),
            .I(N__58549));
    LocalMux I__12409 (
            .O(N__58549),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n669 ));
    InMux I__12408 (
            .O(N__58546),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18306 ));
    CascadeMux I__12407 (
            .O(N__58543),
            .I(N__58540));
    InMux I__12406 (
            .O(N__58540),
            .I(N__58537));
    LocalMux I__12405 (
            .O(N__58537),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n718 ));
    InMux I__12404 (
            .O(N__58534),
            .I(N__58531));
    LocalMux I__12403 (
            .O(N__58531),
            .I(N__58528));
    Span12Mux_v I__12402 (
            .O(N__58528),
            .I(N__58525));
    Odrv12 I__12401 (
            .O(N__58525),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589 ));
    InMux I__12400 (
            .O(N__58522),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18307 ));
    CascadeMux I__12399 (
            .O(N__58519),
            .I(N__58516));
    InMux I__12398 (
            .O(N__58516),
            .I(N__58513));
    LocalMux I__12397 (
            .O(N__58513),
            .I(N__58509));
    InMux I__12396 (
            .O(N__58512),
            .I(N__58506));
    Sp12to4 I__12395 (
            .O(N__58509),
            .I(N__58503));
    LocalMux I__12394 (
            .O(N__58506),
            .I(N__58500));
    Span12Mux_s11_v I__12393 (
            .O(N__58503),
            .I(N__58497));
    Span12Mux_s11_v I__12392 (
            .O(N__58500),
            .I(N__58494));
    Odrv12 I__12391 (
            .O(N__58497),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30 ));
    Odrv12 I__12390 (
            .O(N__58494),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30 ));
    InMux I__12389 (
            .O(N__58489),
            .I(N__58482));
    InMux I__12388 (
            .O(N__58488),
            .I(N__58482));
    InMux I__12387 (
            .O(N__58487),
            .I(N__58479));
    LocalMux I__12386 (
            .O(N__58482),
            .I(N__58476));
    LocalMux I__12385 (
            .O(N__58479),
            .I(N__58473));
    Span4Mux_h I__12384 (
            .O(N__58476),
            .I(N__58470));
    Span12Mux_h I__12383 (
            .O(N__58473),
            .I(N__58467));
    Span4Mux_v I__12382 (
            .O(N__58470),
            .I(N__58464));
    Odrv12 I__12381 (
            .O(N__58467),
            .I(Add_add_temp_34_adj_2386));
    Odrv4 I__12380 (
            .O(N__58464),
            .I(Add_add_temp_34_adj_2386));
    InMux I__12379 (
            .O(N__58459),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15942 ));
    InMux I__12378 (
            .O(N__58456),
            .I(N__58453));
    LocalMux I__12377 (
            .O(N__58453),
            .I(N__58447));
    CascadeMux I__12376 (
            .O(N__58452),
            .I(N__58443));
    CascadeMux I__12375 (
            .O(N__58451),
            .I(N__58439));
    CascadeMux I__12374 (
            .O(N__58450),
            .I(N__58435));
    Span4Mux_v I__12373 (
            .O(N__58447),
            .I(N__58430));
    InMux I__12372 (
            .O(N__58446),
            .I(N__58415));
    InMux I__12371 (
            .O(N__58443),
            .I(N__58415));
    InMux I__12370 (
            .O(N__58442),
            .I(N__58415));
    InMux I__12369 (
            .O(N__58439),
            .I(N__58415));
    InMux I__12368 (
            .O(N__58438),
            .I(N__58415));
    InMux I__12367 (
            .O(N__58435),
            .I(N__58415));
    InMux I__12366 (
            .O(N__58434),
            .I(N__58415));
    InMux I__12365 (
            .O(N__58433),
            .I(N__58412));
    Odrv4 I__12364 (
            .O(N__58430),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31 ));
    LocalMux I__12363 (
            .O(N__58415),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31 ));
    LocalMux I__12362 (
            .O(N__58412),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31 ));
    CascadeMux I__12361 (
            .O(N__58405),
            .I(N__58400));
    CascadeMux I__12360 (
            .O(N__58404),
            .I(N__58396));
    CascadeMux I__12359 (
            .O(N__58403),
            .I(N__58392));
    InMux I__12358 (
            .O(N__58400),
            .I(N__58381));
    InMux I__12357 (
            .O(N__58399),
            .I(N__58381));
    InMux I__12356 (
            .O(N__58396),
            .I(N__58381));
    InMux I__12355 (
            .O(N__58395),
            .I(N__58381));
    InMux I__12354 (
            .O(N__58392),
            .I(N__58381));
    LocalMux I__12353 (
            .O(N__58381),
            .I(N__58378));
    Span4Mux_v I__12352 (
            .O(N__58378),
            .I(N__58375));
    Odrv4 I__12351 (
            .O(N__58375),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31 ));
    InMux I__12350 (
            .O(N__58372),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15943 ));
    InMux I__12349 (
            .O(N__58369),
            .I(N__58364));
    InMux I__12348 (
            .O(N__58368),
            .I(N__58361));
    InMux I__12347 (
            .O(N__58367),
            .I(N__58358));
    LocalMux I__12346 (
            .O(N__58364),
            .I(N__58353));
    LocalMux I__12345 (
            .O(N__58361),
            .I(N__58353));
    LocalMux I__12344 (
            .O(N__58358),
            .I(N__58350));
    Span4Mux_v I__12343 (
            .O(N__58353),
            .I(N__58347));
    Span4Mux_v I__12342 (
            .O(N__58350),
            .I(N__58344));
    Odrv4 I__12341 (
            .O(N__58347),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31 ));
    Odrv4 I__12340 (
            .O(N__58344),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31 ));
    InMux I__12339 (
            .O(N__58339),
            .I(N__58336));
    LocalMux I__12338 (
            .O(N__58336),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n81 ));
    InMux I__12337 (
            .O(N__58333),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18294 ));
    InMux I__12336 (
            .O(N__58330),
            .I(N__58327));
    LocalMux I__12335 (
            .O(N__58327),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n130 ));
    InMux I__12334 (
            .O(N__58324),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18295 ));
    InMux I__12333 (
            .O(N__58321),
            .I(N__58318));
    LocalMux I__12332 (
            .O(N__58318),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n179 ));
    InMux I__12331 (
            .O(N__58315),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18296 ));
    CascadeMux I__12330 (
            .O(N__58312),
            .I(N__58309));
    InMux I__12329 (
            .O(N__58309),
            .I(N__58306));
    LocalMux I__12328 (
            .O(N__58306),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n228 ));
    InMux I__12327 (
            .O(N__58303),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18297 ));
    InMux I__12326 (
            .O(N__58300),
            .I(N__58297));
    LocalMux I__12325 (
            .O(N__58297),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n277 ));
    InMux I__12324 (
            .O(N__58294),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18298 ));
    CascadeMux I__12323 (
            .O(N__58291),
            .I(N__58288));
    InMux I__12322 (
            .O(N__58288),
            .I(N__58285));
    LocalMux I__12321 (
            .O(N__58285),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588 ));
    InMux I__12320 (
            .O(N__58282),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18299 ));
    InMux I__12319 (
            .O(N__58279),
            .I(N__58275));
    InMux I__12318 (
            .O(N__58278),
            .I(N__58272));
    LocalMux I__12317 (
            .O(N__58275),
            .I(N__58269));
    LocalMux I__12316 (
            .O(N__58272),
            .I(N__58266));
    Span4Mux_v I__12315 (
            .O(N__58269),
            .I(N__58263));
    Span4Mux_h I__12314 (
            .O(N__58266),
            .I(N__58260));
    Odrv4 I__12313 (
            .O(N__58263),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23 ));
    Odrv4 I__12312 (
            .O(N__58260),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23 ));
    CascadeMux I__12311 (
            .O(N__58255),
            .I(N__58252));
    InMux I__12310 (
            .O(N__58252),
            .I(N__58249));
    LocalMux I__12309 (
            .O(N__58249),
            .I(N__58246));
    Span4Mux_h I__12308 (
            .O(N__58246),
            .I(N__58243));
    Odrv4 I__12307 (
            .O(N__58243),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27 ));
    InMux I__12306 (
            .O(N__58240),
            .I(N__58235));
    InMux I__12305 (
            .O(N__58239),
            .I(N__58232));
    InMux I__12304 (
            .O(N__58238),
            .I(N__58229));
    LocalMux I__12303 (
            .O(N__58235),
            .I(N__58222));
    LocalMux I__12302 (
            .O(N__58232),
            .I(N__58222));
    LocalMux I__12301 (
            .O(N__58229),
            .I(N__58222));
    Span4Mux_v I__12300 (
            .O(N__58222),
            .I(N__58219));
    Odrv4 I__12299 (
            .O(N__58219),
            .I(Add_add_temp_27_adj_2393));
    InMux I__12298 (
            .O(N__58216),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15935 ));
    CascadeMux I__12297 (
            .O(N__58213),
            .I(N__58209));
    InMux I__12296 (
            .O(N__58212),
            .I(N__58206));
    InMux I__12295 (
            .O(N__58209),
            .I(N__58203));
    LocalMux I__12294 (
            .O(N__58206),
            .I(N__58200));
    LocalMux I__12293 (
            .O(N__58203),
            .I(N__58197));
    Span4Mux_v I__12292 (
            .O(N__58200),
            .I(N__58194));
    Span4Mux_v I__12291 (
            .O(N__58197),
            .I(N__58191));
    Odrv4 I__12290 (
            .O(N__58194),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24 ));
    Odrv4 I__12289 (
            .O(N__58191),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24 ));
    CascadeMux I__12288 (
            .O(N__58186),
            .I(N__58183));
    InMux I__12287 (
            .O(N__58183),
            .I(N__58180));
    LocalMux I__12286 (
            .O(N__58180),
            .I(N__58177));
    Span4Mux_v I__12285 (
            .O(N__58177),
            .I(N__58174));
    Odrv4 I__12284 (
            .O(N__58174),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28 ));
    InMux I__12283 (
            .O(N__58171),
            .I(N__58164));
    InMux I__12282 (
            .O(N__58170),
            .I(N__58164));
    InMux I__12281 (
            .O(N__58169),
            .I(N__58161));
    LocalMux I__12280 (
            .O(N__58164),
            .I(N__58156));
    LocalMux I__12279 (
            .O(N__58161),
            .I(N__58156));
    Span4Mux_v I__12278 (
            .O(N__58156),
            .I(N__58153));
    Odrv4 I__12277 (
            .O(N__58153),
            .I(Add_add_temp_28_adj_2392));
    InMux I__12276 (
            .O(N__58150),
            .I(bfn_21_26_0_));
    InMux I__12275 (
            .O(N__58147),
            .I(N__58144));
    LocalMux I__12274 (
            .O(N__58144),
            .I(N__58141));
    Span4Mux_h I__12273 (
            .O(N__58141),
            .I(N__58137));
    InMux I__12272 (
            .O(N__58140),
            .I(N__58134));
    Sp12to4 I__12271 (
            .O(N__58137),
            .I(N__58129));
    LocalMux I__12270 (
            .O(N__58134),
            .I(N__58129));
    Odrv12 I__12269 (
            .O(N__58129),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25 ));
    CascadeMux I__12268 (
            .O(N__58126),
            .I(N__58123));
    InMux I__12267 (
            .O(N__58123),
            .I(N__58120));
    LocalMux I__12266 (
            .O(N__58120),
            .I(N__58117));
    Span4Mux_v I__12265 (
            .O(N__58117),
            .I(N__58114));
    Odrv4 I__12264 (
            .O(N__58114),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29 ));
    InMux I__12263 (
            .O(N__58111),
            .I(N__58106));
    InMux I__12262 (
            .O(N__58110),
            .I(N__58101));
    InMux I__12261 (
            .O(N__58109),
            .I(N__58101));
    LocalMux I__12260 (
            .O(N__58106),
            .I(N__58098));
    LocalMux I__12259 (
            .O(N__58101),
            .I(N__58095));
    Sp12to4 I__12258 (
            .O(N__58098),
            .I(N__58092));
    Span4Mux_v I__12257 (
            .O(N__58095),
            .I(N__58089));
    Odrv12 I__12256 (
            .O(N__58092),
            .I(Add_add_temp_29_adj_2391));
    Odrv4 I__12255 (
            .O(N__58089),
            .I(Add_add_temp_29_adj_2391));
    InMux I__12254 (
            .O(N__58084),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15937 ));
    InMux I__12253 (
            .O(N__58081),
            .I(N__58077));
    InMux I__12252 (
            .O(N__58080),
            .I(N__58074));
    LocalMux I__12251 (
            .O(N__58077),
            .I(N__58071));
    LocalMux I__12250 (
            .O(N__58074),
            .I(N__58068));
    Span12Mux_v I__12249 (
            .O(N__58071),
            .I(N__58065));
    Span4Mux_v I__12248 (
            .O(N__58068),
            .I(N__58062));
    Odrv12 I__12247 (
            .O(N__58065),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26 ));
    Odrv4 I__12246 (
            .O(N__58062),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26 ));
    CascadeMux I__12245 (
            .O(N__58057),
            .I(N__58054));
    InMux I__12244 (
            .O(N__58054),
            .I(N__58051));
    LocalMux I__12243 (
            .O(N__58051),
            .I(N__58048));
    Span4Mux_v I__12242 (
            .O(N__58048),
            .I(N__58045));
    Odrv4 I__12241 (
            .O(N__58045),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30 ));
    InMux I__12240 (
            .O(N__58042),
            .I(N__58035));
    InMux I__12239 (
            .O(N__58041),
            .I(N__58035));
    InMux I__12238 (
            .O(N__58040),
            .I(N__58032));
    LocalMux I__12237 (
            .O(N__58035),
            .I(N__58029));
    LocalMux I__12236 (
            .O(N__58032),
            .I(N__58026));
    Span4Mux_v I__12235 (
            .O(N__58029),
            .I(N__58021));
    Span4Mux_v I__12234 (
            .O(N__58026),
            .I(N__58021));
    Odrv4 I__12233 (
            .O(N__58021),
            .I(Add_add_temp_30_adj_2390));
    InMux I__12232 (
            .O(N__58018),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15938 ));
    InMux I__12231 (
            .O(N__58015),
            .I(N__58012));
    LocalMux I__12230 (
            .O(N__58012),
            .I(N__58008));
    CascadeMux I__12229 (
            .O(N__58011),
            .I(N__58005));
    Span4Mux_v I__12228 (
            .O(N__58008),
            .I(N__58002));
    InMux I__12227 (
            .O(N__58005),
            .I(N__57999));
    Span4Mux_h I__12226 (
            .O(N__58002),
            .I(N__57994));
    LocalMux I__12225 (
            .O(N__57999),
            .I(N__57994));
    Span4Mux_v I__12224 (
            .O(N__57994),
            .I(N__57991));
    Odrv4 I__12223 (
            .O(N__57991),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27 ));
    InMux I__12222 (
            .O(N__57988),
            .I(N__57981));
    InMux I__12221 (
            .O(N__57987),
            .I(N__57981));
    InMux I__12220 (
            .O(N__57986),
            .I(N__57978));
    LocalMux I__12219 (
            .O(N__57981),
            .I(N__57973));
    LocalMux I__12218 (
            .O(N__57978),
            .I(N__57973));
    Span4Mux_v I__12217 (
            .O(N__57973),
            .I(N__57970));
    Odrv4 I__12216 (
            .O(N__57970),
            .I(Add_add_temp_31_adj_2389));
    InMux I__12215 (
            .O(N__57967),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15939 ));
    InMux I__12214 (
            .O(N__57964),
            .I(N__57960));
    CascadeMux I__12213 (
            .O(N__57963),
            .I(N__57957));
    LocalMux I__12212 (
            .O(N__57960),
            .I(N__57954));
    InMux I__12211 (
            .O(N__57957),
            .I(N__57951));
    Span4Mux_v I__12210 (
            .O(N__57954),
            .I(N__57948));
    LocalMux I__12209 (
            .O(N__57951),
            .I(N__57945));
    Odrv4 I__12208 (
            .O(N__57948),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28 ));
    Odrv12 I__12207 (
            .O(N__57945),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28 ));
    InMux I__12206 (
            .O(N__57940),
            .I(N__57935));
    InMux I__12205 (
            .O(N__57939),
            .I(N__57932));
    InMux I__12204 (
            .O(N__57938),
            .I(N__57929));
    LocalMux I__12203 (
            .O(N__57935),
            .I(N__57922));
    LocalMux I__12202 (
            .O(N__57932),
            .I(N__57922));
    LocalMux I__12201 (
            .O(N__57929),
            .I(N__57922));
    Span4Mux_v I__12200 (
            .O(N__57922),
            .I(N__57919));
    Odrv4 I__12199 (
            .O(N__57919),
            .I(Add_add_temp_32_adj_2388));
    InMux I__12198 (
            .O(N__57916),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15940 ));
    InMux I__12197 (
            .O(N__57913),
            .I(N__57910));
    LocalMux I__12196 (
            .O(N__57910),
            .I(N__57906));
    InMux I__12195 (
            .O(N__57909),
            .I(N__57903));
    Span4Mux_v I__12194 (
            .O(N__57906),
            .I(N__57898));
    LocalMux I__12193 (
            .O(N__57903),
            .I(N__57898));
    Span4Mux_h I__12192 (
            .O(N__57898),
            .I(N__57895));
    Span4Mux_v I__12191 (
            .O(N__57895),
            .I(N__57892));
    Odrv4 I__12190 (
            .O(N__57892),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29 ));
    CascadeMux I__12189 (
            .O(N__57889),
            .I(N__57884));
    InMux I__12188 (
            .O(N__57888),
            .I(N__57879));
    InMux I__12187 (
            .O(N__57887),
            .I(N__57879));
    InMux I__12186 (
            .O(N__57884),
            .I(N__57876));
    LocalMux I__12185 (
            .O(N__57879),
            .I(N__57871));
    LocalMux I__12184 (
            .O(N__57876),
            .I(N__57871));
    Span12Mux_v I__12183 (
            .O(N__57871),
            .I(N__57868));
    Odrv12 I__12182 (
            .O(N__57868),
            .I(Add_add_temp_33_adj_2387));
    InMux I__12181 (
            .O(N__57865),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15941 ));
    InMux I__12180 (
            .O(N__57862),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15927 ));
    InMux I__12179 (
            .O(N__57859),
            .I(N__57856));
    LocalMux I__12178 (
            .O(N__57856),
            .I(N__57853));
    Span4Mux_h I__12177 (
            .O(N__57853),
            .I(N__57849));
    InMux I__12176 (
            .O(N__57852),
            .I(N__57846));
    Odrv4 I__12175 (
            .O(N__57849),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16 ));
    LocalMux I__12174 (
            .O(N__57846),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16 ));
    CascadeMux I__12173 (
            .O(N__57841),
            .I(N__57838));
    InMux I__12172 (
            .O(N__57838),
            .I(N__57835));
    LocalMux I__12171 (
            .O(N__57835),
            .I(N__57832));
    Span4Mux_v I__12170 (
            .O(N__57832),
            .I(N__57829));
    Span4Mux_h I__12169 (
            .O(N__57829),
            .I(N__57826));
    Odrv4 I__12168 (
            .O(N__57826),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20 ));
    InMux I__12167 (
            .O(N__57823),
            .I(bfn_21_25_0_));
    InMux I__12166 (
            .O(N__57820),
            .I(N__57817));
    LocalMux I__12165 (
            .O(N__57817),
            .I(N__57814));
    Span4Mux_h I__12164 (
            .O(N__57814),
            .I(N__57810));
    InMux I__12163 (
            .O(N__57813),
            .I(N__57807));
    Odrv4 I__12162 (
            .O(N__57810),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17 ));
    LocalMux I__12161 (
            .O(N__57807),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17 ));
    CascadeMux I__12160 (
            .O(N__57802),
            .I(N__57799));
    InMux I__12159 (
            .O(N__57799),
            .I(N__57796));
    LocalMux I__12158 (
            .O(N__57796),
            .I(N__57793));
    Span4Mux_v I__12157 (
            .O(N__57793),
            .I(N__57790));
    Odrv4 I__12156 (
            .O(N__57790),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21 ));
    InMux I__12155 (
            .O(N__57787),
            .I(N__57782));
    InMux I__12154 (
            .O(N__57786),
            .I(N__57779));
    InMux I__12153 (
            .O(N__57785),
            .I(N__57776));
    LocalMux I__12152 (
            .O(N__57782),
            .I(N__57773));
    LocalMux I__12151 (
            .O(N__57779),
            .I(N__57770));
    LocalMux I__12150 (
            .O(N__57776),
            .I(N__57767));
    Span4Mux_v I__12149 (
            .O(N__57773),
            .I(N__57762));
    Span4Mux_h I__12148 (
            .O(N__57770),
            .I(N__57762));
    Span4Mux_h I__12147 (
            .O(N__57767),
            .I(N__57759));
    Odrv4 I__12146 (
            .O(N__57762),
            .I(Add_add_temp_21_adj_2399));
    Odrv4 I__12145 (
            .O(N__57759),
            .I(Add_add_temp_21_adj_2399));
    InMux I__12144 (
            .O(N__57754),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15929 ));
    InMux I__12143 (
            .O(N__57751),
            .I(N__57748));
    LocalMux I__12142 (
            .O(N__57748),
            .I(N__57745));
    Span4Mux_v I__12141 (
            .O(N__57745),
            .I(N__57741));
    InMux I__12140 (
            .O(N__57744),
            .I(N__57738));
    Odrv4 I__12139 (
            .O(N__57741),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18 ));
    LocalMux I__12138 (
            .O(N__57738),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18 ));
    CascadeMux I__12137 (
            .O(N__57733),
            .I(N__57730));
    InMux I__12136 (
            .O(N__57730),
            .I(N__57727));
    LocalMux I__12135 (
            .O(N__57727),
            .I(N__57724));
    Span4Mux_v I__12134 (
            .O(N__57724),
            .I(N__57721));
    Odrv4 I__12133 (
            .O(N__57721),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22 ));
    CascadeMux I__12132 (
            .O(N__57718),
            .I(N__57713));
    InMux I__12131 (
            .O(N__57717),
            .I(N__57710));
    InMux I__12130 (
            .O(N__57716),
            .I(N__57707));
    InMux I__12129 (
            .O(N__57713),
            .I(N__57704));
    LocalMux I__12128 (
            .O(N__57710),
            .I(N__57699));
    LocalMux I__12127 (
            .O(N__57707),
            .I(N__57699));
    LocalMux I__12126 (
            .O(N__57704),
            .I(N__57696));
    Span4Mux_v I__12125 (
            .O(N__57699),
            .I(N__57693));
    Odrv12 I__12124 (
            .O(N__57696),
            .I(Add_add_temp_22_adj_2398));
    Odrv4 I__12123 (
            .O(N__57693),
            .I(Add_add_temp_22_adj_2398));
    InMux I__12122 (
            .O(N__57688),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15930 ));
    InMux I__12121 (
            .O(N__57685),
            .I(N__57681));
    InMux I__12120 (
            .O(N__57684),
            .I(N__57678));
    LocalMux I__12119 (
            .O(N__57681),
            .I(N__57675));
    LocalMux I__12118 (
            .O(N__57678),
            .I(N__57672));
    Span4Mux_h I__12117 (
            .O(N__57675),
            .I(N__57669));
    Span4Mux_h I__12116 (
            .O(N__57672),
            .I(N__57666));
    Sp12to4 I__12115 (
            .O(N__57669),
            .I(N__57661));
    Sp12to4 I__12114 (
            .O(N__57666),
            .I(N__57661));
    Odrv12 I__12113 (
            .O(N__57661),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19 ));
    CascadeMux I__12112 (
            .O(N__57658),
            .I(N__57655));
    InMux I__12111 (
            .O(N__57655),
            .I(N__57652));
    LocalMux I__12110 (
            .O(N__57652),
            .I(N__57649));
    Span4Mux_v I__12109 (
            .O(N__57649),
            .I(N__57646));
    Sp12to4 I__12108 (
            .O(N__57646),
            .I(N__57643));
    Odrv12 I__12107 (
            .O(N__57643),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23 ));
    InMux I__12106 (
            .O(N__57640),
            .I(N__57636));
    InMux I__12105 (
            .O(N__57639),
            .I(N__57632));
    LocalMux I__12104 (
            .O(N__57636),
            .I(N__57629));
    InMux I__12103 (
            .O(N__57635),
            .I(N__57626));
    LocalMux I__12102 (
            .O(N__57632),
            .I(N__57623));
    Span4Mux_h I__12101 (
            .O(N__57629),
            .I(N__57620));
    LocalMux I__12100 (
            .O(N__57626),
            .I(N__57615));
    Span4Mux_h I__12099 (
            .O(N__57623),
            .I(N__57615));
    Span4Mux_v I__12098 (
            .O(N__57620),
            .I(N__57612));
    Span4Mux_v I__12097 (
            .O(N__57615),
            .I(N__57609));
    Odrv4 I__12096 (
            .O(N__57612),
            .I(Add_add_temp_23_adj_2397));
    Odrv4 I__12095 (
            .O(N__57609),
            .I(Add_add_temp_23_adj_2397));
    InMux I__12094 (
            .O(N__57604),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15931 ));
    InMux I__12093 (
            .O(N__57601),
            .I(N__57597));
    InMux I__12092 (
            .O(N__57600),
            .I(N__57594));
    LocalMux I__12091 (
            .O(N__57597),
            .I(N__57591));
    LocalMux I__12090 (
            .O(N__57594),
            .I(N__57588));
    Span4Mux_v I__12089 (
            .O(N__57591),
            .I(N__57585));
    Span4Mux_v I__12088 (
            .O(N__57588),
            .I(N__57582));
    Odrv4 I__12087 (
            .O(N__57585),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20 ));
    Odrv4 I__12086 (
            .O(N__57582),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20 ));
    CascadeMux I__12085 (
            .O(N__57577),
            .I(N__57574));
    InMux I__12084 (
            .O(N__57574),
            .I(N__57571));
    LocalMux I__12083 (
            .O(N__57571),
            .I(N__57568));
    Span4Mux_v I__12082 (
            .O(N__57568),
            .I(N__57565));
    Odrv4 I__12081 (
            .O(N__57565),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24 ));
    InMux I__12080 (
            .O(N__57562),
            .I(N__57558));
    InMux I__12079 (
            .O(N__57561),
            .I(N__57555));
    LocalMux I__12078 (
            .O(N__57558),
            .I(N__57552));
    LocalMux I__12077 (
            .O(N__57555),
            .I(N__57548));
    Span4Mux_v I__12076 (
            .O(N__57552),
            .I(N__57545));
    InMux I__12075 (
            .O(N__57551),
            .I(N__57542));
    Sp12to4 I__12074 (
            .O(N__57548),
            .I(N__57535));
    Sp12to4 I__12073 (
            .O(N__57545),
            .I(N__57535));
    LocalMux I__12072 (
            .O(N__57542),
            .I(N__57535));
    Odrv12 I__12071 (
            .O(N__57535),
            .I(Add_add_temp_24_adj_2396));
    InMux I__12070 (
            .O(N__57532),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15932 ));
    InMux I__12069 (
            .O(N__57529),
            .I(N__57526));
    LocalMux I__12068 (
            .O(N__57526),
            .I(N__57522));
    InMux I__12067 (
            .O(N__57525),
            .I(N__57519));
    Span4Mux_h I__12066 (
            .O(N__57522),
            .I(N__57514));
    LocalMux I__12065 (
            .O(N__57519),
            .I(N__57514));
    Span4Mux_v I__12064 (
            .O(N__57514),
            .I(N__57511));
    Odrv4 I__12063 (
            .O(N__57511),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21 ));
    CascadeMux I__12062 (
            .O(N__57508),
            .I(N__57505));
    InMux I__12061 (
            .O(N__57505),
            .I(N__57502));
    LocalMux I__12060 (
            .O(N__57502),
            .I(N__57499));
    Span4Mux_h I__12059 (
            .O(N__57499),
            .I(N__57496));
    Odrv4 I__12058 (
            .O(N__57496),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25 ));
    InMux I__12057 (
            .O(N__57493),
            .I(N__57488));
    InMux I__12056 (
            .O(N__57492),
            .I(N__57485));
    InMux I__12055 (
            .O(N__57491),
            .I(N__57482));
    LocalMux I__12054 (
            .O(N__57488),
            .I(N__57479));
    LocalMux I__12053 (
            .O(N__57485),
            .I(N__57474));
    LocalMux I__12052 (
            .O(N__57482),
            .I(N__57474));
    Span4Mux_h I__12051 (
            .O(N__57479),
            .I(N__57469));
    Span4Mux_v I__12050 (
            .O(N__57474),
            .I(N__57469));
    Odrv4 I__12049 (
            .O(N__57469),
            .I(Add_add_temp_25_adj_2395));
    InMux I__12048 (
            .O(N__57466),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15933 ));
    CascadeMux I__12047 (
            .O(N__57463),
            .I(N__57460));
    InMux I__12046 (
            .O(N__57460),
            .I(N__57457));
    LocalMux I__12045 (
            .O(N__57457),
            .I(N__57453));
    InMux I__12044 (
            .O(N__57456),
            .I(N__57450));
    Span4Mux_v I__12043 (
            .O(N__57453),
            .I(N__57447));
    LocalMux I__12042 (
            .O(N__57450),
            .I(N__57444));
    Odrv4 I__12041 (
            .O(N__57447),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22 ));
    Odrv12 I__12040 (
            .O(N__57444),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22 ));
    CascadeMux I__12039 (
            .O(N__57439),
            .I(N__57436));
    InMux I__12038 (
            .O(N__57436),
            .I(N__57433));
    LocalMux I__12037 (
            .O(N__57433),
            .I(N__57430));
    Span12Mux_h I__12036 (
            .O(N__57430),
            .I(N__57427));
    Odrv12 I__12035 (
            .O(N__57427),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26 ));
    CascadeMux I__12034 (
            .O(N__57424),
            .I(N__57421));
    InMux I__12033 (
            .O(N__57421),
            .I(N__57416));
    InMux I__12032 (
            .O(N__57420),
            .I(N__57411));
    InMux I__12031 (
            .O(N__57419),
            .I(N__57411));
    LocalMux I__12030 (
            .O(N__57416),
            .I(N__57408));
    LocalMux I__12029 (
            .O(N__57411),
            .I(N__57405));
    Span4Mux_h I__12028 (
            .O(N__57408),
            .I(N__57402));
    Span4Mux_v I__12027 (
            .O(N__57405),
            .I(N__57399));
    Span4Mux_v I__12026 (
            .O(N__57402),
            .I(N__57396));
    Span4Mux_h I__12025 (
            .O(N__57399),
            .I(N__57393));
    Odrv4 I__12024 (
            .O(N__57396),
            .I(Add_add_temp_26_adj_2394));
    Odrv4 I__12023 (
            .O(N__57393),
            .I(Add_add_temp_26_adj_2394));
    InMux I__12022 (
            .O(N__57388),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15934 ));
    InMux I__12021 (
            .O(N__57385),
            .I(N__57381));
    InMux I__12020 (
            .O(N__57384),
            .I(N__57378));
    LocalMux I__12019 (
            .O(N__57381),
            .I(N__57375));
    LocalMux I__12018 (
            .O(N__57378),
            .I(N__57372));
    Odrv4 I__12017 (
            .O(N__57375),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8 ));
    Odrv12 I__12016 (
            .O(N__57372),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8 ));
    CascadeMux I__12015 (
            .O(N__57367),
            .I(N__57364));
    InMux I__12014 (
            .O(N__57364),
            .I(N__57361));
    LocalMux I__12013 (
            .O(N__57361),
            .I(N__57358));
    Span4Mux_v I__12012 (
            .O(N__57358),
            .I(N__57355));
    Odrv4 I__12011 (
            .O(N__57355),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12 ));
    InMux I__12010 (
            .O(N__57352),
            .I(bfn_21_24_0_));
    InMux I__12009 (
            .O(N__57349),
            .I(N__57346));
    LocalMux I__12008 (
            .O(N__57346),
            .I(N__57343));
    Odrv12 I__12007 (
            .O(N__57343),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13 ));
    CascadeMux I__12006 (
            .O(N__57340),
            .I(N__57337));
    InMux I__12005 (
            .O(N__57337),
            .I(N__57334));
    LocalMux I__12004 (
            .O(N__57334),
            .I(N__57330));
    InMux I__12003 (
            .O(N__57333),
            .I(N__57327));
    Span4Mux_v I__12002 (
            .O(N__57330),
            .I(N__57324));
    LocalMux I__12001 (
            .O(N__57327),
            .I(N__57321));
    Odrv4 I__12000 (
            .O(N__57324),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9 ));
    Odrv4 I__11999 (
            .O(N__57321),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9 ));
    InMux I__11998 (
            .O(N__57316),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15921 ));
    InMux I__11997 (
            .O(N__57313),
            .I(N__57310));
    LocalMux I__11996 (
            .O(N__57310),
            .I(N__57307));
    Odrv4 I__11995 (
            .O(N__57307),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14 ));
    CascadeMux I__11994 (
            .O(N__57304),
            .I(N__57301));
    InMux I__11993 (
            .O(N__57301),
            .I(N__57298));
    LocalMux I__11992 (
            .O(N__57298),
            .I(N__57294));
    InMux I__11991 (
            .O(N__57297),
            .I(N__57291));
    Span4Mux_v I__11990 (
            .O(N__57294),
            .I(N__57288));
    LocalMux I__11989 (
            .O(N__57291),
            .I(N__57285));
    Odrv4 I__11988 (
            .O(N__57288),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10 ));
    Odrv4 I__11987 (
            .O(N__57285),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10 ));
    InMux I__11986 (
            .O(N__57280),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15922 ));
    InMux I__11985 (
            .O(N__57277),
            .I(N__57273));
    CascadeMux I__11984 (
            .O(N__57276),
            .I(N__57270));
    LocalMux I__11983 (
            .O(N__57273),
            .I(N__57267));
    InMux I__11982 (
            .O(N__57270),
            .I(N__57264));
    Span4Mux_v I__11981 (
            .O(N__57267),
            .I(N__57261));
    LocalMux I__11980 (
            .O(N__57264),
            .I(N__57258));
    Odrv4 I__11979 (
            .O(N__57261),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11 ));
    Odrv4 I__11978 (
            .O(N__57258),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11 ));
    CascadeMux I__11977 (
            .O(N__57253),
            .I(N__57250));
    InMux I__11976 (
            .O(N__57250),
            .I(N__57247));
    LocalMux I__11975 (
            .O(N__57247),
            .I(N__57244));
    Span4Mux_h I__11974 (
            .O(N__57244),
            .I(N__57241));
    Odrv4 I__11973 (
            .O(N__57241),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15 ));
    InMux I__11972 (
            .O(N__57238),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15923 ));
    InMux I__11971 (
            .O(N__57235),
            .I(N__57232));
    LocalMux I__11970 (
            .O(N__57232),
            .I(N__57229));
    Span4Mux_v I__11969 (
            .O(N__57229),
            .I(N__57226));
    Odrv4 I__11968 (
            .O(N__57226),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16 ));
    CascadeMux I__11967 (
            .O(N__57223),
            .I(N__57220));
    InMux I__11966 (
            .O(N__57220),
            .I(N__57216));
    InMux I__11965 (
            .O(N__57219),
            .I(N__57213));
    LocalMux I__11964 (
            .O(N__57216),
            .I(N__57210));
    LocalMux I__11963 (
            .O(N__57213),
            .I(N__57207));
    Odrv4 I__11962 (
            .O(N__57210),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12 ));
    Odrv12 I__11961 (
            .O(N__57207),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12 ));
    InMux I__11960 (
            .O(N__57202),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15924 ));
    InMux I__11959 (
            .O(N__57199),
            .I(N__57196));
    LocalMux I__11958 (
            .O(N__57196),
            .I(N__57192));
    InMux I__11957 (
            .O(N__57195),
            .I(N__57189));
    Span12Mux_s10_v I__11956 (
            .O(N__57192),
            .I(N__57186));
    LocalMux I__11955 (
            .O(N__57189),
            .I(N__57183));
    Odrv12 I__11954 (
            .O(N__57186),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13 ));
    Odrv12 I__11953 (
            .O(N__57183),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13 ));
    CascadeMux I__11952 (
            .O(N__57178),
            .I(N__57175));
    InMux I__11951 (
            .O(N__57175),
            .I(N__57172));
    LocalMux I__11950 (
            .O(N__57172),
            .I(N__57169));
    Span4Mux_h I__11949 (
            .O(N__57169),
            .I(N__57166));
    Odrv4 I__11948 (
            .O(N__57166),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17 ));
    InMux I__11947 (
            .O(N__57163),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15925 ));
    InMux I__11946 (
            .O(N__57160),
            .I(N__57157));
    LocalMux I__11945 (
            .O(N__57157),
            .I(N__57154));
    Span4Mux_h I__11944 (
            .O(N__57154),
            .I(N__57150));
    InMux I__11943 (
            .O(N__57153),
            .I(N__57147));
    Span4Mux_v I__11942 (
            .O(N__57150),
            .I(N__57144));
    LocalMux I__11941 (
            .O(N__57147),
            .I(N__57141));
    Odrv4 I__11940 (
            .O(N__57144),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14 ));
    Odrv4 I__11939 (
            .O(N__57141),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14 ));
    CascadeMux I__11938 (
            .O(N__57136),
            .I(N__57133));
    InMux I__11937 (
            .O(N__57133),
            .I(N__57130));
    LocalMux I__11936 (
            .O(N__57130),
            .I(N__57127));
    Span4Mux_h I__11935 (
            .O(N__57127),
            .I(N__57124));
    Odrv4 I__11934 (
            .O(N__57124),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18 ));
    InMux I__11933 (
            .O(N__57121),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15926 ));
    InMux I__11932 (
            .O(N__57118),
            .I(N__57115));
    LocalMux I__11931 (
            .O(N__57115),
            .I(N__57111));
    InMux I__11930 (
            .O(N__57114),
            .I(N__57108));
    Span4Mux_h I__11929 (
            .O(N__57111),
            .I(N__57103));
    LocalMux I__11928 (
            .O(N__57108),
            .I(N__57103));
    Span4Mux_v I__11927 (
            .O(N__57103),
            .I(N__57100));
    Odrv4 I__11926 (
            .O(N__57100),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15 ));
    CascadeMux I__11925 (
            .O(N__57097),
            .I(N__57094));
    InMux I__11924 (
            .O(N__57094),
            .I(N__57091));
    LocalMux I__11923 (
            .O(N__57091),
            .I(N__57088));
    Span4Mux_h I__11922 (
            .O(N__57088),
            .I(N__57085));
    Odrv4 I__11921 (
            .O(N__57085),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19 ));
    InMux I__11920 (
            .O(N__57082),
            .I(N__57079));
    LocalMux I__11919 (
            .O(N__57079),
            .I(N__57076));
    Odrv12 I__11918 (
            .O(N__57076),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0 ));
    CascadeMux I__11917 (
            .O(N__57073),
            .I(N__57070));
    InMux I__11916 (
            .O(N__57070),
            .I(N__57067));
    LocalMux I__11915 (
            .O(N__57067),
            .I(N__57064));
    Odrv4 I__11914 (
            .O(N__57064),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4 ));
    InMux I__11913 (
            .O(N__57061),
            .I(N__57058));
    LocalMux I__11912 (
            .O(N__57058),
            .I(N__57055));
    Odrv12 I__11911 (
            .O(N__57055),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5 ));
    CascadeMux I__11910 (
            .O(N__57052),
            .I(N__57049));
    InMux I__11909 (
            .O(N__57049),
            .I(N__57046));
    LocalMux I__11908 (
            .O(N__57046),
            .I(N__57043));
    Odrv12 I__11907 (
            .O(N__57043),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1 ));
    InMux I__11906 (
            .O(N__57040),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15913 ));
    InMux I__11905 (
            .O(N__57037),
            .I(N__57034));
    LocalMux I__11904 (
            .O(N__57034),
            .I(N__57031));
    Odrv4 I__11903 (
            .O(N__57031),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2 ));
    CascadeMux I__11902 (
            .O(N__57028),
            .I(N__57025));
    InMux I__11901 (
            .O(N__57025),
            .I(N__57022));
    LocalMux I__11900 (
            .O(N__57022),
            .I(N__57019));
    Span4Mux_v I__11899 (
            .O(N__57019),
            .I(N__57016));
    Odrv4 I__11898 (
            .O(N__57016),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6 ));
    InMux I__11897 (
            .O(N__57013),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15914 ));
    InMux I__11896 (
            .O(N__57010),
            .I(N__57007));
    LocalMux I__11895 (
            .O(N__57007),
            .I(N__57004));
    Odrv12 I__11894 (
            .O(N__57004),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3 ));
    CascadeMux I__11893 (
            .O(N__57001),
            .I(N__56998));
    InMux I__11892 (
            .O(N__56998),
            .I(N__56995));
    LocalMux I__11891 (
            .O(N__56995),
            .I(N__56992));
    Odrv12 I__11890 (
            .O(N__56992),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7 ));
    InMux I__11889 (
            .O(N__56989),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15915 ));
    InMux I__11888 (
            .O(N__56986),
            .I(N__56983));
    LocalMux I__11887 (
            .O(N__56983),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4 ));
    CascadeMux I__11886 (
            .O(N__56980),
            .I(N__56977));
    InMux I__11885 (
            .O(N__56977),
            .I(N__56974));
    LocalMux I__11884 (
            .O(N__56974),
            .I(N__56971));
    Odrv4 I__11883 (
            .O(N__56971),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8 ));
    InMux I__11882 (
            .O(N__56968),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15916 ));
    InMux I__11881 (
            .O(N__56965),
            .I(N__56962));
    LocalMux I__11880 (
            .O(N__56962),
            .I(N__56959));
    Odrv12 I__11879 (
            .O(N__56959),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5 ));
    CascadeMux I__11878 (
            .O(N__56956),
            .I(N__56953));
    InMux I__11877 (
            .O(N__56953),
            .I(N__56950));
    LocalMux I__11876 (
            .O(N__56950),
            .I(N__56947));
    Odrv4 I__11875 (
            .O(N__56947),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9 ));
    InMux I__11874 (
            .O(N__56944),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15917 ));
    InMux I__11873 (
            .O(N__56941),
            .I(N__56938));
    LocalMux I__11872 (
            .O(N__56938),
            .I(N__56935));
    Odrv4 I__11871 (
            .O(N__56935),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6 ));
    CascadeMux I__11870 (
            .O(N__56932),
            .I(N__56929));
    InMux I__11869 (
            .O(N__56929),
            .I(N__56926));
    LocalMux I__11868 (
            .O(N__56926),
            .I(N__56923));
    Odrv4 I__11867 (
            .O(N__56923),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10 ));
    InMux I__11866 (
            .O(N__56920),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15918 ));
    InMux I__11865 (
            .O(N__56917),
            .I(N__56914));
    LocalMux I__11864 (
            .O(N__56914),
            .I(N__56910));
    InMux I__11863 (
            .O(N__56913),
            .I(N__56907));
    Span4Mux_v I__11862 (
            .O(N__56910),
            .I(N__56904));
    LocalMux I__11861 (
            .O(N__56907),
            .I(N__56901));
    Odrv4 I__11860 (
            .O(N__56904),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0 ));
    Odrv4 I__11859 (
            .O(N__56901),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0 ));
    CascadeMux I__11858 (
            .O(N__56896),
            .I(N__56893));
    InMux I__11857 (
            .O(N__56893),
            .I(N__56890));
    LocalMux I__11856 (
            .O(N__56890),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11 ));
    InMux I__11855 (
            .O(N__56887),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15919 ));
    InMux I__11854 (
            .O(N__56884),
            .I(N__56881));
    LocalMux I__11853 (
            .O(N__56881),
            .I(N__56878));
    Span4Mux_h I__11852 (
            .O(N__56878),
            .I(N__56875));
    Odrv4 I__11851 (
            .O(N__56875),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n400 ));
    InMux I__11850 (
            .O(N__56872),
            .I(bfn_21_22_0_));
    InMux I__11849 (
            .O(N__56869),
            .I(N__56866));
    LocalMux I__11848 (
            .O(N__56866),
            .I(N__56863));
    Span4Mux_h I__11847 (
            .O(N__56863),
            .I(N__56860));
    Odrv4 I__11846 (
            .O(N__56860),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n449 ));
    InMux I__11845 (
            .O(N__56857),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18182 ));
    InMux I__11844 (
            .O(N__56854),
            .I(N__56851));
    LocalMux I__11843 (
            .O(N__56851),
            .I(N__56848));
    Span12Mux_h I__11842 (
            .O(N__56848),
            .I(N__56845));
    Odrv12 I__11841 (
            .O(N__56845),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n498 ));
    InMux I__11840 (
            .O(N__56842),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18183 ));
    InMux I__11839 (
            .O(N__56839),
            .I(N__56836));
    LocalMux I__11838 (
            .O(N__56836),
            .I(N__56833));
    Span4Mux_h I__11837 (
            .O(N__56833),
            .I(N__56830));
    Odrv4 I__11836 (
            .O(N__56830),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n547 ));
    InMux I__11835 (
            .O(N__56827),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18184 ));
    InMux I__11834 (
            .O(N__56824),
            .I(N__56814));
    InMux I__11833 (
            .O(N__56823),
            .I(N__56794));
    InMux I__11832 (
            .O(N__56822),
            .I(N__56794));
    InMux I__11831 (
            .O(N__56821),
            .I(N__56794));
    InMux I__11830 (
            .O(N__56820),
            .I(N__56785));
    InMux I__11829 (
            .O(N__56819),
            .I(N__56785));
    InMux I__11828 (
            .O(N__56818),
            .I(N__56785));
    InMux I__11827 (
            .O(N__56817),
            .I(N__56785));
    LocalMux I__11826 (
            .O(N__56814),
            .I(N__56775));
    InMux I__11825 (
            .O(N__56813),
            .I(N__56766));
    InMux I__11824 (
            .O(N__56812),
            .I(N__56766));
    InMux I__11823 (
            .O(N__56811),
            .I(N__56766));
    InMux I__11822 (
            .O(N__56810),
            .I(N__56766));
    InMux I__11821 (
            .O(N__56809),
            .I(N__56757));
    InMux I__11820 (
            .O(N__56808),
            .I(N__56757));
    InMux I__11819 (
            .O(N__56807),
            .I(N__56757));
    InMux I__11818 (
            .O(N__56806),
            .I(N__56757));
    InMux I__11817 (
            .O(N__56805),
            .I(N__56752));
    InMux I__11816 (
            .O(N__56804),
            .I(N__56752));
    InMux I__11815 (
            .O(N__56803),
            .I(N__56745));
    InMux I__11814 (
            .O(N__56802),
            .I(N__56745));
    InMux I__11813 (
            .O(N__56801),
            .I(N__56745));
    LocalMux I__11812 (
            .O(N__56794),
            .I(N__56740));
    LocalMux I__11811 (
            .O(N__56785),
            .I(N__56740));
    InMux I__11810 (
            .O(N__56784),
            .I(N__56733));
    InMux I__11809 (
            .O(N__56783),
            .I(N__56733));
    InMux I__11808 (
            .O(N__56782),
            .I(N__56733));
    InMux I__11807 (
            .O(N__56781),
            .I(N__56724));
    InMux I__11806 (
            .O(N__56780),
            .I(N__56724));
    InMux I__11805 (
            .O(N__56779),
            .I(N__56724));
    InMux I__11804 (
            .O(N__56778),
            .I(N__56724));
    Odrv4 I__11803 (
            .O(N__56775),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11802 (
            .O(N__56766),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11801 (
            .O(N__56757),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11800 (
            .O(N__56752),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11799 (
            .O(N__56745),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    Odrv12 I__11798 (
            .O(N__56740),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11797 (
            .O(N__56733),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    LocalMux I__11796 (
            .O(N__56724),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ));
    InMux I__11795 (
            .O(N__56707),
            .I(N__56704));
    LocalMux I__11794 (
            .O(N__56704),
            .I(N__56701));
    Span4Mux_h I__11793 (
            .O(N__56701),
            .I(N__56698));
    Odrv4 I__11792 (
            .O(N__56698),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n596 ));
    InMux I__11791 (
            .O(N__56695),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18185 ));
    CascadeMux I__11790 (
            .O(N__56692),
            .I(N__56689));
    InMux I__11789 (
            .O(N__56689),
            .I(N__56686));
    LocalMux I__11788 (
            .O(N__56686),
            .I(N__56683));
    Span4Mux_v I__11787 (
            .O(N__56683),
            .I(N__56680));
    Odrv4 I__11786 (
            .O(N__56680),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n645 ));
    InMux I__11785 (
            .O(N__56677),
            .I(N__56671));
    InMux I__11784 (
            .O(N__56676),
            .I(N__56671));
    LocalMux I__11783 (
            .O(N__56671),
            .I(N__56668));
    Span4Mux_v I__11782 (
            .O(N__56668),
            .I(N__56665));
    Odrv4 I__11781 (
            .O(N__56665),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n691 ));
    InMux I__11780 (
            .O(N__56662),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18186 ));
    InMux I__11779 (
            .O(N__56659),
            .I(N__56656));
    LocalMux I__11778 (
            .O(N__56656),
            .I(N__56653));
    Span4Mux_v I__11777 (
            .O(N__56653),
            .I(N__56650));
    Odrv4 I__11776 (
            .O(N__56650),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n694 ));
    CascadeMux I__11775 (
            .O(N__56647),
            .I(N__56644));
    InMux I__11774 (
            .O(N__56644),
            .I(N__56641));
    LocalMux I__11773 (
            .O(N__56641),
            .I(N__56638));
    Span4Mux_v I__11772 (
            .O(N__56638),
            .I(N__56635));
    Odrv4 I__11771 (
            .O(N__56635),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n742 ));
    InMux I__11770 (
            .O(N__56632),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18187 ));
    InMux I__11769 (
            .O(N__56629),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743 ));
    CascadeMux I__11768 (
            .O(N__56626),
            .I(N__56623));
    InMux I__11767 (
            .O(N__56623),
            .I(N__56620));
    LocalMux I__11766 (
            .O(N__56620),
            .I(N__56617));
    Span4Mux_h I__11765 (
            .O(N__56617),
            .I(N__56614));
    Odrv4 I__11764 (
            .O(N__56614),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO ));
    CascadeMux I__11763 (
            .O(N__56611),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_ ));
    InMux I__11762 (
            .O(N__56608),
            .I(N__56605));
    LocalMux I__11761 (
            .O(N__56605),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19308 ));
    InMux I__11760 (
            .O(N__56602),
            .I(N__56599));
    LocalMux I__11759 (
            .O(N__56599),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n57 ));
    InMux I__11758 (
            .O(N__56596),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18174 ));
    CascadeMux I__11757 (
            .O(N__56593),
            .I(N__56590));
    InMux I__11756 (
            .O(N__56590),
            .I(N__56587));
    LocalMux I__11755 (
            .O(N__56587),
            .I(N__56584));
    Span4Mux_v I__11754 (
            .O(N__56584),
            .I(N__56581));
    Span4Mux_v I__11753 (
            .O(N__56581),
            .I(N__56578));
    Odrv4 I__11752 (
            .O(N__56578),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n106 ));
    InMux I__11751 (
            .O(N__56575),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18175 ));
    InMux I__11750 (
            .O(N__56572),
            .I(N__56569));
    LocalMux I__11749 (
            .O(N__56569),
            .I(N__56566));
    Span4Mux_h I__11748 (
            .O(N__56566),
            .I(N__56563));
    Odrv4 I__11747 (
            .O(N__56563),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n155 ));
    InMux I__11746 (
            .O(N__56560),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18176 ));
    InMux I__11745 (
            .O(N__56557),
            .I(N__56554));
    LocalMux I__11744 (
            .O(N__56554),
            .I(N__56551));
    Span4Mux_v I__11743 (
            .O(N__56551),
            .I(N__56548));
    Odrv4 I__11742 (
            .O(N__56548),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n204 ));
    InMux I__11741 (
            .O(N__56545),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18177 ));
    InMux I__11740 (
            .O(N__56542),
            .I(N__56539));
    LocalMux I__11739 (
            .O(N__56539),
            .I(N__56536));
    Span4Mux_v I__11738 (
            .O(N__56536),
            .I(N__56533));
    Odrv4 I__11737 (
            .O(N__56533),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n253 ));
    InMux I__11736 (
            .O(N__56530),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18178 ));
    InMux I__11735 (
            .O(N__56527),
            .I(N__56524));
    LocalMux I__11734 (
            .O(N__56524),
            .I(N__56521));
    Span4Mux_v I__11733 (
            .O(N__56521),
            .I(N__56518));
    Sp12to4 I__11732 (
            .O(N__56518),
            .I(N__56515));
    Odrv12 I__11731 (
            .O(N__56515),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n302 ));
    InMux I__11730 (
            .O(N__56512),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18179 ));
    InMux I__11729 (
            .O(N__56509),
            .I(N__56506));
    LocalMux I__11728 (
            .O(N__56506),
            .I(N__56503));
    Span4Mux_h I__11727 (
            .O(N__56503),
            .I(N__56500));
    Odrv4 I__11726 (
            .O(N__56500),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n351 ));
    InMux I__11725 (
            .O(N__56497),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18180 ));
    InMux I__11724 (
            .O(N__56494),
            .I(N__56485));
    InMux I__11723 (
            .O(N__56493),
            .I(N__56485));
    InMux I__11722 (
            .O(N__56492),
            .I(N__56485));
    LocalMux I__11721 (
            .O(N__56485),
            .I(N__56473));
    InMux I__11720 (
            .O(N__56484),
            .I(N__56464));
    InMux I__11719 (
            .O(N__56483),
            .I(N__56464));
    InMux I__11718 (
            .O(N__56482),
            .I(N__56464));
    InMux I__11717 (
            .O(N__56481),
            .I(N__56464));
    CascadeMux I__11716 (
            .O(N__56480),
            .I(N__56451));
    CascadeMux I__11715 (
            .O(N__56479),
            .I(N__56444));
    InMux I__11714 (
            .O(N__56478),
            .I(N__56433));
    InMux I__11713 (
            .O(N__56477),
            .I(N__56433));
    InMux I__11712 (
            .O(N__56476),
            .I(N__56433));
    Span4Mux_v I__11711 (
            .O(N__56473),
            .I(N__56428));
    LocalMux I__11710 (
            .O(N__56464),
            .I(N__56428));
    InMux I__11709 (
            .O(N__56463),
            .I(N__56425));
    InMux I__11708 (
            .O(N__56462),
            .I(N__56412));
    InMux I__11707 (
            .O(N__56461),
            .I(N__56412));
    InMux I__11706 (
            .O(N__56460),
            .I(N__56412));
    InMux I__11705 (
            .O(N__56459),
            .I(N__56412));
    InMux I__11704 (
            .O(N__56458),
            .I(N__56412));
    InMux I__11703 (
            .O(N__56457),
            .I(N__56412));
    InMux I__11702 (
            .O(N__56456),
            .I(N__56399));
    InMux I__11701 (
            .O(N__56455),
            .I(N__56399));
    InMux I__11700 (
            .O(N__56454),
            .I(N__56399));
    InMux I__11699 (
            .O(N__56451),
            .I(N__56399));
    InMux I__11698 (
            .O(N__56450),
            .I(N__56399));
    InMux I__11697 (
            .O(N__56449),
            .I(N__56399));
    InMux I__11696 (
            .O(N__56448),
            .I(N__56390));
    InMux I__11695 (
            .O(N__56447),
            .I(N__56390));
    InMux I__11694 (
            .O(N__56444),
            .I(N__56390));
    InMux I__11693 (
            .O(N__56443),
            .I(N__56390));
    InMux I__11692 (
            .O(N__56442),
            .I(N__56383));
    InMux I__11691 (
            .O(N__56441),
            .I(N__56383));
    InMux I__11690 (
            .O(N__56440),
            .I(N__56383));
    LocalMux I__11689 (
            .O(N__56433),
            .I(Saturate_out1_31__N_266_adj_2417));
    Odrv4 I__11688 (
            .O(N__56428),
            .I(Saturate_out1_31__N_266_adj_2417));
    LocalMux I__11687 (
            .O(N__56425),
            .I(Saturate_out1_31__N_266_adj_2417));
    LocalMux I__11686 (
            .O(N__56412),
            .I(Saturate_out1_31__N_266_adj_2417));
    LocalMux I__11685 (
            .O(N__56399),
            .I(Saturate_out1_31__N_266_adj_2417));
    LocalMux I__11684 (
            .O(N__56390),
            .I(Saturate_out1_31__N_266_adj_2417));
    LocalMux I__11683 (
            .O(N__56383),
            .I(Saturate_out1_31__N_266_adj_2417));
    InMux I__11682 (
            .O(N__56368),
            .I(N__56353));
    InMux I__11681 (
            .O(N__56367),
            .I(N__56353));
    InMux I__11680 (
            .O(N__56366),
            .I(N__56353));
    CascadeMux I__11679 (
            .O(N__56365),
            .I(N__56349));
    CascadeMux I__11678 (
            .O(N__56364),
            .I(N__56346));
    InMux I__11677 (
            .O(N__56363),
            .I(N__56335));
    InMux I__11676 (
            .O(N__56362),
            .I(N__56335));
    InMux I__11675 (
            .O(N__56361),
            .I(N__56335));
    CascadeMux I__11674 (
            .O(N__56360),
            .I(N__56332));
    LocalMux I__11673 (
            .O(N__56353),
            .I(N__56326));
    InMux I__11672 (
            .O(N__56352),
            .I(N__56313));
    InMux I__11671 (
            .O(N__56349),
            .I(N__56313));
    InMux I__11670 (
            .O(N__56346),
            .I(N__56313));
    InMux I__11669 (
            .O(N__56345),
            .I(N__56313));
    InMux I__11668 (
            .O(N__56344),
            .I(N__56313));
    InMux I__11667 (
            .O(N__56343),
            .I(N__56313));
    InMux I__11666 (
            .O(N__56342),
            .I(N__56310));
    LocalMux I__11665 (
            .O(N__56335),
            .I(N__56294));
    InMux I__11664 (
            .O(N__56332),
            .I(N__56285));
    InMux I__11663 (
            .O(N__56331),
            .I(N__56285));
    InMux I__11662 (
            .O(N__56330),
            .I(N__56285));
    InMux I__11661 (
            .O(N__56329),
            .I(N__56285));
    Span4Mux_v I__11660 (
            .O(N__56326),
            .I(N__56278));
    LocalMux I__11659 (
            .O(N__56313),
            .I(N__56278));
    LocalMux I__11658 (
            .O(N__56310),
            .I(N__56278));
    InMux I__11657 (
            .O(N__56309),
            .I(N__56269));
    InMux I__11656 (
            .O(N__56308),
            .I(N__56269));
    InMux I__11655 (
            .O(N__56307),
            .I(N__56269));
    InMux I__11654 (
            .O(N__56306),
            .I(N__56269));
    InMux I__11653 (
            .O(N__56305),
            .I(N__56260));
    InMux I__11652 (
            .O(N__56304),
            .I(N__56260));
    InMux I__11651 (
            .O(N__56303),
            .I(N__56260));
    InMux I__11650 (
            .O(N__56302),
            .I(N__56260));
    InMux I__11649 (
            .O(N__56301),
            .I(N__56251));
    InMux I__11648 (
            .O(N__56300),
            .I(N__56251));
    InMux I__11647 (
            .O(N__56299),
            .I(N__56251));
    InMux I__11646 (
            .O(N__56298),
            .I(N__56251));
    InMux I__11645 (
            .O(N__56297),
            .I(N__56248));
    Odrv4 I__11644 (
            .O(N__56294),
            .I(Saturate_out1_31__N_267_adj_2418));
    LocalMux I__11643 (
            .O(N__56285),
            .I(Saturate_out1_31__N_267_adj_2418));
    Odrv4 I__11642 (
            .O(N__56278),
            .I(Saturate_out1_31__N_267_adj_2418));
    LocalMux I__11641 (
            .O(N__56269),
            .I(Saturate_out1_31__N_267_adj_2418));
    LocalMux I__11640 (
            .O(N__56260),
            .I(Saturate_out1_31__N_267_adj_2418));
    LocalMux I__11639 (
            .O(N__56251),
            .I(Saturate_out1_31__N_267_adj_2418));
    LocalMux I__11638 (
            .O(N__56248),
            .I(Saturate_out1_31__N_267_adj_2418));
    CascadeMux I__11637 (
            .O(N__56233),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_ ));
    CascadeMux I__11636 (
            .O(N__56230),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_ ));
    InMux I__11635 (
            .O(N__56227),
            .I(N__56224));
    LocalMux I__11634 (
            .O(N__56224),
            .I(N__56221));
    Span4Mux_v I__11633 (
            .O(N__56221),
            .I(N__56218));
    Odrv4 I__11632 (
            .O(N__56218),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492 ));
    CascadeMux I__11631 (
            .O(N__56215),
            .I(N__56211));
    CascadeMux I__11630 (
            .O(N__56214),
            .I(N__56208));
    InMux I__11629 (
            .O(N__56211),
            .I(N__56201));
    InMux I__11628 (
            .O(N__56208),
            .I(N__56198));
    CascadeMux I__11627 (
            .O(N__56207),
            .I(N__56194));
    CascadeMux I__11626 (
            .O(N__56206),
            .I(N__56191));
    CascadeMux I__11625 (
            .O(N__56205),
            .I(N__56186));
    CascadeMux I__11624 (
            .O(N__56204),
            .I(N__56183));
    LocalMux I__11623 (
            .O(N__56201),
            .I(N__56179));
    LocalMux I__11622 (
            .O(N__56198),
            .I(N__56176));
    CascadeMux I__11621 (
            .O(N__56197),
            .I(N__56173));
    InMux I__11620 (
            .O(N__56194),
            .I(N__56170));
    InMux I__11619 (
            .O(N__56191),
            .I(N__56167));
    CascadeMux I__11618 (
            .O(N__56190),
            .I(N__56164));
    CascadeMux I__11617 (
            .O(N__56189),
            .I(N__56161));
    InMux I__11616 (
            .O(N__56186),
            .I(N__56157));
    InMux I__11615 (
            .O(N__56183),
            .I(N__56154));
    CascadeMux I__11614 (
            .O(N__56182),
            .I(N__56151));
    Span4Mux_v I__11613 (
            .O(N__56179),
            .I(N__56142));
    Span4Mux_h I__11612 (
            .O(N__56176),
            .I(N__56139));
    InMux I__11611 (
            .O(N__56173),
            .I(N__56136));
    LocalMux I__11610 (
            .O(N__56170),
            .I(N__56131));
    LocalMux I__11609 (
            .O(N__56167),
            .I(N__56131));
    InMux I__11608 (
            .O(N__56164),
            .I(N__56128));
    InMux I__11607 (
            .O(N__56161),
            .I(N__56125));
    CascadeMux I__11606 (
            .O(N__56160),
            .I(N__56122));
    LocalMux I__11605 (
            .O(N__56157),
            .I(N__56116));
    LocalMux I__11604 (
            .O(N__56154),
            .I(N__56116));
    InMux I__11603 (
            .O(N__56151),
            .I(N__56113));
    CascadeMux I__11602 (
            .O(N__56150),
            .I(N__56110));
    CascadeMux I__11601 (
            .O(N__56149),
            .I(N__56107));
    CascadeMux I__11600 (
            .O(N__56148),
            .I(N__56103));
    CascadeMux I__11599 (
            .O(N__56147),
            .I(N__56099));
    CascadeMux I__11598 (
            .O(N__56146),
            .I(N__56095));
    CascadeMux I__11597 (
            .O(N__56145),
            .I(N__56091));
    Span4Mux_v I__11596 (
            .O(N__56142),
            .I(N__56083));
    Span4Mux_v I__11595 (
            .O(N__56139),
            .I(N__56083));
    LocalMux I__11594 (
            .O(N__56136),
            .I(N__56083));
    Span4Mux_v I__11593 (
            .O(N__56131),
            .I(N__56076));
    LocalMux I__11592 (
            .O(N__56128),
            .I(N__56076));
    LocalMux I__11591 (
            .O(N__56125),
            .I(N__56076));
    InMux I__11590 (
            .O(N__56122),
            .I(N__56073));
    InMux I__11589 (
            .O(N__56121),
            .I(N__56070));
    Span4Mux_v I__11588 (
            .O(N__56116),
            .I(N__56065));
    LocalMux I__11587 (
            .O(N__56113),
            .I(N__56065));
    InMux I__11586 (
            .O(N__56110),
            .I(N__56062));
    InMux I__11585 (
            .O(N__56107),
            .I(N__56059));
    InMux I__11584 (
            .O(N__56106),
            .I(N__56042));
    InMux I__11583 (
            .O(N__56103),
            .I(N__56042));
    InMux I__11582 (
            .O(N__56102),
            .I(N__56042));
    InMux I__11581 (
            .O(N__56099),
            .I(N__56042));
    InMux I__11580 (
            .O(N__56098),
            .I(N__56042));
    InMux I__11579 (
            .O(N__56095),
            .I(N__56042));
    InMux I__11578 (
            .O(N__56094),
            .I(N__56042));
    InMux I__11577 (
            .O(N__56091),
            .I(N__56042));
    CascadeMux I__11576 (
            .O(N__56090),
            .I(N__56039));
    Span4Mux_h I__11575 (
            .O(N__56083),
            .I(N__56035));
    Span4Mux_v I__11574 (
            .O(N__56076),
            .I(N__56030));
    LocalMux I__11573 (
            .O(N__56073),
            .I(N__56030));
    LocalMux I__11572 (
            .O(N__56070),
            .I(N__56027));
    Span4Mux_v I__11571 (
            .O(N__56065),
            .I(N__56020));
    LocalMux I__11570 (
            .O(N__56062),
            .I(N__56020));
    LocalMux I__11569 (
            .O(N__56059),
            .I(N__56020));
    LocalMux I__11568 (
            .O(N__56042),
            .I(N__56017));
    InMux I__11567 (
            .O(N__56039),
            .I(N__56014));
    CascadeMux I__11566 (
            .O(N__56038),
            .I(N__56010));
    Span4Mux_v I__11565 (
            .O(N__56035),
            .I(N__56007));
    Span4Mux_v I__11564 (
            .O(N__56030),
            .I(N__56004));
    Span4Mux_h I__11563 (
            .O(N__56027),
            .I(N__55995));
    Span4Mux_v I__11562 (
            .O(N__56020),
            .I(N__55995));
    Span4Mux_v I__11561 (
            .O(N__56017),
            .I(N__55995));
    LocalMux I__11560 (
            .O(N__56014),
            .I(N__55995));
    InMux I__11559 (
            .O(N__56013),
            .I(N__55990));
    InMux I__11558 (
            .O(N__56010),
            .I(N__55990));
    Odrv4 I__11557 (
            .O(N__56007),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n129 ));
    Odrv4 I__11556 (
            .O(N__56004),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n129 ));
    Odrv4 I__11555 (
            .O(N__55995),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n129 ));
    LocalMux I__11554 (
            .O(N__55990),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n129 ));
    InMux I__11553 (
            .O(N__55981),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17744 ));
    InMux I__11552 (
            .O(N__55978),
            .I(N__55975));
    LocalMux I__11551 (
            .O(N__55975),
            .I(N__55972));
    Span4Mux_v I__11550 (
            .O(N__55972),
            .I(N__55969));
    Odrv4 I__11549 (
            .O(N__55969),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469 ));
    CascadeMux I__11548 (
            .O(N__55966),
            .I(N__55961));
    CascadeMux I__11547 (
            .O(N__55965),
            .I(N__55957));
    CascadeMux I__11546 (
            .O(N__55964),
            .I(N__55953));
    InMux I__11545 (
            .O(N__55961),
            .I(N__55950));
    InMux I__11544 (
            .O(N__55960),
            .I(N__55947));
    InMux I__11543 (
            .O(N__55957),
            .I(N__55941));
    CascadeMux I__11542 (
            .O(N__55956),
            .I(N__55936));
    InMux I__11541 (
            .O(N__55953),
            .I(N__55933));
    LocalMux I__11540 (
            .O(N__55950),
            .I(N__55928));
    LocalMux I__11539 (
            .O(N__55947),
            .I(N__55928));
    CascadeMux I__11538 (
            .O(N__55946),
            .I(N__55925));
    CascadeMux I__11537 (
            .O(N__55945),
            .I(N__55922));
    CascadeMux I__11536 (
            .O(N__55944),
            .I(N__55919));
    LocalMux I__11535 (
            .O(N__55941),
            .I(N__55912));
    CascadeMux I__11534 (
            .O(N__55940),
            .I(N__55909));
    CascadeMux I__11533 (
            .O(N__55939),
            .I(N__55906));
    InMux I__11532 (
            .O(N__55936),
            .I(N__55903));
    LocalMux I__11531 (
            .O(N__55933),
            .I(N__55900));
    Span4Mux_v I__11530 (
            .O(N__55928),
            .I(N__55897));
    InMux I__11529 (
            .O(N__55925),
            .I(N__55894));
    InMux I__11528 (
            .O(N__55922),
            .I(N__55891));
    InMux I__11527 (
            .O(N__55919),
            .I(N__55888));
    CascadeMux I__11526 (
            .O(N__55918),
            .I(N__55885));
    CascadeMux I__11525 (
            .O(N__55917),
            .I(N__55882));
    CascadeMux I__11524 (
            .O(N__55916),
            .I(N__55879));
    CascadeMux I__11523 (
            .O(N__55915),
            .I(N__55876));
    Span4Mux_v I__11522 (
            .O(N__55912),
            .I(N__55869));
    InMux I__11521 (
            .O(N__55909),
            .I(N__55866));
    InMux I__11520 (
            .O(N__55906),
            .I(N__55863));
    LocalMux I__11519 (
            .O(N__55903),
            .I(N__55860));
    Span4Mux_h I__11518 (
            .O(N__55900),
            .I(N__55849));
    Span4Mux_h I__11517 (
            .O(N__55897),
            .I(N__55849));
    LocalMux I__11516 (
            .O(N__55894),
            .I(N__55849));
    LocalMux I__11515 (
            .O(N__55891),
            .I(N__55849));
    LocalMux I__11514 (
            .O(N__55888),
            .I(N__55849));
    InMux I__11513 (
            .O(N__55885),
            .I(N__55846));
    InMux I__11512 (
            .O(N__55882),
            .I(N__55843));
    InMux I__11511 (
            .O(N__55879),
            .I(N__55840));
    InMux I__11510 (
            .O(N__55876),
            .I(N__55836));
    CascadeMux I__11509 (
            .O(N__55875),
            .I(N__55832));
    CascadeMux I__11508 (
            .O(N__55874),
            .I(N__55828));
    CascadeMux I__11507 (
            .O(N__55873),
            .I(N__55824));
    CascadeMux I__11506 (
            .O(N__55872),
            .I(N__55820));
    Sp12to4 I__11505 (
            .O(N__55869),
            .I(N__55813));
    LocalMux I__11504 (
            .O(N__55866),
            .I(N__55813));
    LocalMux I__11503 (
            .O(N__55863),
            .I(N__55813));
    Span4Mux_h I__11502 (
            .O(N__55860),
            .I(N__55806));
    Span4Mux_v I__11501 (
            .O(N__55849),
            .I(N__55806));
    LocalMux I__11500 (
            .O(N__55846),
            .I(N__55806));
    LocalMux I__11499 (
            .O(N__55843),
            .I(N__55803));
    LocalMux I__11498 (
            .O(N__55840),
            .I(N__55800));
    InMux I__11497 (
            .O(N__55839),
            .I(N__55797));
    LocalMux I__11496 (
            .O(N__55836),
            .I(N__55794));
    InMux I__11495 (
            .O(N__55835),
            .I(N__55777));
    InMux I__11494 (
            .O(N__55832),
            .I(N__55777));
    InMux I__11493 (
            .O(N__55831),
            .I(N__55777));
    InMux I__11492 (
            .O(N__55828),
            .I(N__55777));
    InMux I__11491 (
            .O(N__55827),
            .I(N__55777));
    InMux I__11490 (
            .O(N__55824),
            .I(N__55777));
    InMux I__11489 (
            .O(N__55823),
            .I(N__55777));
    InMux I__11488 (
            .O(N__55820),
            .I(N__55777));
    Span12Mux_h I__11487 (
            .O(N__55813),
            .I(N__55774));
    Span4Mux_v I__11486 (
            .O(N__55806),
            .I(N__55769));
    Span4Mux_h I__11485 (
            .O(N__55803),
            .I(N__55769));
    Span4Mux_v I__11484 (
            .O(N__55800),
            .I(N__55760));
    LocalMux I__11483 (
            .O(N__55797),
            .I(N__55760));
    Span4Mux_v I__11482 (
            .O(N__55794),
            .I(N__55760));
    LocalMux I__11481 (
            .O(N__55777),
            .I(N__55760));
    Odrv12 I__11480 (
            .O(N__55774),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n132 ));
    Odrv4 I__11479 (
            .O(N__55769),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n132 ));
    Odrv4 I__11478 (
            .O(N__55760),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n132 ));
    InMux I__11477 (
            .O(N__55753),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17745 ));
    InMux I__11476 (
            .O(N__55750),
            .I(N__55747));
    LocalMux I__11475 (
            .O(N__55747),
            .I(N__55744));
    Span4Mux_v I__11474 (
            .O(N__55744),
            .I(N__55741));
    Odrv4 I__11473 (
            .O(N__55741),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454 ));
    CascadeMux I__11472 (
            .O(N__55738),
            .I(N__55733));
    CascadeMux I__11471 (
            .O(N__55737),
            .I(N__55730));
    CascadeMux I__11470 (
            .O(N__55736),
            .I(N__55726));
    InMux I__11469 (
            .O(N__55733),
            .I(N__55719));
    InMux I__11468 (
            .O(N__55730),
            .I(N__55714));
    CascadeMux I__11467 (
            .O(N__55729),
            .I(N__55711));
    InMux I__11466 (
            .O(N__55726),
            .I(N__55708));
    CascadeMux I__11465 (
            .O(N__55725),
            .I(N__55705));
    CascadeMux I__11464 (
            .O(N__55724),
            .I(N__55702));
    CascadeMux I__11463 (
            .O(N__55723),
            .I(N__55699));
    CascadeMux I__11462 (
            .O(N__55722),
            .I(N__55694));
    LocalMux I__11461 (
            .O(N__55719),
            .I(N__55691));
    CascadeMux I__11460 (
            .O(N__55718),
            .I(N__55688));
    CascadeMux I__11459 (
            .O(N__55717),
            .I(N__55685));
    LocalMux I__11458 (
            .O(N__55714),
            .I(N__55682));
    InMux I__11457 (
            .O(N__55711),
            .I(N__55679));
    LocalMux I__11456 (
            .O(N__55708),
            .I(N__55676));
    InMux I__11455 (
            .O(N__55705),
            .I(N__55673));
    InMux I__11454 (
            .O(N__55702),
            .I(N__55670));
    InMux I__11453 (
            .O(N__55699),
            .I(N__55667));
    CascadeMux I__11452 (
            .O(N__55698),
            .I(N__55664));
    CascadeMux I__11451 (
            .O(N__55697),
            .I(N__55660));
    InMux I__11450 (
            .O(N__55694),
            .I(N__55656));
    Span4Mux_v I__11449 (
            .O(N__55691),
            .I(N__55653));
    InMux I__11448 (
            .O(N__55688),
            .I(N__55650));
    InMux I__11447 (
            .O(N__55685),
            .I(N__55647));
    Span4Mux_v I__11446 (
            .O(N__55682),
            .I(N__55642));
    LocalMux I__11445 (
            .O(N__55679),
            .I(N__55642));
    Span4Mux_v I__11444 (
            .O(N__55676),
            .I(N__55633));
    LocalMux I__11443 (
            .O(N__55673),
            .I(N__55633));
    LocalMux I__11442 (
            .O(N__55670),
            .I(N__55633));
    LocalMux I__11441 (
            .O(N__55667),
            .I(N__55633));
    InMux I__11440 (
            .O(N__55664),
            .I(N__55630));
    InMux I__11439 (
            .O(N__55663),
            .I(N__55627));
    InMux I__11438 (
            .O(N__55660),
            .I(N__55624));
    CascadeMux I__11437 (
            .O(N__55659),
            .I(N__55621));
    LocalMux I__11436 (
            .O(N__55656),
            .I(N__55612));
    Span4Mux_v I__11435 (
            .O(N__55653),
            .I(N__55605));
    LocalMux I__11434 (
            .O(N__55650),
            .I(N__55605));
    LocalMux I__11433 (
            .O(N__55647),
            .I(N__55605));
    Span4Mux_h I__11432 (
            .O(N__55642),
            .I(N__55598));
    Span4Mux_v I__11431 (
            .O(N__55633),
            .I(N__55598));
    LocalMux I__11430 (
            .O(N__55630),
            .I(N__55598));
    LocalMux I__11429 (
            .O(N__55627),
            .I(N__55595));
    LocalMux I__11428 (
            .O(N__55624),
            .I(N__55592));
    InMux I__11427 (
            .O(N__55621),
            .I(N__55589));
    CascadeMux I__11426 (
            .O(N__55620),
            .I(N__55586));
    CascadeMux I__11425 (
            .O(N__55619),
            .I(N__55583));
    CascadeMux I__11424 (
            .O(N__55618),
            .I(N__55579));
    CascadeMux I__11423 (
            .O(N__55617),
            .I(N__55576));
    CascadeMux I__11422 (
            .O(N__55616),
            .I(N__55573));
    CascadeMux I__11421 (
            .O(N__55615),
            .I(N__55570));
    Span12Mux_h I__11420 (
            .O(N__55612),
            .I(N__55567));
    Span4Mux_h I__11419 (
            .O(N__55605),
            .I(N__55564));
    Span4Mux_v I__11418 (
            .O(N__55598),
            .I(N__55557));
    Span4Mux_v I__11417 (
            .O(N__55595),
            .I(N__55557));
    Span4Mux_h I__11416 (
            .O(N__55592),
            .I(N__55557));
    LocalMux I__11415 (
            .O(N__55589),
            .I(N__55554));
    InMux I__11414 (
            .O(N__55586),
            .I(N__55549));
    InMux I__11413 (
            .O(N__55583),
            .I(N__55549));
    InMux I__11412 (
            .O(N__55582),
            .I(N__55540));
    InMux I__11411 (
            .O(N__55579),
            .I(N__55540));
    InMux I__11410 (
            .O(N__55576),
            .I(N__55540));
    InMux I__11409 (
            .O(N__55573),
            .I(N__55540));
    InMux I__11408 (
            .O(N__55570),
            .I(N__55537));
    Odrv12 I__11407 (
            .O(N__55567),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    Odrv4 I__11406 (
            .O(N__55564),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    Odrv4 I__11405 (
            .O(N__55557),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    Odrv4 I__11404 (
            .O(N__55554),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    LocalMux I__11403 (
            .O(N__55549),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    LocalMux I__11402 (
            .O(N__55540),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    LocalMux I__11401 (
            .O(N__55537),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ));
    InMux I__11400 (
            .O(N__55522),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17746 ));
    CascadeMux I__11399 (
            .O(N__55519),
            .I(N__55516));
    InMux I__11398 (
            .O(N__55516),
            .I(N__55513));
    LocalMux I__11397 (
            .O(N__55513),
            .I(N__55506));
    InMux I__11396 (
            .O(N__55512),
            .I(N__55497));
    InMux I__11395 (
            .O(N__55511),
            .I(N__55497));
    InMux I__11394 (
            .O(N__55510),
            .I(N__55497));
    InMux I__11393 (
            .O(N__55509),
            .I(N__55497));
    Span4Mux_v I__11392 (
            .O(N__55506),
            .I(N__55481));
    LocalMux I__11391 (
            .O(N__55497),
            .I(N__55481));
    InMux I__11390 (
            .O(N__55496),
            .I(N__55472));
    InMux I__11389 (
            .O(N__55495),
            .I(N__55472));
    InMux I__11388 (
            .O(N__55494),
            .I(N__55472));
    InMux I__11387 (
            .O(N__55493),
            .I(N__55472));
    InMux I__11386 (
            .O(N__55492),
            .I(N__55465));
    InMux I__11385 (
            .O(N__55491),
            .I(N__55465));
    InMux I__11384 (
            .O(N__55490),
            .I(N__55465));
    InMux I__11383 (
            .O(N__55489),
            .I(N__55456));
    InMux I__11382 (
            .O(N__55488),
            .I(N__55456));
    InMux I__11381 (
            .O(N__55487),
            .I(N__55456));
    InMux I__11380 (
            .O(N__55486),
            .I(N__55456));
    Span4Mux_h I__11379 (
            .O(N__55481),
            .I(N__55435));
    LocalMux I__11378 (
            .O(N__55472),
            .I(N__55435));
    LocalMux I__11377 (
            .O(N__55465),
            .I(N__55435));
    LocalMux I__11376 (
            .O(N__55456),
            .I(N__55435));
    InMux I__11375 (
            .O(N__55455),
            .I(N__55430));
    InMux I__11374 (
            .O(N__55454),
            .I(N__55430));
    InMux I__11373 (
            .O(N__55453),
            .I(N__55423));
    InMux I__11372 (
            .O(N__55452),
            .I(N__55423));
    InMux I__11371 (
            .O(N__55451),
            .I(N__55423));
    InMux I__11370 (
            .O(N__55450),
            .I(N__55416));
    InMux I__11369 (
            .O(N__55449),
            .I(N__55416));
    InMux I__11368 (
            .O(N__55448),
            .I(N__55416));
    InMux I__11367 (
            .O(N__55447),
            .I(N__55407));
    InMux I__11366 (
            .O(N__55446),
            .I(N__55407));
    InMux I__11365 (
            .O(N__55445),
            .I(N__55407));
    InMux I__11364 (
            .O(N__55444),
            .I(N__55407));
    Span4Mux_v I__11363 (
            .O(N__55435),
            .I(N__55404));
    LocalMux I__11362 (
            .O(N__55430),
            .I(N__55395));
    LocalMux I__11361 (
            .O(N__55423),
            .I(N__55395));
    LocalMux I__11360 (
            .O(N__55416),
            .I(N__55395));
    LocalMux I__11359 (
            .O(N__55407),
            .I(N__55395));
    Odrv4 I__11358 (
            .O(N__55404),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201 ));
    Odrv12 I__11357 (
            .O(N__55395),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201 ));
    InMux I__11356 (
            .O(N__55390),
            .I(N__55387));
    LocalMux I__11355 (
            .O(N__55387),
            .I(N__55384));
    Span4Mux_v I__11354 (
            .O(N__55384),
            .I(N__55381));
    Odrv4 I__11353 (
            .O(N__55381),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434 ));
    CascadeMux I__11352 (
            .O(N__55378),
            .I(N__55374));
    CascadeMux I__11351 (
            .O(N__55377),
            .I(N__55371));
    InMux I__11350 (
            .O(N__55374),
            .I(N__55367));
    InMux I__11349 (
            .O(N__55371),
            .I(N__55360));
    InMux I__11348 (
            .O(N__55370),
            .I(N__55357));
    LocalMux I__11347 (
            .O(N__55367),
            .I(N__55353));
    CascadeMux I__11346 (
            .O(N__55366),
            .I(N__55350));
    CascadeMux I__11345 (
            .O(N__55365),
            .I(N__55345));
    CascadeMux I__11344 (
            .O(N__55364),
            .I(N__55342));
    CascadeMux I__11343 (
            .O(N__55363),
            .I(N__55338));
    LocalMux I__11342 (
            .O(N__55360),
            .I(N__55334));
    LocalMux I__11341 (
            .O(N__55357),
            .I(N__55331));
    CascadeMux I__11340 (
            .O(N__55356),
            .I(N__55328));
    Span4Mux_v I__11339 (
            .O(N__55353),
            .I(N__55325));
    InMux I__11338 (
            .O(N__55350),
            .I(N__55322));
    CascadeMux I__11337 (
            .O(N__55349),
            .I(N__55319));
    CascadeMux I__11336 (
            .O(N__55348),
            .I(N__55316));
    InMux I__11335 (
            .O(N__55345),
            .I(N__55313));
    InMux I__11334 (
            .O(N__55342),
            .I(N__55310));
    CascadeMux I__11333 (
            .O(N__55341),
            .I(N__55307));
    InMux I__11332 (
            .O(N__55338),
            .I(N__55303));
    CascadeMux I__11331 (
            .O(N__55337),
            .I(N__55300));
    Span4Mux_v I__11330 (
            .O(N__55334),
            .I(N__55297));
    Span4Mux_h I__11329 (
            .O(N__55331),
            .I(N__55294));
    InMux I__11328 (
            .O(N__55328),
            .I(N__55291));
    Span4Mux_h I__11327 (
            .O(N__55325),
            .I(N__55286));
    LocalMux I__11326 (
            .O(N__55322),
            .I(N__55286));
    InMux I__11325 (
            .O(N__55319),
            .I(N__55283));
    InMux I__11324 (
            .O(N__55316),
            .I(N__55280));
    LocalMux I__11323 (
            .O(N__55313),
            .I(N__55275));
    LocalMux I__11322 (
            .O(N__55310),
            .I(N__55275));
    InMux I__11321 (
            .O(N__55307),
            .I(N__55272));
    CascadeMux I__11320 (
            .O(N__55306),
            .I(N__55269));
    LocalMux I__11319 (
            .O(N__55303),
            .I(N__55263));
    InMux I__11318 (
            .O(N__55300),
            .I(N__55260));
    Span4Mux_v I__11317 (
            .O(N__55297),
            .I(N__55253));
    Span4Mux_v I__11316 (
            .O(N__55294),
            .I(N__55253));
    LocalMux I__11315 (
            .O(N__55291),
            .I(N__55253));
    Span4Mux_h I__11314 (
            .O(N__55286),
            .I(N__55242));
    LocalMux I__11313 (
            .O(N__55283),
            .I(N__55242));
    LocalMux I__11312 (
            .O(N__55280),
            .I(N__55242));
    Span4Mux_h I__11311 (
            .O(N__55275),
            .I(N__55242));
    LocalMux I__11310 (
            .O(N__55272),
            .I(N__55242));
    InMux I__11309 (
            .O(N__55269),
            .I(N__55239));
    InMux I__11308 (
            .O(N__55268),
            .I(N__55234));
    InMux I__11307 (
            .O(N__55267),
            .I(N__55234));
    CascadeMux I__11306 (
            .O(N__55266),
            .I(N__55230));
    Span12Mux_h I__11305 (
            .O(N__55263),
            .I(N__55224));
    LocalMux I__11304 (
            .O(N__55260),
            .I(N__55224));
    Span4Mux_h I__11303 (
            .O(N__55253),
            .I(N__55221));
    Span4Mux_v I__11302 (
            .O(N__55242),
            .I(N__55216));
    LocalMux I__11301 (
            .O(N__55239),
            .I(N__55216));
    LocalMux I__11300 (
            .O(N__55234),
            .I(N__55213));
    InMux I__11299 (
            .O(N__55233),
            .I(N__55210));
    InMux I__11298 (
            .O(N__55230),
            .I(N__55207));
    InMux I__11297 (
            .O(N__55229),
            .I(N__55204));
    Odrv12 I__11296 (
            .O(N__55224),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    Odrv4 I__11295 (
            .O(N__55221),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    Odrv4 I__11294 (
            .O(N__55216),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    Odrv4 I__11293 (
            .O(N__55213),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    LocalMux I__11292 (
            .O(N__55210),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    LocalMux I__11291 (
            .O(N__55207),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    LocalMux I__11290 (
            .O(N__55204),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ));
    InMux I__11289 (
            .O(N__55189),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17747 ));
    InMux I__11288 (
            .O(N__55186),
            .I(N__55183));
    LocalMux I__11287 (
            .O(N__55183),
            .I(N__55176));
    InMux I__11286 (
            .O(N__55182),
            .I(N__55173));
    InMux I__11285 (
            .O(N__55181),
            .I(N__55170));
    CascadeMux I__11284 (
            .O(N__55180),
            .I(N__55167));
    InMux I__11283 (
            .O(N__55179),
            .I(N__55163));
    Span4Mux_h I__11282 (
            .O(N__55176),
            .I(N__55156));
    LocalMux I__11281 (
            .O(N__55173),
            .I(N__55156));
    LocalMux I__11280 (
            .O(N__55170),
            .I(N__55156));
    InMux I__11279 (
            .O(N__55167),
            .I(N__55152));
    CascadeMux I__11278 (
            .O(N__55166),
            .I(N__55147));
    LocalMux I__11277 (
            .O(N__55163),
            .I(N__55144));
    Span4Mux_v I__11276 (
            .O(N__55156),
            .I(N__55141));
    InMux I__11275 (
            .O(N__55155),
            .I(N__55138));
    LocalMux I__11274 (
            .O(N__55152),
            .I(N__55135));
    InMux I__11273 (
            .O(N__55151),
            .I(N__55132));
    InMux I__11272 (
            .O(N__55150),
            .I(N__55129));
    InMux I__11271 (
            .O(N__55147),
            .I(N__55126));
    Span4Mux_v I__11270 (
            .O(N__55144),
            .I(N__55115));
    Span4Mux_h I__11269 (
            .O(N__55141),
            .I(N__55115));
    LocalMux I__11268 (
            .O(N__55138),
            .I(N__55115));
    Span4Mux_h I__11267 (
            .O(N__55135),
            .I(N__55106));
    LocalMux I__11266 (
            .O(N__55132),
            .I(N__55106));
    LocalMux I__11265 (
            .O(N__55129),
            .I(N__55106));
    LocalMux I__11264 (
            .O(N__55126),
            .I(N__55106));
    InMux I__11263 (
            .O(N__55125),
            .I(N__55103));
    InMux I__11262 (
            .O(N__55124),
            .I(N__55100));
    InMux I__11261 (
            .O(N__55123),
            .I(N__55097));
    InMux I__11260 (
            .O(N__55122),
            .I(N__55094));
    Span4Mux_v I__11259 (
            .O(N__55115),
            .I(N__55090));
    Span4Mux_v I__11258 (
            .O(N__55106),
            .I(N__55084));
    LocalMux I__11257 (
            .O(N__55103),
            .I(N__55084));
    LocalMux I__11256 (
            .O(N__55100),
            .I(N__55077));
    LocalMux I__11255 (
            .O(N__55097),
            .I(N__55077));
    LocalMux I__11254 (
            .O(N__55094),
            .I(N__55077));
    InMux I__11253 (
            .O(N__55093),
            .I(N__55074));
    Span4Mux_h I__11252 (
            .O(N__55090),
            .I(N__55070));
    InMux I__11251 (
            .O(N__55089),
            .I(N__55067));
    Span4Mux_v I__11250 (
            .O(N__55084),
            .I(N__55060));
    Span4Mux_v I__11249 (
            .O(N__55077),
            .I(N__55060));
    LocalMux I__11248 (
            .O(N__55074),
            .I(N__55060));
    InMux I__11247 (
            .O(N__55073),
            .I(N__55057));
    Odrv4 I__11246 (
            .O(N__55070),
            .I(n141));
    LocalMux I__11245 (
            .O(N__55067),
            .I(n141));
    Odrv4 I__11244 (
            .O(N__55060),
            .I(n141));
    LocalMux I__11243 (
            .O(N__55057),
            .I(n141));
    CascadeMux I__11242 (
            .O(N__55048),
            .I(N__55045));
    InMux I__11241 (
            .O(N__55045),
            .I(N__55042));
    LocalMux I__11240 (
            .O(N__55042),
            .I(N__55039));
    Span4Mux_h I__11239 (
            .O(N__55039),
            .I(N__55036));
    Odrv4 I__11238 (
            .O(N__55036),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429 ));
    InMux I__11237 (
            .O(N__55033),
            .I(N__55027));
    InMux I__11236 (
            .O(N__55032),
            .I(N__55027));
    LocalMux I__11235 (
            .O(N__55027),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n691 ));
    InMux I__11234 (
            .O(N__55024),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17748 ));
    InMux I__11233 (
            .O(N__55021),
            .I(N__55018));
    LocalMux I__11232 (
            .O(N__55018),
            .I(N__55015));
    Span12Mux_v I__11231 (
            .O(N__55015),
            .I(N__55012));
    Odrv12 I__11230 (
            .O(N__55012),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427 ));
    CascadeMux I__11229 (
            .O(N__55009),
            .I(N__55006));
    InMux I__11228 (
            .O(N__55006),
            .I(N__55002));
    CascadeMux I__11227 (
            .O(N__55005),
            .I(N__54998));
    LocalMux I__11226 (
            .O(N__55002),
            .I(N__54993));
    InMux I__11225 (
            .O(N__55001),
            .I(N__54990));
    InMux I__11224 (
            .O(N__54998),
            .I(N__54984));
    InMux I__11223 (
            .O(N__54997),
            .I(N__54981));
    InMux I__11222 (
            .O(N__54996),
            .I(N__54978));
    Span4Mux_v I__11221 (
            .O(N__54993),
            .I(N__54973));
    LocalMux I__11220 (
            .O(N__54990),
            .I(N__54973));
    InMux I__11219 (
            .O(N__54989),
            .I(N__54970));
    InMux I__11218 (
            .O(N__54988),
            .I(N__54966));
    InMux I__11217 (
            .O(N__54987),
            .I(N__54963));
    LocalMux I__11216 (
            .O(N__54984),
            .I(N__54960));
    LocalMux I__11215 (
            .O(N__54981),
            .I(N__54955));
    LocalMux I__11214 (
            .O(N__54978),
            .I(N__54952));
    Span4Mux_v I__11213 (
            .O(N__54973),
            .I(N__54947));
    LocalMux I__11212 (
            .O(N__54970),
            .I(N__54947));
    InMux I__11211 (
            .O(N__54969),
            .I(N__54942));
    LocalMux I__11210 (
            .O(N__54966),
            .I(N__54935));
    LocalMux I__11209 (
            .O(N__54963),
            .I(N__54935));
    Span4Mux_v I__11208 (
            .O(N__54960),
            .I(N__54932));
    InMux I__11207 (
            .O(N__54959),
            .I(N__54929));
    InMux I__11206 (
            .O(N__54958),
            .I(N__54926));
    Span4Mux_h I__11205 (
            .O(N__54955),
            .I(N__54923));
    Span4Mux_h I__11204 (
            .O(N__54952),
            .I(N__54918));
    Span4Mux_h I__11203 (
            .O(N__54947),
            .I(N__54918));
    InMux I__11202 (
            .O(N__54946),
            .I(N__54915));
    CascadeMux I__11201 (
            .O(N__54945),
            .I(N__54911));
    LocalMux I__11200 (
            .O(N__54942),
            .I(N__54908));
    InMux I__11199 (
            .O(N__54941),
            .I(N__54905));
    InMux I__11198 (
            .O(N__54940),
            .I(N__54902));
    Span4Mux_v I__11197 (
            .O(N__54935),
            .I(N__54895));
    Span4Mux_h I__11196 (
            .O(N__54932),
            .I(N__54895));
    LocalMux I__11195 (
            .O(N__54929),
            .I(N__54895));
    LocalMux I__11194 (
            .O(N__54926),
            .I(N__54886));
    Sp12to4 I__11193 (
            .O(N__54923),
            .I(N__54886));
    Sp12to4 I__11192 (
            .O(N__54918),
            .I(N__54886));
    LocalMux I__11191 (
            .O(N__54915),
            .I(N__54886));
    InMux I__11190 (
            .O(N__54914),
            .I(N__54883));
    InMux I__11189 (
            .O(N__54911),
            .I(N__54880));
    Span4Mux_v I__11188 (
            .O(N__54908),
            .I(N__54873));
    LocalMux I__11187 (
            .O(N__54905),
            .I(N__54873));
    LocalMux I__11186 (
            .O(N__54902),
            .I(N__54873));
    Odrv4 I__11185 (
            .O(N__54895),
            .I(n146));
    Odrv12 I__11184 (
            .O(N__54886),
            .I(n146));
    LocalMux I__11183 (
            .O(N__54883),
            .I(n146));
    LocalMux I__11182 (
            .O(N__54880),
            .I(n146));
    Odrv4 I__11181 (
            .O(N__54873),
            .I(n146));
    CascadeMux I__11180 (
            .O(N__54862),
            .I(N__54859));
    InMux I__11179 (
            .O(N__54859),
            .I(N__54856));
    LocalMux I__11178 (
            .O(N__54856),
            .I(N__54853));
    Span4Mux_v I__11177 (
            .O(N__54853),
            .I(N__54850));
    Odrv4 I__11176 (
            .O(N__54850),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n742 ));
    InMux I__11175 (
            .O(N__54847),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17749 ));
    InMux I__11174 (
            .O(N__54844),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n743 ));
    CascadeMux I__11173 (
            .O(N__54841),
            .I(N__54838));
    InMux I__11172 (
            .O(N__54838),
            .I(N__54835));
    LocalMux I__11171 (
            .O(N__54835),
            .I(N__54832));
    Span4Mux_h I__11170 (
            .O(N__54832),
            .I(N__54829));
    Odrv4 I__11169 (
            .O(N__54829),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO ));
    InMux I__11168 (
            .O(N__54826),
            .I(N__54823));
    LocalMux I__11167 (
            .O(N__54823),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n57 ));
    InMux I__11166 (
            .O(N__54820),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17736 ));
    InMux I__11165 (
            .O(N__54817),
            .I(N__54814));
    LocalMux I__11164 (
            .O(N__54814),
            .I(N__54810));
    CascadeMux I__11163 (
            .O(N__54813),
            .I(N__54807));
    Span4Mux_v I__11162 (
            .O(N__54810),
            .I(N__54793));
    InMux I__11161 (
            .O(N__54807),
            .I(N__54790));
    CascadeMux I__11160 (
            .O(N__54806),
            .I(N__54787));
    CascadeMux I__11159 (
            .O(N__54805),
            .I(N__54784));
    CascadeMux I__11158 (
            .O(N__54804),
            .I(N__54781));
    CascadeMux I__11157 (
            .O(N__54803),
            .I(N__54778));
    CascadeMux I__11156 (
            .O(N__54802),
            .I(N__54775));
    InMux I__11155 (
            .O(N__54801),
            .I(N__54765));
    CascadeMux I__11154 (
            .O(N__54800),
            .I(N__54762));
    CascadeMux I__11153 (
            .O(N__54799),
            .I(N__54758));
    CascadeMux I__11152 (
            .O(N__54798),
            .I(N__54754));
    CascadeMux I__11151 (
            .O(N__54797),
            .I(N__54751));
    CascadeMux I__11150 (
            .O(N__54796),
            .I(N__54747));
    Span4Mux_h I__11149 (
            .O(N__54793),
            .I(N__54742));
    LocalMux I__11148 (
            .O(N__54790),
            .I(N__54742));
    InMux I__11147 (
            .O(N__54787),
            .I(N__54739));
    InMux I__11146 (
            .O(N__54784),
            .I(N__54736));
    InMux I__11145 (
            .O(N__54781),
            .I(N__54733));
    InMux I__11144 (
            .O(N__54778),
            .I(N__54730));
    InMux I__11143 (
            .O(N__54775),
            .I(N__54727));
    CascadeMux I__11142 (
            .O(N__54774),
            .I(N__54724));
    CascadeMux I__11141 (
            .O(N__54773),
            .I(N__54721));
    CascadeMux I__11140 (
            .O(N__54772),
            .I(N__54718));
    CascadeMux I__11139 (
            .O(N__54771),
            .I(N__54715));
    CascadeMux I__11138 (
            .O(N__54770),
            .I(N__54710));
    CascadeMux I__11137 (
            .O(N__54769),
            .I(N__54706));
    CascadeMux I__11136 (
            .O(N__54768),
            .I(N__54702));
    LocalMux I__11135 (
            .O(N__54765),
            .I(N__54699));
    InMux I__11134 (
            .O(N__54762),
            .I(N__54696));
    InMux I__11133 (
            .O(N__54761),
            .I(N__54681));
    InMux I__11132 (
            .O(N__54758),
            .I(N__54681));
    InMux I__11131 (
            .O(N__54757),
            .I(N__54681));
    InMux I__11130 (
            .O(N__54754),
            .I(N__54681));
    InMux I__11129 (
            .O(N__54751),
            .I(N__54681));
    InMux I__11128 (
            .O(N__54750),
            .I(N__54681));
    InMux I__11127 (
            .O(N__54747),
            .I(N__54681));
    Span4Mux_v I__11126 (
            .O(N__54742),
            .I(N__54675));
    LocalMux I__11125 (
            .O(N__54739),
            .I(N__54675));
    LocalMux I__11124 (
            .O(N__54736),
            .I(N__54672));
    LocalMux I__11123 (
            .O(N__54733),
            .I(N__54665));
    LocalMux I__11122 (
            .O(N__54730),
            .I(N__54665));
    LocalMux I__11121 (
            .O(N__54727),
            .I(N__54665));
    InMux I__11120 (
            .O(N__54724),
            .I(N__54662));
    InMux I__11119 (
            .O(N__54721),
            .I(N__54659));
    InMux I__11118 (
            .O(N__54718),
            .I(N__54656));
    InMux I__11117 (
            .O(N__54715),
            .I(N__54653));
    CascadeMux I__11116 (
            .O(N__54714),
            .I(N__54650));
    InMux I__11115 (
            .O(N__54713),
            .I(N__54637));
    InMux I__11114 (
            .O(N__54710),
            .I(N__54637));
    InMux I__11113 (
            .O(N__54709),
            .I(N__54637));
    InMux I__11112 (
            .O(N__54706),
            .I(N__54637));
    InMux I__11111 (
            .O(N__54705),
            .I(N__54637));
    InMux I__11110 (
            .O(N__54702),
            .I(N__54637));
    Span4Mux_v I__11109 (
            .O(N__54699),
            .I(N__54632));
    LocalMux I__11108 (
            .O(N__54696),
            .I(N__54632));
    LocalMux I__11107 (
            .O(N__54681),
            .I(N__54629));
    CascadeMux I__11106 (
            .O(N__54680),
            .I(N__54626));
    Span4Mux_v I__11105 (
            .O(N__54675),
            .I(N__54620));
    Span4Mux_h I__11104 (
            .O(N__54672),
            .I(N__54620));
    Span4Mux_v I__11103 (
            .O(N__54665),
            .I(N__54609));
    LocalMux I__11102 (
            .O(N__54662),
            .I(N__54609));
    LocalMux I__11101 (
            .O(N__54659),
            .I(N__54609));
    LocalMux I__11100 (
            .O(N__54656),
            .I(N__54609));
    LocalMux I__11099 (
            .O(N__54653),
            .I(N__54609));
    InMux I__11098 (
            .O(N__54650),
            .I(N__54606));
    LocalMux I__11097 (
            .O(N__54637),
            .I(N__54599));
    Span4Mux_v I__11096 (
            .O(N__54632),
            .I(N__54599));
    Span4Mux_v I__11095 (
            .O(N__54629),
            .I(N__54599));
    InMux I__11094 (
            .O(N__54626),
            .I(N__54596));
    CascadeMux I__11093 (
            .O(N__54625),
            .I(N__54593));
    Span4Mux_v I__11092 (
            .O(N__54620),
            .I(N__54590));
    Span4Mux_v I__11091 (
            .O(N__54609),
            .I(N__54585));
    LocalMux I__11090 (
            .O(N__54606),
            .I(N__54585));
    Span4Mux_h I__11089 (
            .O(N__54599),
            .I(N__54580));
    LocalMux I__11088 (
            .O(N__54596),
            .I(N__54580));
    InMux I__11087 (
            .O(N__54593),
            .I(N__54577));
    Odrv4 I__11086 (
            .O(N__54590),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n108 ));
    Odrv4 I__11085 (
            .O(N__54585),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n108 ));
    Odrv4 I__11084 (
            .O(N__54580),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n108 ));
    LocalMux I__11083 (
            .O(N__54577),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n108 ));
    CascadeMux I__11082 (
            .O(N__54568),
            .I(N__54565));
    InMux I__11081 (
            .O(N__54565),
            .I(N__54562));
    LocalMux I__11080 (
            .O(N__54562),
            .I(N__54559));
    Span4Mux_v I__11079 (
            .O(N__54559),
            .I(N__54556));
    Odrv4 I__11078 (
            .O(N__54556),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n106 ));
    InMux I__11077 (
            .O(N__54553),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17737 ));
    InMux I__11076 (
            .O(N__54550),
            .I(N__54547));
    LocalMux I__11075 (
            .O(N__54547),
            .I(N__54544));
    Span4Mux_v I__11074 (
            .O(N__54544),
            .I(N__54541));
    Odrv4 I__11073 (
            .O(N__54541),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369 ));
    CascadeMux I__11072 (
            .O(N__54538),
            .I(N__54535));
    InMux I__11071 (
            .O(N__54535),
            .I(N__54531));
    CascadeMux I__11070 (
            .O(N__54534),
            .I(N__54527));
    LocalMux I__11069 (
            .O(N__54531),
            .I(N__54522));
    CascadeMux I__11068 (
            .O(N__54530),
            .I(N__54518));
    InMux I__11067 (
            .O(N__54527),
            .I(N__54513));
    CascadeMux I__11066 (
            .O(N__54526),
            .I(N__54505));
    CascadeMux I__11065 (
            .O(N__54525),
            .I(N__54502));
    Span4Mux_v I__11064 (
            .O(N__54522),
            .I(N__54494));
    InMux I__11063 (
            .O(N__54521),
            .I(N__54491));
    InMux I__11062 (
            .O(N__54518),
            .I(N__54488));
    CascadeMux I__11061 (
            .O(N__54517),
            .I(N__54485));
    CascadeMux I__11060 (
            .O(N__54516),
            .I(N__54482));
    LocalMux I__11059 (
            .O(N__54513),
            .I(N__54477));
    CascadeMux I__11058 (
            .O(N__54512),
            .I(N__54474));
    CascadeMux I__11057 (
            .O(N__54511),
            .I(N__54470));
    CascadeMux I__11056 (
            .O(N__54510),
            .I(N__54466));
    CascadeMux I__11055 (
            .O(N__54509),
            .I(N__54463));
    InMux I__11054 (
            .O(N__54508),
            .I(N__54460));
    InMux I__11053 (
            .O(N__54505),
            .I(N__54457));
    InMux I__11052 (
            .O(N__54502),
            .I(N__54454));
    CascadeMux I__11051 (
            .O(N__54501),
            .I(N__54451));
    CascadeMux I__11050 (
            .O(N__54500),
            .I(N__54446));
    CascadeMux I__11049 (
            .O(N__54499),
            .I(N__54442));
    CascadeMux I__11048 (
            .O(N__54498),
            .I(N__54438));
    CascadeMux I__11047 (
            .O(N__54497),
            .I(N__54434));
    Span4Mux_h I__11046 (
            .O(N__54494),
            .I(N__54426));
    LocalMux I__11045 (
            .O(N__54491),
            .I(N__54426));
    LocalMux I__11044 (
            .O(N__54488),
            .I(N__54426));
    InMux I__11043 (
            .O(N__54485),
            .I(N__54423));
    InMux I__11042 (
            .O(N__54482),
            .I(N__54420));
    CascadeMux I__11041 (
            .O(N__54481),
            .I(N__54417));
    CascadeMux I__11040 (
            .O(N__54480),
            .I(N__54414));
    Span4Mux_v I__11039 (
            .O(N__54477),
            .I(N__54411));
    InMux I__11038 (
            .O(N__54474),
            .I(N__54400));
    InMux I__11037 (
            .O(N__54473),
            .I(N__54400));
    InMux I__11036 (
            .O(N__54470),
            .I(N__54400));
    InMux I__11035 (
            .O(N__54469),
            .I(N__54400));
    InMux I__11034 (
            .O(N__54466),
            .I(N__54400));
    InMux I__11033 (
            .O(N__54463),
            .I(N__54397));
    LocalMux I__11032 (
            .O(N__54460),
            .I(N__54390));
    LocalMux I__11031 (
            .O(N__54457),
            .I(N__54390));
    LocalMux I__11030 (
            .O(N__54454),
            .I(N__54390));
    InMux I__11029 (
            .O(N__54451),
            .I(N__54387));
    InMux I__11028 (
            .O(N__54450),
            .I(N__54383));
    InMux I__11027 (
            .O(N__54449),
            .I(N__54374));
    InMux I__11026 (
            .O(N__54446),
            .I(N__54374));
    InMux I__11025 (
            .O(N__54445),
            .I(N__54374));
    InMux I__11024 (
            .O(N__54442),
            .I(N__54374));
    InMux I__11023 (
            .O(N__54441),
            .I(N__54365));
    InMux I__11022 (
            .O(N__54438),
            .I(N__54365));
    InMux I__11021 (
            .O(N__54437),
            .I(N__54365));
    InMux I__11020 (
            .O(N__54434),
            .I(N__54365));
    InMux I__11019 (
            .O(N__54433),
            .I(N__54362));
    Span4Mux_v I__11018 (
            .O(N__54426),
            .I(N__54355));
    LocalMux I__11017 (
            .O(N__54423),
            .I(N__54355));
    LocalMux I__11016 (
            .O(N__54420),
            .I(N__54355));
    InMux I__11015 (
            .O(N__54417),
            .I(N__54352));
    InMux I__11014 (
            .O(N__54414),
            .I(N__54349));
    Span4Mux_v I__11013 (
            .O(N__54411),
            .I(N__54344));
    LocalMux I__11012 (
            .O(N__54400),
            .I(N__54344));
    LocalMux I__11011 (
            .O(N__54397),
            .I(N__54341));
    Span4Mux_v I__11010 (
            .O(N__54390),
            .I(N__54336));
    LocalMux I__11009 (
            .O(N__54387),
            .I(N__54336));
    CascadeMux I__11008 (
            .O(N__54386),
            .I(N__54333));
    LocalMux I__11007 (
            .O(N__54383),
            .I(N__54324));
    LocalMux I__11006 (
            .O(N__54374),
            .I(N__54324));
    LocalMux I__11005 (
            .O(N__54365),
            .I(N__54324));
    LocalMux I__11004 (
            .O(N__54362),
            .I(N__54324));
    Span4Mux_v I__11003 (
            .O(N__54355),
            .I(N__54317));
    LocalMux I__11002 (
            .O(N__54352),
            .I(N__54317));
    LocalMux I__11001 (
            .O(N__54349),
            .I(N__54317));
    Span4Mux_v I__11000 (
            .O(N__54344),
            .I(N__54312));
    Span4Mux_v I__10999 (
            .O(N__54341),
            .I(N__54312));
    Span4Mux_v I__10998 (
            .O(N__54336),
            .I(N__54309));
    InMux I__10997 (
            .O(N__54333),
            .I(N__54306));
    Span12Mux_h I__10996 (
            .O(N__54324),
            .I(N__54303));
    Span4Mux_v I__10995 (
            .O(N__54317),
            .I(N__54300));
    Sp12to4 I__10994 (
            .O(N__54312),
            .I(N__54293));
    Sp12to4 I__10993 (
            .O(N__54309),
            .I(N__54293));
    LocalMux I__10992 (
            .O(N__54306),
            .I(N__54293));
    Odrv12 I__10991 (
            .O(N__54303),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n111 ));
    Odrv4 I__10990 (
            .O(N__54300),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n111 ));
    Odrv12 I__10989 (
            .O(N__54293),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n111 ));
    InMux I__10988 (
            .O(N__54286),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17738 ));
    InMux I__10987 (
            .O(N__54283),
            .I(N__54280));
    LocalMux I__10986 (
            .O(N__54280),
            .I(N__54277));
    Span4Mux_h I__10985 (
            .O(N__54277),
            .I(N__54274));
    Odrv4 I__10984 (
            .O(N__54274),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361 ));
    CascadeMux I__10983 (
            .O(N__54271),
            .I(N__54268));
    InMux I__10982 (
            .O(N__54268),
            .I(N__54265));
    LocalMux I__10981 (
            .O(N__54265),
            .I(N__54261));
    CascadeMux I__10980 (
            .O(N__54264),
            .I(N__54258));
    Span4Mux_v I__10979 (
            .O(N__54261),
            .I(N__54245));
    InMux I__10978 (
            .O(N__54258),
            .I(N__54242));
    CascadeMux I__10977 (
            .O(N__54257),
            .I(N__54239));
    CascadeMux I__10976 (
            .O(N__54256),
            .I(N__54236));
    CascadeMux I__10975 (
            .O(N__54255),
            .I(N__54233));
    CascadeMux I__10974 (
            .O(N__54254),
            .I(N__54229));
    CascadeMux I__10973 (
            .O(N__54253),
            .I(N__54225));
    CascadeMux I__10972 (
            .O(N__54252),
            .I(N__54221));
    CascadeMux I__10971 (
            .O(N__54251),
            .I(N__54217));
    CascadeMux I__10970 (
            .O(N__54250),
            .I(N__54214));
    CascadeMux I__10969 (
            .O(N__54249),
            .I(N__54211));
    CascadeMux I__10968 (
            .O(N__54248),
            .I(N__54208));
    Span4Mux_v I__10967 (
            .O(N__54245),
            .I(N__54202));
    LocalMux I__10966 (
            .O(N__54242),
            .I(N__54202));
    InMux I__10965 (
            .O(N__54239),
            .I(N__54199));
    InMux I__10964 (
            .O(N__54236),
            .I(N__54196));
    InMux I__10963 (
            .O(N__54233),
            .I(N__54190));
    InMux I__10962 (
            .O(N__54232),
            .I(N__54177));
    InMux I__10961 (
            .O(N__54229),
            .I(N__54177));
    InMux I__10960 (
            .O(N__54228),
            .I(N__54177));
    InMux I__10959 (
            .O(N__54225),
            .I(N__54177));
    InMux I__10958 (
            .O(N__54224),
            .I(N__54177));
    InMux I__10957 (
            .O(N__54221),
            .I(N__54177));
    CascadeMux I__10956 (
            .O(N__54220),
            .I(N__54172));
    InMux I__10955 (
            .O(N__54217),
            .I(N__54169));
    InMux I__10954 (
            .O(N__54214),
            .I(N__54166));
    InMux I__10953 (
            .O(N__54211),
            .I(N__54163));
    InMux I__10952 (
            .O(N__54208),
            .I(N__54160));
    CascadeMux I__10951 (
            .O(N__54207),
            .I(N__54157));
    Span4Mux_h I__10950 (
            .O(N__54202),
            .I(N__54153));
    LocalMux I__10949 (
            .O(N__54199),
            .I(N__54148));
    LocalMux I__10948 (
            .O(N__54196),
            .I(N__54148));
    CascadeMux I__10947 (
            .O(N__54195),
            .I(N__54145));
    CascadeMux I__10946 (
            .O(N__54194),
            .I(N__54142));
    CascadeMux I__10945 (
            .O(N__54193),
            .I(N__54139));
    LocalMux I__10944 (
            .O(N__54190),
            .I(N__54132));
    LocalMux I__10943 (
            .O(N__54177),
            .I(N__54129));
    InMux I__10942 (
            .O(N__54176),
            .I(N__54126));
    InMux I__10941 (
            .O(N__54175),
            .I(N__54123));
    InMux I__10940 (
            .O(N__54172),
            .I(N__54120));
    LocalMux I__10939 (
            .O(N__54169),
            .I(N__54111));
    LocalMux I__10938 (
            .O(N__54166),
            .I(N__54111));
    LocalMux I__10937 (
            .O(N__54163),
            .I(N__54111));
    LocalMux I__10936 (
            .O(N__54160),
            .I(N__54111));
    InMux I__10935 (
            .O(N__54157),
            .I(N__54108));
    CascadeMux I__10934 (
            .O(N__54156),
            .I(N__54105));
    Span4Mux_v I__10933 (
            .O(N__54153),
            .I(N__54100));
    Span4Mux_h I__10932 (
            .O(N__54148),
            .I(N__54100));
    InMux I__10931 (
            .O(N__54145),
            .I(N__54091));
    InMux I__10930 (
            .O(N__54142),
            .I(N__54091));
    InMux I__10929 (
            .O(N__54139),
            .I(N__54091));
    InMux I__10928 (
            .O(N__54138),
            .I(N__54091));
    CascadeMux I__10927 (
            .O(N__54137),
            .I(N__54088));
    CascadeMux I__10926 (
            .O(N__54136),
            .I(N__54085));
    CascadeMux I__10925 (
            .O(N__54135),
            .I(N__54081));
    Span4Mux_h I__10924 (
            .O(N__54132),
            .I(N__54077));
    Span4Mux_v I__10923 (
            .O(N__54129),
            .I(N__54070));
    LocalMux I__10922 (
            .O(N__54126),
            .I(N__54070));
    LocalMux I__10921 (
            .O(N__54123),
            .I(N__54070));
    LocalMux I__10920 (
            .O(N__54120),
            .I(N__54063));
    Span4Mux_v I__10919 (
            .O(N__54111),
            .I(N__54063));
    LocalMux I__10918 (
            .O(N__54108),
            .I(N__54063));
    InMux I__10917 (
            .O(N__54105),
            .I(N__54060));
    Span4Mux_v I__10916 (
            .O(N__54100),
            .I(N__54055));
    LocalMux I__10915 (
            .O(N__54091),
            .I(N__54055));
    InMux I__10914 (
            .O(N__54088),
            .I(N__54046));
    InMux I__10913 (
            .O(N__54085),
            .I(N__54046));
    InMux I__10912 (
            .O(N__54084),
            .I(N__54046));
    InMux I__10911 (
            .O(N__54081),
            .I(N__54046));
    CascadeMux I__10910 (
            .O(N__54080),
            .I(N__54043));
    Span4Mux_v I__10909 (
            .O(N__54077),
            .I(N__54038));
    Span4Mux_h I__10908 (
            .O(N__54070),
            .I(N__54038));
    Span4Mux_v I__10907 (
            .O(N__54063),
            .I(N__54033));
    LocalMux I__10906 (
            .O(N__54060),
            .I(N__54033));
    Sp12to4 I__10905 (
            .O(N__54055),
            .I(N__54028));
    LocalMux I__10904 (
            .O(N__54046),
            .I(N__54028));
    InMux I__10903 (
            .O(N__54043),
            .I(N__54025));
    Odrv4 I__10902 (
            .O(N__54038),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n114 ));
    Odrv4 I__10901 (
            .O(N__54033),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n114 ));
    Odrv12 I__10900 (
            .O(N__54028),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n114 ));
    LocalMux I__10899 (
            .O(N__54025),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n114 ));
    InMux I__10898 (
            .O(N__54016),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17739 ));
    InMux I__10897 (
            .O(N__54013),
            .I(N__54010));
    LocalMux I__10896 (
            .O(N__54010),
            .I(N__54007));
    Span4Mux_h I__10895 (
            .O(N__54007),
            .I(N__54004));
    Odrv4 I__10894 (
            .O(N__54004),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n253 ));
    CascadeMux I__10893 (
            .O(N__54001),
            .I(N__53996));
    CascadeMux I__10892 (
            .O(N__54000),
            .I(N__53993));
    CascadeMux I__10891 (
            .O(N__53999),
            .I(N__53987));
    InMux I__10890 (
            .O(N__53996),
            .I(N__53983));
    InMux I__10889 (
            .O(N__53993),
            .I(N__53980));
    CascadeMux I__10888 (
            .O(N__53992),
            .I(N__53977));
    CascadeMux I__10887 (
            .O(N__53991),
            .I(N__53974));
    CascadeMux I__10886 (
            .O(N__53990),
            .I(N__53971));
    InMux I__10885 (
            .O(N__53987),
            .I(N__53966));
    CascadeMux I__10884 (
            .O(N__53986),
            .I(N__53963));
    LocalMux I__10883 (
            .O(N__53983),
            .I(N__53958));
    LocalMux I__10882 (
            .O(N__53980),
            .I(N__53958));
    InMux I__10881 (
            .O(N__53977),
            .I(N__53955));
    InMux I__10880 (
            .O(N__53974),
            .I(N__53952));
    InMux I__10879 (
            .O(N__53971),
            .I(N__53949));
    CascadeMux I__10878 (
            .O(N__53970),
            .I(N__53946));
    CascadeMux I__10877 (
            .O(N__53969),
            .I(N__53943));
    LocalMux I__10876 (
            .O(N__53966),
            .I(N__53934));
    InMux I__10875 (
            .O(N__53963),
            .I(N__53931));
    Span4Mux_v I__10874 (
            .O(N__53958),
            .I(N__53922));
    LocalMux I__10873 (
            .O(N__53955),
            .I(N__53922));
    LocalMux I__10872 (
            .O(N__53952),
            .I(N__53922));
    LocalMux I__10871 (
            .O(N__53949),
            .I(N__53922));
    InMux I__10870 (
            .O(N__53946),
            .I(N__53919));
    InMux I__10869 (
            .O(N__53943),
            .I(N__53916));
    CascadeMux I__10868 (
            .O(N__53942),
            .I(N__53912));
    CascadeMux I__10867 (
            .O(N__53941),
            .I(N__53908));
    CascadeMux I__10866 (
            .O(N__53940),
            .I(N__53904));
    CascadeMux I__10865 (
            .O(N__53939),
            .I(N__53900));
    CascadeMux I__10864 (
            .O(N__53938),
            .I(N__53897));
    CascadeMux I__10863 (
            .O(N__53937),
            .I(N__53894));
    Span4Mux_v I__10862 (
            .O(N__53934),
            .I(N__53889));
    LocalMux I__10861 (
            .O(N__53931),
            .I(N__53889));
    Span4Mux_v I__10860 (
            .O(N__53922),
            .I(N__53876));
    LocalMux I__10859 (
            .O(N__53919),
            .I(N__53876));
    LocalMux I__10858 (
            .O(N__53916),
            .I(N__53873));
    InMux I__10857 (
            .O(N__53915),
            .I(N__53870));
    InMux I__10856 (
            .O(N__53912),
            .I(N__53867));
    InMux I__10855 (
            .O(N__53911),
            .I(N__53854));
    InMux I__10854 (
            .O(N__53908),
            .I(N__53854));
    InMux I__10853 (
            .O(N__53907),
            .I(N__53854));
    InMux I__10852 (
            .O(N__53904),
            .I(N__53854));
    InMux I__10851 (
            .O(N__53903),
            .I(N__53854));
    InMux I__10850 (
            .O(N__53900),
            .I(N__53854));
    InMux I__10849 (
            .O(N__53897),
            .I(N__53851));
    InMux I__10848 (
            .O(N__53894),
            .I(N__53848));
    Span4Mux_h I__10847 (
            .O(N__53889),
            .I(N__53845));
    InMux I__10846 (
            .O(N__53888),
            .I(N__53842));
    CascadeMux I__10845 (
            .O(N__53887),
            .I(N__53839));
    CascadeMux I__10844 (
            .O(N__53886),
            .I(N__53836));
    CascadeMux I__10843 (
            .O(N__53885),
            .I(N__53833));
    CascadeMux I__10842 (
            .O(N__53884),
            .I(N__53829));
    CascadeMux I__10841 (
            .O(N__53883),
            .I(N__53826));
    CascadeMux I__10840 (
            .O(N__53882),
            .I(N__53823));
    CascadeMux I__10839 (
            .O(N__53881),
            .I(N__53820));
    Span4Mux_v I__10838 (
            .O(N__53876),
            .I(N__53816));
    Span4Mux_v I__10837 (
            .O(N__53873),
            .I(N__53805));
    LocalMux I__10836 (
            .O(N__53870),
            .I(N__53805));
    LocalMux I__10835 (
            .O(N__53867),
            .I(N__53805));
    LocalMux I__10834 (
            .O(N__53854),
            .I(N__53805));
    LocalMux I__10833 (
            .O(N__53851),
            .I(N__53805));
    LocalMux I__10832 (
            .O(N__53848),
            .I(N__53802));
    Span4Mux_v I__10831 (
            .O(N__53845),
            .I(N__53799));
    LocalMux I__10830 (
            .O(N__53842),
            .I(N__53796));
    InMux I__10829 (
            .O(N__53839),
            .I(N__53785));
    InMux I__10828 (
            .O(N__53836),
            .I(N__53785));
    InMux I__10827 (
            .O(N__53833),
            .I(N__53785));
    InMux I__10826 (
            .O(N__53832),
            .I(N__53785));
    InMux I__10825 (
            .O(N__53829),
            .I(N__53785));
    InMux I__10824 (
            .O(N__53826),
            .I(N__53778));
    InMux I__10823 (
            .O(N__53823),
            .I(N__53778));
    InMux I__10822 (
            .O(N__53820),
            .I(N__53778));
    CascadeMux I__10821 (
            .O(N__53819),
            .I(N__53775));
    Span4Mux_h I__10820 (
            .O(N__53816),
            .I(N__53772));
    Span4Mux_v I__10819 (
            .O(N__53805),
            .I(N__53769));
    Span4Mux_h I__10818 (
            .O(N__53802),
            .I(N__53766));
    Span4Mux_v I__10817 (
            .O(N__53799),
            .I(N__53757));
    Span4Mux_h I__10816 (
            .O(N__53796),
            .I(N__53757));
    LocalMux I__10815 (
            .O(N__53785),
            .I(N__53757));
    LocalMux I__10814 (
            .O(N__53778),
            .I(N__53757));
    InMux I__10813 (
            .O(N__53775),
            .I(N__53754));
    Odrv4 I__10812 (
            .O(N__53772),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ));
    Odrv4 I__10811 (
            .O(N__53769),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ));
    Odrv4 I__10810 (
            .O(N__53766),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ));
    Odrv4 I__10809 (
            .O(N__53757),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ));
    LocalMux I__10808 (
            .O(N__53754),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ));
    InMux I__10807 (
            .O(N__53743),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17740 ));
    InMux I__10806 (
            .O(N__53740),
            .I(N__53737));
    LocalMux I__10805 (
            .O(N__53737),
            .I(N__53734));
    Span4Mux_h I__10804 (
            .O(N__53734),
            .I(N__53731));
    Odrv4 I__10803 (
            .O(N__53731),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364 ));
    CascadeMux I__10802 (
            .O(N__53728),
            .I(N__53725));
    InMux I__10801 (
            .O(N__53725),
            .I(N__53719));
    CascadeMux I__10800 (
            .O(N__53724),
            .I(N__53716));
    CascadeMux I__10799 (
            .O(N__53723),
            .I(N__53712));
    CascadeMux I__10798 (
            .O(N__53722),
            .I(N__53708));
    LocalMux I__10797 (
            .O(N__53719),
            .I(N__53702));
    InMux I__10796 (
            .O(N__53716),
            .I(N__53699));
    CascadeMux I__10795 (
            .O(N__53715),
            .I(N__53696));
    InMux I__10794 (
            .O(N__53712),
            .I(N__53690));
    CascadeMux I__10793 (
            .O(N__53711),
            .I(N__53687));
    InMux I__10792 (
            .O(N__53708),
            .I(N__53684));
    CascadeMux I__10791 (
            .O(N__53707),
            .I(N__53681));
    CascadeMux I__10790 (
            .O(N__53706),
            .I(N__53677));
    InMux I__10789 (
            .O(N__53705),
            .I(N__53674));
    Span4Mux_v I__10788 (
            .O(N__53702),
            .I(N__53669));
    LocalMux I__10787 (
            .O(N__53699),
            .I(N__53669));
    InMux I__10786 (
            .O(N__53696),
            .I(N__53666));
    CascadeMux I__10785 (
            .O(N__53695),
            .I(N__53662));
    CascadeMux I__10784 (
            .O(N__53694),
            .I(N__53658));
    CascadeMux I__10783 (
            .O(N__53693),
            .I(N__53654));
    LocalMux I__10782 (
            .O(N__53690),
            .I(N__53651));
    InMux I__10781 (
            .O(N__53687),
            .I(N__53647));
    LocalMux I__10780 (
            .O(N__53684),
            .I(N__53644));
    InMux I__10779 (
            .O(N__53681),
            .I(N__53641));
    InMux I__10778 (
            .O(N__53680),
            .I(N__53638));
    InMux I__10777 (
            .O(N__53677),
            .I(N__53633));
    LocalMux I__10776 (
            .O(N__53674),
            .I(N__53630));
    Span4Mux_h I__10775 (
            .O(N__53669),
            .I(N__53625));
    LocalMux I__10774 (
            .O(N__53666),
            .I(N__53625));
    InMux I__10773 (
            .O(N__53665),
            .I(N__53612));
    InMux I__10772 (
            .O(N__53662),
            .I(N__53612));
    InMux I__10771 (
            .O(N__53661),
            .I(N__53612));
    InMux I__10770 (
            .O(N__53658),
            .I(N__53612));
    InMux I__10769 (
            .O(N__53657),
            .I(N__53612));
    InMux I__10768 (
            .O(N__53654),
            .I(N__53612));
    Span4Mux_v I__10767 (
            .O(N__53651),
            .I(N__53604));
    InMux I__10766 (
            .O(N__53650),
            .I(N__53601));
    LocalMux I__10765 (
            .O(N__53647),
            .I(N__53592));
    Span4Mux_h I__10764 (
            .O(N__53644),
            .I(N__53592));
    LocalMux I__10763 (
            .O(N__53641),
            .I(N__53592));
    LocalMux I__10762 (
            .O(N__53638),
            .I(N__53592));
    InMux I__10761 (
            .O(N__53637),
            .I(N__53589));
    CascadeMux I__10760 (
            .O(N__53636),
            .I(N__53586));
    LocalMux I__10759 (
            .O(N__53633),
            .I(N__53582));
    Span4Mux_v I__10758 (
            .O(N__53630),
            .I(N__53575));
    Span4Mux_h I__10757 (
            .O(N__53625),
            .I(N__53575));
    LocalMux I__10756 (
            .O(N__53612),
            .I(N__53575));
    InMux I__10755 (
            .O(N__53611),
            .I(N__53572));
    CascadeMux I__10754 (
            .O(N__53610),
            .I(N__53569));
    CascadeMux I__10753 (
            .O(N__53609),
            .I(N__53564));
    CascadeMux I__10752 (
            .O(N__53608),
            .I(N__53560));
    CascadeMux I__10751 (
            .O(N__53607),
            .I(N__53556));
    Span4Mux_h I__10750 (
            .O(N__53604),
            .I(N__53547));
    LocalMux I__10749 (
            .O(N__53601),
            .I(N__53547));
    Span4Mux_v I__10748 (
            .O(N__53592),
            .I(N__53547));
    LocalMux I__10747 (
            .O(N__53589),
            .I(N__53547));
    InMux I__10746 (
            .O(N__53586),
            .I(N__53544));
    CascadeMux I__10745 (
            .O(N__53585),
            .I(N__53541));
    Span4Mux_v I__10744 (
            .O(N__53582),
            .I(N__53534));
    Span4Mux_v I__10743 (
            .O(N__53575),
            .I(N__53534));
    LocalMux I__10742 (
            .O(N__53572),
            .I(N__53534));
    InMux I__10741 (
            .O(N__53569),
            .I(N__53529));
    InMux I__10740 (
            .O(N__53568),
            .I(N__53529));
    InMux I__10739 (
            .O(N__53567),
            .I(N__53516));
    InMux I__10738 (
            .O(N__53564),
            .I(N__53516));
    InMux I__10737 (
            .O(N__53563),
            .I(N__53516));
    InMux I__10736 (
            .O(N__53560),
            .I(N__53516));
    InMux I__10735 (
            .O(N__53559),
            .I(N__53516));
    InMux I__10734 (
            .O(N__53556),
            .I(N__53516));
    Span4Mux_v I__10733 (
            .O(N__53547),
            .I(N__53511));
    LocalMux I__10732 (
            .O(N__53544),
            .I(N__53511));
    InMux I__10731 (
            .O(N__53541),
            .I(N__53508));
    Sp12to4 I__10730 (
            .O(N__53534),
            .I(N__53501));
    LocalMux I__10729 (
            .O(N__53529),
            .I(N__53501));
    LocalMux I__10728 (
            .O(N__53516),
            .I(N__53501));
    Odrv4 I__10727 (
            .O(N__53511),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n120 ));
    LocalMux I__10726 (
            .O(N__53508),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n120 ));
    Odrv12 I__10725 (
            .O(N__53501),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n120 ));
    InMux I__10724 (
            .O(N__53494),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17741 ));
    InMux I__10723 (
            .O(N__53491),
            .I(N__53488));
    LocalMux I__10722 (
            .O(N__53488),
            .I(N__53485));
    Span4Mux_v I__10721 (
            .O(N__53485),
            .I(N__53482));
    Odrv4 I__10720 (
            .O(N__53482),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n351 ));
    InMux I__10719 (
            .O(N__53479),
            .I(N__53475));
    CascadeMux I__10718 (
            .O(N__53478),
            .I(N__53471));
    LocalMux I__10717 (
            .O(N__53475),
            .I(N__53461));
    InMux I__10716 (
            .O(N__53474),
            .I(N__53458));
    InMux I__10715 (
            .O(N__53471),
            .I(N__53455));
    CascadeMux I__10714 (
            .O(N__53470),
            .I(N__53452));
    CascadeMux I__10713 (
            .O(N__53469),
            .I(N__53449));
    CascadeMux I__10712 (
            .O(N__53468),
            .I(N__53446));
    CascadeMux I__10711 (
            .O(N__53467),
            .I(N__53442));
    CascadeMux I__10710 (
            .O(N__53466),
            .I(N__53439));
    CascadeMux I__10709 (
            .O(N__53465),
            .I(N__53435));
    CascadeMux I__10708 (
            .O(N__53464),
            .I(N__53431));
    Span4Mux_v I__10707 (
            .O(N__53461),
            .I(N__53423));
    LocalMux I__10706 (
            .O(N__53458),
            .I(N__53420));
    LocalMux I__10705 (
            .O(N__53455),
            .I(N__53417));
    InMux I__10704 (
            .O(N__53452),
            .I(N__53414));
    InMux I__10703 (
            .O(N__53449),
            .I(N__53411));
    InMux I__10702 (
            .O(N__53446),
            .I(N__53405));
    InMux I__10701 (
            .O(N__53445),
            .I(N__53390));
    InMux I__10700 (
            .O(N__53442),
            .I(N__53390));
    InMux I__10699 (
            .O(N__53439),
            .I(N__53390));
    InMux I__10698 (
            .O(N__53438),
            .I(N__53390));
    InMux I__10697 (
            .O(N__53435),
            .I(N__53390));
    InMux I__10696 (
            .O(N__53434),
            .I(N__53390));
    InMux I__10695 (
            .O(N__53431),
            .I(N__53390));
    CascadeMux I__10694 (
            .O(N__53430),
            .I(N__53387));
    CascadeMux I__10693 (
            .O(N__53429),
            .I(N__53383));
    CascadeMux I__10692 (
            .O(N__53428),
            .I(N__53379));
    CascadeMux I__10691 (
            .O(N__53427),
            .I(N__53374));
    InMux I__10690 (
            .O(N__53426),
            .I(N__53370));
    Span4Mux_v I__10689 (
            .O(N__53423),
            .I(N__53364));
    Span4Mux_v I__10688 (
            .O(N__53420),
            .I(N__53364));
    Span4Mux_h I__10687 (
            .O(N__53417),
            .I(N__53359));
    LocalMux I__10686 (
            .O(N__53414),
            .I(N__53359));
    LocalMux I__10685 (
            .O(N__53411),
            .I(N__53356));
    CascadeMux I__10684 (
            .O(N__53410),
            .I(N__53353));
    CascadeMux I__10683 (
            .O(N__53409),
            .I(N__53350));
    CascadeMux I__10682 (
            .O(N__53408),
            .I(N__53347));
    LocalMux I__10681 (
            .O(N__53405),
            .I(N__53342));
    LocalMux I__10680 (
            .O(N__53390),
            .I(N__53342));
    InMux I__10679 (
            .O(N__53387),
            .I(N__53329));
    InMux I__10678 (
            .O(N__53386),
            .I(N__53329));
    InMux I__10677 (
            .O(N__53383),
            .I(N__53329));
    InMux I__10676 (
            .O(N__53382),
            .I(N__53329));
    InMux I__10675 (
            .O(N__53379),
            .I(N__53329));
    InMux I__10674 (
            .O(N__53378),
            .I(N__53329));
    InMux I__10673 (
            .O(N__53377),
            .I(N__53326));
    InMux I__10672 (
            .O(N__53374),
            .I(N__53323));
    CascadeMux I__10671 (
            .O(N__53373),
            .I(N__53320));
    LocalMux I__10670 (
            .O(N__53370),
            .I(N__53317));
    CascadeMux I__10669 (
            .O(N__53369),
            .I(N__53313));
    Span4Mux_h I__10668 (
            .O(N__53364),
            .I(N__53306));
    Span4Mux_v I__10667 (
            .O(N__53359),
            .I(N__53306));
    Span4Mux_v I__10666 (
            .O(N__53356),
            .I(N__53306));
    InMux I__10665 (
            .O(N__53353),
            .I(N__53303));
    InMux I__10664 (
            .O(N__53350),
            .I(N__53300));
    InMux I__10663 (
            .O(N__53347),
            .I(N__53297));
    Span4Mux_v I__10662 (
            .O(N__53342),
            .I(N__53288));
    LocalMux I__10661 (
            .O(N__53329),
            .I(N__53288));
    LocalMux I__10660 (
            .O(N__53326),
            .I(N__53288));
    LocalMux I__10659 (
            .O(N__53323),
            .I(N__53288));
    InMux I__10658 (
            .O(N__53320),
            .I(N__53285));
    Span4Mux_v I__10657 (
            .O(N__53317),
            .I(N__53281));
    InMux I__10656 (
            .O(N__53316),
            .I(N__53278));
    InMux I__10655 (
            .O(N__53313),
            .I(N__53275));
    Span4Mux_h I__10654 (
            .O(N__53306),
            .I(N__53262));
    LocalMux I__10653 (
            .O(N__53303),
            .I(N__53262));
    LocalMux I__10652 (
            .O(N__53300),
            .I(N__53262));
    LocalMux I__10651 (
            .O(N__53297),
            .I(N__53262));
    Span4Mux_v I__10650 (
            .O(N__53288),
            .I(N__53262));
    LocalMux I__10649 (
            .O(N__53285),
            .I(N__53262));
    CascadeMux I__10648 (
            .O(N__53284),
            .I(N__53259));
    Span4Mux_h I__10647 (
            .O(N__53281),
            .I(N__53254));
    LocalMux I__10646 (
            .O(N__53278),
            .I(N__53254));
    LocalMux I__10645 (
            .O(N__53275),
            .I(N__53251));
    Span4Mux_v I__10644 (
            .O(N__53262),
            .I(N__53248));
    InMux I__10643 (
            .O(N__53259),
            .I(N__53245));
    Span4Mux_v I__10642 (
            .O(N__53254),
            .I(N__53242));
    Span4Mux_v I__10641 (
            .O(N__53251),
            .I(N__53239));
    Sp12to4 I__10640 (
            .O(N__53248),
            .I(N__53234));
    LocalMux I__10639 (
            .O(N__53245),
            .I(N__53234));
    Odrv4 I__10638 (
            .O(N__53242),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n123 ));
    Odrv4 I__10637 (
            .O(N__53239),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n123 ));
    Odrv12 I__10636 (
            .O(N__53234),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n123 ));
    InMux I__10635 (
            .O(N__53227),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17742 ));
    InMux I__10634 (
            .O(N__53224),
            .I(N__53221));
    LocalMux I__10633 (
            .O(N__53221),
            .I(N__53218));
    Odrv12 I__10632 (
            .O(N__53218),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511 ));
    CascadeMux I__10631 (
            .O(N__53215),
            .I(N__53212));
    InMux I__10630 (
            .O(N__53212),
            .I(N__53207));
    CascadeMux I__10629 (
            .O(N__53211),
            .I(N__53203));
    CascadeMux I__10628 (
            .O(N__53210),
            .I(N__53191));
    LocalMux I__10627 (
            .O(N__53207),
            .I(N__53186));
    InMux I__10626 (
            .O(N__53206),
            .I(N__53183));
    InMux I__10625 (
            .O(N__53203),
            .I(N__53180));
    CascadeMux I__10624 (
            .O(N__53202),
            .I(N__53177));
    CascadeMux I__10623 (
            .O(N__53201),
            .I(N__53174));
    CascadeMux I__10622 (
            .O(N__53200),
            .I(N__53171));
    CascadeMux I__10621 (
            .O(N__53199),
            .I(N__53166));
    CascadeMux I__10620 (
            .O(N__53198),
            .I(N__53162));
    CascadeMux I__10619 (
            .O(N__53197),
            .I(N__53158));
    CascadeMux I__10618 (
            .O(N__53196),
            .I(N__53155));
    CascadeMux I__10617 (
            .O(N__53195),
            .I(N__53151));
    CascadeMux I__10616 (
            .O(N__53194),
            .I(N__53148));
    InMux I__10615 (
            .O(N__53191),
            .I(N__53144));
    CascadeMux I__10614 (
            .O(N__53190),
            .I(N__53141));
    CascadeMux I__10613 (
            .O(N__53189),
            .I(N__53137));
    Span4Mux_h I__10612 (
            .O(N__53186),
            .I(N__53131));
    LocalMux I__10611 (
            .O(N__53183),
            .I(N__53131));
    LocalMux I__10610 (
            .O(N__53180),
            .I(N__53127));
    InMux I__10609 (
            .O(N__53177),
            .I(N__53124));
    InMux I__10608 (
            .O(N__53174),
            .I(N__53121));
    InMux I__10607 (
            .O(N__53171),
            .I(N__53116));
    InMux I__10606 (
            .O(N__53170),
            .I(N__53116));
    InMux I__10605 (
            .O(N__53169),
            .I(N__53103));
    InMux I__10604 (
            .O(N__53166),
            .I(N__53103));
    InMux I__10603 (
            .O(N__53165),
            .I(N__53103));
    InMux I__10602 (
            .O(N__53162),
            .I(N__53103));
    InMux I__10601 (
            .O(N__53161),
            .I(N__53103));
    InMux I__10600 (
            .O(N__53158),
            .I(N__53103));
    InMux I__10599 (
            .O(N__53155),
            .I(N__53100));
    InMux I__10598 (
            .O(N__53154),
            .I(N__53093));
    InMux I__10597 (
            .O(N__53151),
            .I(N__53093));
    InMux I__10596 (
            .O(N__53148),
            .I(N__53093));
    InMux I__10595 (
            .O(N__53147),
            .I(N__53090));
    LocalMux I__10594 (
            .O(N__53144),
            .I(N__53085));
    InMux I__10593 (
            .O(N__53141),
            .I(N__53082));
    CascadeMux I__10592 (
            .O(N__53140),
            .I(N__53079));
    InMux I__10591 (
            .O(N__53137),
            .I(N__53076));
    CascadeMux I__10590 (
            .O(N__53136),
            .I(N__53072));
    Span4Mux_v I__10589 (
            .O(N__53131),
            .I(N__53069));
    InMux I__10588 (
            .O(N__53130),
            .I(N__53066));
    Span4Mux_h I__10587 (
            .O(N__53127),
            .I(N__53059));
    LocalMux I__10586 (
            .O(N__53124),
            .I(N__53059));
    LocalMux I__10585 (
            .O(N__53121),
            .I(N__53059));
    LocalMux I__10584 (
            .O(N__53116),
            .I(N__53048));
    LocalMux I__10583 (
            .O(N__53103),
            .I(N__53048));
    LocalMux I__10582 (
            .O(N__53100),
            .I(N__53048));
    LocalMux I__10581 (
            .O(N__53093),
            .I(N__53048));
    LocalMux I__10580 (
            .O(N__53090),
            .I(N__53048));
    InMux I__10579 (
            .O(N__53089),
            .I(N__53045));
    CascadeMux I__10578 (
            .O(N__53088),
            .I(N__53042));
    Span4Mux_v I__10577 (
            .O(N__53085),
            .I(N__53037));
    LocalMux I__10576 (
            .O(N__53082),
            .I(N__53037));
    InMux I__10575 (
            .O(N__53079),
            .I(N__53034));
    LocalMux I__10574 (
            .O(N__53076),
            .I(N__53031));
    CascadeMux I__10573 (
            .O(N__53075),
            .I(N__53028));
    InMux I__10572 (
            .O(N__53072),
            .I(N__53025));
    Span4Mux_h I__10571 (
            .O(N__53069),
            .I(N__53020));
    LocalMux I__10570 (
            .O(N__53066),
            .I(N__53020));
    Span4Mux_v I__10569 (
            .O(N__53059),
            .I(N__53013));
    Span4Mux_v I__10568 (
            .O(N__53048),
            .I(N__53013));
    LocalMux I__10567 (
            .O(N__53045),
            .I(N__53013));
    InMux I__10566 (
            .O(N__53042),
            .I(N__53010));
    Span4Mux_h I__10565 (
            .O(N__53037),
            .I(N__53005));
    LocalMux I__10564 (
            .O(N__53034),
            .I(N__53005));
    Span4Mux_h I__10563 (
            .O(N__53031),
            .I(N__53002));
    InMux I__10562 (
            .O(N__53028),
            .I(N__52999));
    LocalMux I__10561 (
            .O(N__53025),
            .I(N__52996));
    Span4Mux_v I__10560 (
            .O(N__53020),
            .I(N__52989));
    Span4Mux_v I__10559 (
            .O(N__53013),
            .I(N__52989));
    LocalMux I__10558 (
            .O(N__53010),
            .I(N__52989));
    Span4Mux_v I__10557 (
            .O(N__53005),
            .I(N__52986));
    Span4Mux_v I__10556 (
            .O(N__53002),
            .I(N__52981));
    LocalMux I__10555 (
            .O(N__52999),
            .I(N__52981));
    Span12Mux_h I__10554 (
            .O(N__52996),
            .I(N__52978));
    Span4Mux_h I__10553 (
            .O(N__52989),
            .I(N__52975));
    Span4Mux_v I__10552 (
            .O(N__52986),
            .I(N__52970));
    Span4Mux_h I__10551 (
            .O(N__52981),
            .I(N__52970));
    Odrv12 I__10550 (
            .O(N__52978),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n126 ));
    Odrv4 I__10549 (
            .O(N__52975),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n126 ));
    Odrv4 I__10548 (
            .O(N__52970),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n126 ));
    InMux I__10547 (
            .O(N__52963),
            .I(bfn_21_18_0_));
    CascadeMux I__10546 (
            .O(N__52960),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_ ));
    CascadeMux I__10545 (
            .O(N__52957),
            .I(N__52954));
    InMux I__10544 (
            .O(N__52954),
            .I(N__52951));
    LocalMux I__10543 (
            .O(N__52951),
            .I(N__52948));
    Span4Mux_v I__10542 (
            .O(N__52948),
            .I(N__52945));
    Odrv4 I__10541 (
            .O(N__52945),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20604 ));
    CascadeMux I__10540 (
            .O(N__52942),
            .I(N__52939));
    InMux I__10539 (
            .O(N__52939),
            .I(N__52936));
    LocalMux I__10538 (
            .O(N__52936),
            .I(N__52933));
    Span4Mux_v I__10537 (
            .O(N__52933),
            .I(N__52930));
    Sp12to4 I__10536 (
            .O(N__52930),
            .I(N__52925));
    InMux I__10535 (
            .O(N__52929),
            .I(N__52922));
    InMux I__10534 (
            .O(N__52928),
            .I(N__52919));
    Span12Mux_h I__10533 (
            .O(N__52925),
            .I(N__52912));
    LocalMux I__10532 (
            .O(N__52922),
            .I(N__52912));
    LocalMux I__10531 (
            .O(N__52919),
            .I(N__52912));
    Odrv12 I__10530 (
            .O(N__52912),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25 ));
    InMux I__10529 (
            .O(N__52909),
            .I(N__52906));
    LocalMux I__10528 (
            .O(N__52906),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20588 ));
    InMux I__10527 (
            .O(N__52903),
            .I(N__52900));
    LocalMux I__10526 (
            .O(N__52900),
            .I(N__52897));
    Span4Mux_h I__10525 (
            .O(N__52897),
            .I(N__52894));
    Odrv4 I__10524 (
            .O(N__52894),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896 ));
    CascadeMux I__10523 (
            .O(N__52891),
            .I(\foc.Out_31__N_333_cascade_ ));
    InMux I__10522 (
            .O(N__52888),
            .I(N__52885));
    LocalMux I__10521 (
            .O(N__52885),
            .I(N__52882));
    Span4Mux_h I__10520 (
            .O(N__52882),
            .I(N__52879));
    Odrv4 I__10519 (
            .O(N__52879),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920 ));
    InMux I__10518 (
            .O(N__52876),
            .I(N__52867));
    InMux I__10517 (
            .O(N__52875),
            .I(N__52867));
    InMux I__10516 (
            .O(N__52874),
            .I(N__52867));
    LocalMux I__10515 (
            .O(N__52867),
            .I(N__52864));
    Span12Mux_v I__10514 (
            .O(N__52864),
            .I(N__52861));
    Odrv12 I__10513 (
            .O(N__52861),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30 ));
    CascadeMux I__10512 (
            .O(N__52858),
            .I(N__52854));
    CascadeMux I__10511 (
            .O(N__52857),
            .I(N__52851));
    InMux I__10510 (
            .O(N__52854),
            .I(N__52846));
    InMux I__10509 (
            .O(N__52851),
            .I(N__52846));
    LocalMux I__10508 (
            .O(N__52846),
            .I(N__52843));
    Span4Mux_v I__10507 (
            .O(N__52843),
            .I(N__52839));
    InMux I__10506 (
            .O(N__52842),
            .I(N__52836));
    Sp12to4 I__10505 (
            .O(N__52839),
            .I(N__52831));
    LocalMux I__10504 (
            .O(N__52836),
            .I(N__52831));
    Span12Mux_h I__10503 (
            .O(N__52831),
            .I(N__52828));
    Odrv12 I__10502 (
            .O(N__52828),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29 ));
    InMux I__10501 (
            .O(N__52825),
            .I(N__52819));
    InMux I__10500 (
            .O(N__52824),
            .I(N__52819));
    LocalMux I__10499 (
            .O(N__52819),
            .I(N__52816));
    Span4Mux_h I__10498 (
            .O(N__52816),
            .I(N__52813));
    Span4Mux_v I__10497 (
            .O(N__52813),
            .I(N__52810));
    Span4Mux_v I__10496 (
            .O(N__52810),
            .I(N__52807));
    Odrv4 I__10495 (
            .O(N__52807),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31 ));
    CascadeMux I__10494 (
            .O(N__52804),
            .I(\foc.Out_31__N_332_cascade_ ));
    InMux I__10493 (
            .O(N__52801),
            .I(N__52798));
    LocalMux I__10492 (
            .O(N__52798),
            .I(\foc.qVoltage_9 ));
    InMux I__10491 (
            .O(N__52795),
            .I(N__52789));
    InMux I__10490 (
            .O(N__52794),
            .I(N__52789));
    LocalMux I__10489 (
            .O(N__52789),
            .I(N__52786));
    Span4Mux_h I__10488 (
            .O(N__52786),
            .I(N__52782));
    InMux I__10487 (
            .O(N__52785),
            .I(N__52779));
    Span4Mux_v I__10486 (
            .O(N__52782),
            .I(N__52776));
    LocalMux I__10485 (
            .O(N__52779),
            .I(N__52773));
    Sp12to4 I__10484 (
            .O(N__52776),
            .I(N__52767));
    Span12Mux_h I__10483 (
            .O(N__52773),
            .I(N__52767));
    InMux I__10482 (
            .O(N__52772),
            .I(N__52764));
    Odrv12 I__10481 (
            .O(N__52767),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18 ));
    LocalMux I__10480 (
            .O(N__52764),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18 ));
    CascadeMux I__10479 (
            .O(N__52759),
            .I(\foc.qVoltage_14_cascade_ ));
    InMux I__10478 (
            .O(N__52756),
            .I(N__52750));
    InMux I__10477 (
            .O(N__52755),
            .I(N__52750));
    LocalMux I__10476 (
            .O(N__52750),
            .I(N__52747));
    Span4Mux_h I__10475 (
            .O(N__52747),
            .I(N__52742));
    InMux I__10474 (
            .O(N__52746),
            .I(N__52739));
    InMux I__10473 (
            .O(N__52745),
            .I(N__52736));
    Sp12to4 I__10472 (
            .O(N__52742),
            .I(N__52729));
    LocalMux I__10471 (
            .O(N__52739),
            .I(N__52729));
    LocalMux I__10470 (
            .O(N__52736),
            .I(N__52729));
    Odrv12 I__10469 (
            .O(N__52729),
            .I(\foc.preSatVoltage_23 ));
    InMux I__10468 (
            .O(N__52726),
            .I(N__52723));
    LocalMux I__10467 (
            .O(N__52723),
            .I(N__52719));
    InMux I__10466 (
            .O(N__52722),
            .I(N__52716));
    Span4Mux_v I__10465 (
            .O(N__52719),
            .I(N__52713));
    LocalMux I__10464 (
            .O(N__52716),
            .I(N__52710));
    Span4Mux_h I__10463 (
            .O(N__52713),
            .I(N__52705));
    Span4Mux_v I__10462 (
            .O(N__52710),
            .I(N__52705));
    Span4Mux_h I__10461 (
            .O(N__52705),
            .I(N__52700));
    InMux I__10460 (
            .O(N__52704),
            .I(N__52697));
    InMux I__10459 (
            .O(N__52703),
            .I(N__52694));
    Sp12to4 I__10458 (
            .O(N__52700),
            .I(N__52687));
    LocalMux I__10457 (
            .O(N__52697),
            .I(N__52687));
    LocalMux I__10456 (
            .O(N__52694),
            .I(N__52687));
    Odrv12 I__10455 (
            .O(N__52687),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24 ));
    InMux I__10454 (
            .O(N__52684),
            .I(N__52681));
    LocalMux I__10453 (
            .O(N__52681),
            .I(\foc.qVoltage_15 ));
    CascadeMux I__10452 (
            .O(N__52678),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_ ));
    InMux I__10451 (
            .O(N__52675),
            .I(N__52672));
    LocalMux I__10450 (
            .O(N__52672),
            .I(\foc.dVoltage_15 ));
    CascadeMux I__10449 (
            .O(N__52669),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_ ));
    InMux I__10448 (
            .O(N__52666),
            .I(N__52663));
    LocalMux I__10447 (
            .O(N__52663),
            .I(\foc.dVoltage_10 ));
    CascadeMux I__10446 (
            .O(N__52660),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_ ));
    CascadeMux I__10445 (
            .O(N__52657),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_ ));
    CascadeMux I__10444 (
            .O(N__52654),
            .I(\foc.qVoltage_5_cascade_ ));
    InMux I__10443 (
            .O(N__52651),
            .I(N__52645));
    InMux I__10442 (
            .O(N__52650),
            .I(N__52645));
    LocalMux I__10441 (
            .O(N__52645),
            .I(N__52642));
    Span12Mux_v I__10440 (
            .O(N__52642),
            .I(N__52637));
    InMux I__10439 (
            .O(N__52641),
            .I(N__52634));
    InMux I__10438 (
            .O(N__52640),
            .I(N__52631));
    Odrv12 I__10437 (
            .O(N__52637),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14 ));
    LocalMux I__10436 (
            .O(N__52634),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14 ));
    LocalMux I__10435 (
            .O(N__52631),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14 ));
    InMux I__10434 (
            .O(N__52624),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17560 ));
    CascadeMux I__10433 (
            .O(N__52621),
            .I(N__52618));
    InMux I__10432 (
            .O(N__52618),
            .I(N__52615));
    LocalMux I__10431 (
            .O(N__52615),
            .I(N__52612));
    Odrv12 I__10430 (
            .O(N__52612),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441 ));
    InMux I__10429 (
            .O(N__52609),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17561 ));
    InMux I__10428 (
            .O(N__52606),
            .I(N__52603));
    LocalMux I__10427 (
            .O(N__52603),
            .I(N__52600));
    Odrv4 I__10426 (
            .O(N__52600),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376 ));
    InMux I__10425 (
            .O(N__52597),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17562 ));
    CascadeMux I__10424 (
            .O(N__52594),
            .I(N__52591));
    InMux I__10423 (
            .O(N__52591),
            .I(N__52588));
    LocalMux I__10422 (
            .O(N__52588),
            .I(N__52585));
    Odrv4 I__10421 (
            .O(N__52585),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n648 ));
    InMux I__10420 (
            .O(N__52582),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17563 ));
    InMux I__10419 (
            .O(N__52579),
            .I(N__52576));
    LocalMux I__10418 (
            .O(N__52576),
            .I(N__52573));
    Span4Mux_h I__10417 (
            .O(N__52573),
            .I(N__52569));
    InMux I__10416 (
            .O(N__52572),
            .I(N__52566));
    Span4Mux_v I__10415 (
            .O(N__52569),
            .I(N__52561));
    LocalMux I__10414 (
            .O(N__52566),
            .I(N__52561));
    Odrv4 I__10413 (
            .O(N__52561),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n745 ));
    CascadeMux I__10412 (
            .O(N__52558),
            .I(N__52555));
    InMux I__10411 (
            .O(N__52555),
            .I(N__52552));
    LocalMux I__10410 (
            .O(N__52552),
            .I(N__52549));
    Odrv4 I__10409 (
            .O(N__52549),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444 ));
    CascadeMux I__10408 (
            .O(N__52546),
            .I(N__52543));
    InMux I__10407 (
            .O(N__52543),
            .I(N__52540));
    LocalMux I__10406 (
            .O(N__52540),
            .I(N__52537));
    Odrv4 I__10405 (
            .O(N__52537),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409 ));
    InMux I__10404 (
            .O(N__52534),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17564 ));
    InMux I__10403 (
            .O(N__52531),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408 ));
    CascadeMux I__10402 (
            .O(N__52528),
            .I(N__52525));
    InMux I__10401 (
            .O(N__52525),
            .I(N__52522));
    LocalMux I__10400 (
            .O(N__52522),
            .I(N__52519));
    Span4Mux_v I__10399 (
            .O(N__52519),
            .I(N__52516));
    Odrv4 I__10398 (
            .O(N__52516),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO ));
    CascadeMux I__10397 (
            .O(N__52513),
            .I(\foc.dVoltage_2_cascade_ ));
    InMux I__10396 (
            .O(N__52510),
            .I(N__52507));
    LocalMux I__10395 (
            .O(N__52507),
            .I(N__52504));
    Odrv4 I__10394 (
            .O(N__52504),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n109 ));
    InMux I__10393 (
            .O(N__52501),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17552 ));
    CascadeMux I__10392 (
            .O(N__52498),
            .I(N__52495));
    InMux I__10391 (
            .O(N__52495),
            .I(N__52492));
    LocalMux I__10390 (
            .O(N__52492),
            .I(N__52489));
    Odrv12 I__10389 (
            .O(N__52489),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n158 ));
    InMux I__10388 (
            .O(N__52486),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17553 ));
    InMux I__10387 (
            .O(N__52483),
            .I(N__52480));
    LocalMux I__10386 (
            .O(N__52480),
            .I(N__52477));
    Odrv4 I__10385 (
            .O(N__52477),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394 ));
    InMux I__10384 (
            .O(N__52474),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17554 ));
    CascadeMux I__10383 (
            .O(N__52471),
            .I(N__52468));
    InMux I__10382 (
            .O(N__52468),
            .I(N__52465));
    LocalMux I__10381 (
            .O(N__52465),
            .I(N__52462));
    Odrv4 I__10380 (
            .O(N__52462),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392 ));
    InMux I__10379 (
            .O(N__52459),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17555 ));
    InMux I__10378 (
            .O(N__52456),
            .I(N__52453));
    LocalMux I__10377 (
            .O(N__52453),
            .I(N__52450));
    Odrv12 I__10376 (
            .O(N__52450),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390 ));
    InMux I__10375 (
            .O(N__52447),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17556 ));
    CascadeMux I__10374 (
            .O(N__52444),
            .I(N__52441));
    InMux I__10373 (
            .O(N__52441),
            .I(N__52438));
    LocalMux I__10372 (
            .O(N__52438),
            .I(N__52435));
    Odrv4 I__10371 (
            .O(N__52435),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n354 ));
    InMux I__10370 (
            .O(N__52432),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17557 ));
    InMux I__10369 (
            .O(N__52429),
            .I(N__52426));
    LocalMux I__10368 (
            .O(N__52426),
            .I(N__52423));
    Odrv12 I__10367 (
            .O(N__52423),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n403 ));
    InMux I__10366 (
            .O(N__52420),
            .I(bfn_21_12_0_));
    CascadeMux I__10365 (
            .O(N__52417),
            .I(N__52414));
    InMux I__10364 (
            .O(N__52414),
            .I(N__52411));
    LocalMux I__10363 (
            .O(N__52411),
            .I(N__52408));
    Odrv12 I__10362 (
            .O(N__52408),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n452 ));
    InMux I__10361 (
            .O(N__52405),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17559 ));
    InMux I__10360 (
            .O(N__52402),
            .I(N__52399));
    LocalMux I__10359 (
            .O(N__52399),
            .I(N__52396));
    Odrv4 I__10358 (
            .O(N__52396),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481 ));
    InMux I__10357 (
            .O(N__52393),
            .I(N__52390));
    LocalMux I__10356 (
            .O(N__52390),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467 ));
    InMux I__10355 (
            .O(N__52387),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17575 ));
    CascadeMux I__10354 (
            .O(N__52384),
            .I(N__52381));
    InMux I__10353 (
            .O(N__52381),
            .I(N__52378));
    LocalMux I__10352 (
            .O(N__52378),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446 ));
    InMux I__10351 (
            .O(N__52375),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17576 ));
    InMux I__10350 (
            .O(N__52372),
            .I(N__52369));
    LocalMux I__10349 (
            .O(N__52369),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355 ));
    InMux I__10348 (
            .O(N__52366),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17577 ));
    CascadeMux I__10347 (
            .O(N__52363),
            .I(N__52360));
    InMux I__10346 (
            .O(N__52360),
            .I(N__52357));
    LocalMux I__10345 (
            .O(N__52357),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n651 ));
    InMux I__10344 (
            .O(N__52354),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17578 ));
    InMux I__10343 (
            .O(N__52351),
            .I(N__52348));
    LocalMux I__10342 (
            .O(N__52348),
            .I(N__52345));
    Span4Mux_v I__10341 (
            .O(N__52345),
            .I(N__52341));
    InMux I__10340 (
            .O(N__52344),
            .I(N__52338));
    Odrv4 I__10339 (
            .O(N__52341),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n749 ));
    LocalMux I__10338 (
            .O(N__52338),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n749 ));
    CascadeMux I__10337 (
            .O(N__52333),
            .I(N__52330));
    InMux I__10336 (
            .O(N__52330),
            .I(N__52327));
    LocalMux I__10335 (
            .O(N__52327),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n700 ));
    InMux I__10334 (
            .O(N__52324),
            .I(N__52321));
    LocalMux I__10333 (
            .O(N__52321),
            .I(N__52318));
    Span4Mux_v I__10332 (
            .O(N__52318),
            .I(N__52315));
    Odrv4 I__10331 (
            .O(N__52315),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407 ));
    InMux I__10330 (
            .O(N__52312),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17579 ));
    InMux I__10329 (
            .O(N__52309),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406 ));
    CascadeMux I__10328 (
            .O(N__52306),
            .I(N__52303));
    InMux I__10327 (
            .O(N__52303),
            .I(N__52300));
    LocalMux I__10326 (
            .O(N__52300),
            .I(N__52297));
    Span4Mux_v I__10325 (
            .O(N__52297),
            .I(N__52294));
    Odrv4 I__10324 (
            .O(N__52294),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO ));
    CascadeMux I__10323 (
            .O(N__52291),
            .I(N__52288));
    InMux I__10322 (
            .O(N__52288),
            .I(N__52285));
    LocalMux I__10321 (
            .O(N__52285),
            .I(N__52282));
    Odrv4 I__10320 (
            .O(N__52282),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495 ));
    InMux I__10319 (
            .O(N__52279),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17551 ));
    CascadeMux I__10318 (
            .O(N__52276),
            .I(N__52273));
    InMux I__10317 (
            .O(N__52273),
            .I(N__52270));
    LocalMux I__10316 (
            .O(N__52270),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n63 ));
    InMux I__10315 (
            .O(N__52267),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17566 ));
    InMux I__10314 (
            .O(N__52264),
            .I(N__52261));
    LocalMux I__10313 (
            .O(N__52261),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442 ));
    InMux I__10312 (
            .O(N__52258),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17567 ));
    InMux I__10311 (
            .O(N__52255),
            .I(N__52252));
    LocalMux I__10310 (
            .O(N__52252),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395 ));
    InMux I__10309 (
            .O(N__52249),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17568 ));
    InMux I__10308 (
            .O(N__52246),
            .I(N__52243));
    LocalMux I__10307 (
            .O(N__52243),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393 ));
    InMux I__10306 (
            .O(N__52240),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17569 ));
    CascadeMux I__10305 (
            .O(N__52237),
            .I(N__52234));
    InMux I__10304 (
            .O(N__52234),
            .I(N__52231));
    LocalMux I__10303 (
            .O(N__52231),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391 ));
    InMux I__10302 (
            .O(N__52228),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17570 ));
    InMux I__10301 (
            .O(N__52225),
            .I(N__52222));
    LocalMux I__10300 (
            .O(N__52222),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n308 ));
    InMux I__10299 (
            .O(N__52219),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17571 ));
    CascadeMux I__10298 (
            .O(N__52216),
            .I(N__52213));
    InMux I__10297 (
            .O(N__52213),
            .I(N__52210));
    LocalMux I__10296 (
            .O(N__52210),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n357 ));
    InMux I__10295 (
            .O(N__52207),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17572 ));
    InMux I__10294 (
            .O(N__52204),
            .I(N__52201));
    LocalMux I__10293 (
            .O(N__52201),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n406 ));
    InMux I__10292 (
            .O(N__52198),
            .I(bfn_21_10_0_));
    CascadeMux I__10291 (
            .O(N__52195),
            .I(N__52192));
    InMux I__10290 (
            .O(N__52192),
            .I(N__52189));
    LocalMux I__10289 (
            .O(N__52189),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n455 ));
    InMux I__10288 (
            .O(N__52186),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17574 ));
    CascadeMux I__10287 (
            .O(N__52183),
            .I(N__52180));
    InMux I__10286 (
            .O(N__52180),
            .I(N__52177));
    LocalMux I__10285 (
            .O(N__52177),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470 ));
    CascadeMux I__10284 (
            .O(N__52174),
            .I(N__52171));
    InMux I__10283 (
            .O(N__52171),
            .I(N__52168));
    LocalMux I__10282 (
            .O(N__52168),
            .I(N__52165));
    Odrv4 I__10281 (
            .O(N__52165),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447 ));
    InMux I__10280 (
            .O(N__52162),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17604 ));
    InMux I__10279 (
            .O(N__52159),
            .I(N__52156));
    LocalMux I__10278 (
            .O(N__52156),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458 ));
    InMux I__10277 (
            .O(N__52153),
            .I(N__52150));
    LocalMux I__10276 (
            .O(N__52150),
            .I(N__52147));
    Odrv4 I__10275 (
            .O(N__52147),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n556 ));
    InMux I__10274 (
            .O(N__52144),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17605 ));
    CascadeMux I__10273 (
            .O(N__52141),
            .I(N__52138));
    InMux I__10272 (
            .O(N__52138),
            .I(N__52135));
    LocalMux I__10271 (
            .O(N__52135),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n559 ));
    CascadeMux I__10270 (
            .O(N__52132),
            .I(N__52129));
    InMux I__10269 (
            .O(N__52129),
            .I(N__52126));
    LocalMux I__10268 (
            .O(N__52126),
            .I(N__52123));
    Odrv4 I__10267 (
            .O(N__52123),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n605 ));
    InMux I__10266 (
            .O(N__52120),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17606 ));
    InMux I__10265 (
            .O(N__52117),
            .I(N__52114));
    LocalMux I__10264 (
            .O(N__52114),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n608 ));
    InMux I__10263 (
            .O(N__52111),
            .I(N__52108));
    LocalMux I__10262 (
            .O(N__52108),
            .I(N__52105));
    Span4Mux_v I__10261 (
            .O(N__52105),
            .I(N__52102));
    Odrv4 I__10260 (
            .O(N__52102),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n654 ));
    InMux I__10259 (
            .O(N__52099),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17607 ));
    CascadeMux I__10258 (
            .O(N__52096),
            .I(N__52093));
    InMux I__10257 (
            .O(N__52093),
            .I(N__52090));
    LocalMux I__10256 (
            .O(N__52090),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n657 ));
    CascadeMux I__10255 (
            .O(N__52087),
            .I(N__52084));
    InMux I__10254 (
            .O(N__52084),
            .I(N__52081));
    LocalMux I__10253 (
            .O(N__52081),
            .I(N__52078));
    Sp12to4 I__10252 (
            .O(N__52078),
            .I(N__52075));
    Odrv12 I__10251 (
            .O(N__52075),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n703 ));
    InMux I__10250 (
            .O(N__52072),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17608 ));
    InMux I__10249 (
            .O(N__52069),
            .I(N__52066));
    LocalMux I__10248 (
            .O(N__52066),
            .I(N__52063));
    Span4Mux_h I__10247 (
            .O(N__52063),
            .I(N__52059));
    InMux I__10246 (
            .O(N__52062),
            .I(N__52056));
    Odrv4 I__10245 (
            .O(N__52059),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n757 ));
    LocalMux I__10244 (
            .O(N__52056),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n757 ));
    CascadeMux I__10243 (
            .O(N__52051),
            .I(N__52048));
    InMux I__10242 (
            .O(N__52048),
            .I(N__52045));
    LocalMux I__10241 (
            .O(N__52045),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n706 ));
    InMux I__10240 (
            .O(N__52042),
            .I(N__52039));
    LocalMux I__10239 (
            .O(N__52039),
            .I(N__52036));
    Span4Mux_v I__10238 (
            .O(N__52036),
            .I(N__52033));
    Odrv4 I__10237 (
            .O(N__52033),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403 ));
    InMux I__10236 (
            .O(N__52030),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17609 ));
    InMux I__10235 (
            .O(N__52027),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n759 ));
    CascadeMux I__10234 (
            .O(N__52024),
            .I(N__52021));
    InMux I__10233 (
            .O(N__52021),
            .I(N__52018));
    LocalMux I__10232 (
            .O(N__52018),
            .I(N__52015));
    Span4Mux_v I__10231 (
            .O(N__52015),
            .I(N__52012));
    Odrv4 I__10230 (
            .O(N__52012),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO ));
    InMux I__10229 (
            .O(N__52009),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17596 ));
    CascadeMux I__10228 (
            .O(N__52006),
            .I(N__52003));
    InMux I__10227 (
            .O(N__52003),
            .I(N__52000));
    LocalMux I__10226 (
            .O(N__52000),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487 ));
    InMux I__10225 (
            .O(N__51997),
            .I(N__51994));
    LocalMux I__10224 (
            .O(N__51994),
            .I(N__51991));
    Odrv4 I__10223 (
            .O(N__51991),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466 ));
    InMux I__10222 (
            .O(N__51988),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17597 ));
    InMux I__10221 (
            .O(N__51985),
            .I(N__51982));
    LocalMux I__10220 (
            .O(N__51982),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486 ));
    CascadeMux I__10219 (
            .O(N__51979),
            .I(N__51976));
    InMux I__10218 (
            .O(N__51976),
            .I(N__51973));
    LocalMux I__10217 (
            .O(N__51973),
            .I(N__51970));
    Odrv4 I__10216 (
            .O(N__51970),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445 ));
    InMux I__10215 (
            .O(N__51967),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17598 ));
    InMux I__10214 (
            .O(N__51964),
            .I(N__51961));
    LocalMux I__10213 (
            .O(N__51961),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485 ));
    CascadeMux I__10212 (
            .O(N__51958),
            .I(N__51955));
    InMux I__10211 (
            .O(N__51955),
            .I(N__51952));
    LocalMux I__10210 (
            .O(N__51952),
            .I(N__51949));
    Odrv4 I__10209 (
            .O(N__51949),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n262 ));
    InMux I__10208 (
            .O(N__51946),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17599 ));
    InMux I__10207 (
            .O(N__51943),
            .I(N__51940));
    LocalMux I__10206 (
            .O(N__51940),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471 ));
    InMux I__10205 (
            .O(N__51937),
            .I(N__51934));
    LocalMux I__10204 (
            .O(N__51934),
            .I(N__51931));
    Odrv4 I__10203 (
            .O(N__51931),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n311 ));
    InMux I__10202 (
            .O(N__51928),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17600 ));
    InMux I__10201 (
            .O(N__51925),
            .I(N__51922));
    LocalMux I__10200 (
            .O(N__51922),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n314 ));
    CascadeMux I__10199 (
            .O(N__51919),
            .I(N__51916));
    InMux I__10198 (
            .O(N__51916),
            .I(N__51913));
    LocalMux I__10197 (
            .O(N__51913),
            .I(N__51910));
    Odrv4 I__10196 (
            .O(N__51910),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484 ));
    InMux I__10195 (
            .O(N__51907),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17601 ));
    InMux I__10194 (
            .O(N__51904),
            .I(N__51901));
    LocalMux I__10193 (
            .O(N__51901),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n363 ));
    InMux I__10192 (
            .O(N__51898),
            .I(N__51895));
    LocalMux I__10191 (
            .O(N__51895),
            .I(N__51892));
    Odrv4 I__10190 (
            .O(N__51892),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483 ));
    InMux I__10189 (
            .O(N__51889),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17602 ));
    InMux I__10188 (
            .O(N__51886),
            .I(N__51883));
    LocalMux I__10187 (
            .O(N__51883),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482 ));
    InMux I__10186 (
            .O(N__51880),
            .I(N__51877));
    LocalMux I__10185 (
            .O(N__51877),
            .I(N__51874));
    Odrv4 I__10184 (
            .O(N__51874),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468 ));
    InMux I__10183 (
            .O(N__51871),
            .I(bfn_21_8_0_));
    InMux I__10182 (
            .O(N__51868),
            .I(N__51865));
    LocalMux I__10181 (
            .O(N__51865),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n476 ));
    InMux I__10180 (
            .O(N__51862),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18317 ));
    InMux I__10179 (
            .O(N__51859),
            .I(N__51856));
    LocalMux I__10178 (
            .O(N__51856),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n525 ));
    InMux I__10177 (
            .O(N__51853),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18318 ));
    InMux I__10176 (
            .O(N__51850),
            .I(N__51847));
    LocalMux I__10175 (
            .O(N__51847),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n574 ));
    InMux I__10174 (
            .O(N__51844),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18319 ));
    InMux I__10173 (
            .O(N__51841),
            .I(N__51838));
    LocalMux I__10172 (
            .O(N__51838),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n623 ));
    InMux I__10171 (
            .O(N__51835),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18320 ));
    CascadeMux I__10170 (
            .O(N__51832),
            .I(N__51829));
    InMux I__10169 (
            .O(N__51829),
            .I(N__51826));
    LocalMux I__10168 (
            .O(N__51826),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n672 ));
    InMux I__10167 (
            .O(N__51823),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18321 ));
    CascadeMux I__10166 (
            .O(N__51820),
            .I(N__51817));
    InMux I__10165 (
            .O(N__51817),
            .I(N__51814));
    LocalMux I__10164 (
            .O(N__51814),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n721 ));
    InMux I__10163 (
            .O(N__51811),
            .I(N__51808));
    LocalMux I__10162 (
            .O(N__51808),
            .I(N__51805));
    Span4Mux_v I__10161 (
            .O(N__51805),
            .I(N__51802));
    Sp12to4 I__10160 (
            .O(N__51802),
            .I(N__51799));
    Odrv12 I__10159 (
            .O(N__51799),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n778 ));
    InMux I__10158 (
            .O(N__51796),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18322 ));
    InMux I__10157 (
            .O(N__51793),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779 ));
    CascadeMux I__10156 (
            .O(N__51790),
            .I(N__51787));
    InMux I__10155 (
            .O(N__51787),
            .I(N__51784));
    LocalMux I__10154 (
            .O(N__51784),
            .I(N__51781));
    Span4Mux_h I__10153 (
            .O(N__51781),
            .I(N__51778));
    Span4Mux_v I__10152 (
            .O(N__51778),
            .I(N__51775));
    Odrv4 I__10151 (
            .O(N__51775),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO ));
    InMux I__10150 (
            .O(N__51772),
            .I(N__51769));
    LocalMux I__10149 (
            .O(N__51769),
            .I(N__51766));
    Odrv4 I__10148 (
            .O(N__51766),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n66 ));
    CascadeMux I__10147 (
            .O(N__51763),
            .I(N__51760));
    InMux I__10146 (
            .O(N__51760),
            .I(N__51757));
    LocalMux I__10145 (
            .O(N__51757),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489 ));
    CascadeMux I__10144 (
            .O(N__51754),
            .I(N__51751));
    InMux I__10143 (
            .O(N__51751),
            .I(N__51748));
    LocalMux I__10142 (
            .O(N__51748),
            .I(N__51745));
    Odrv4 I__10141 (
            .O(N__51745),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488 ));
    InMux I__10140 (
            .O(N__51742),
            .I(N__51739));
    LocalMux I__10139 (
            .O(N__51739),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n84 ));
    InMux I__10138 (
            .O(N__51736),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18309 ));
    InMux I__10137 (
            .O(N__51733),
            .I(N__51730));
    LocalMux I__10136 (
            .O(N__51730),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n133 ));
    InMux I__10135 (
            .O(N__51727),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18310 ));
    InMux I__10134 (
            .O(N__51724),
            .I(N__51721));
    LocalMux I__10133 (
            .O(N__51721),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n182 ));
    InMux I__10132 (
            .O(N__51718),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18311 ));
    InMux I__10131 (
            .O(N__51715),
            .I(N__51712));
    LocalMux I__10130 (
            .O(N__51712),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n231 ));
    InMux I__10129 (
            .O(N__51709),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18312 ));
    InMux I__10128 (
            .O(N__51706),
            .I(N__51703));
    LocalMux I__10127 (
            .O(N__51703),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n280 ));
    InMux I__10126 (
            .O(N__51700),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18313 ));
    InMux I__10125 (
            .O(N__51697),
            .I(N__51694));
    LocalMux I__10124 (
            .O(N__51694),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n329 ));
    InMux I__10123 (
            .O(N__51691),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18314 ));
    InMux I__10122 (
            .O(N__51688),
            .I(N__51685));
    LocalMux I__10121 (
            .O(N__51685),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n378 ));
    InMux I__10120 (
            .O(N__51682),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18315 ));
    InMux I__10119 (
            .O(N__51679),
            .I(N__51676));
    LocalMux I__10118 (
            .O(N__51676),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n427 ));
    InMux I__10117 (
            .O(N__51673),
            .I(bfn_20_29_0_));
    InMux I__10116 (
            .O(N__51670),
            .I(N__51667));
    LocalMux I__10115 (
            .O(N__51667),
            .I(N__51664));
    Odrv4 I__10114 (
            .O(N__51664),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n455 ));
    InMux I__10113 (
            .O(N__51661),
            .I(bfn_20_26_0_));
    InMux I__10112 (
            .O(N__51658),
            .I(N__51655));
    LocalMux I__10111 (
            .O(N__51655),
            .I(N__51652));
    Odrv4 I__10110 (
            .O(N__51652),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n504 ));
    InMux I__10109 (
            .O(N__51649),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18227 ));
    InMux I__10108 (
            .O(N__51646),
            .I(N__51643));
    LocalMux I__10107 (
            .O(N__51643),
            .I(N__51640));
    Odrv12 I__10106 (
            .O(N__51640),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n553 ));
    InMux I__10105 (
            .O(N__51637),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18228 ));
    CascadeMux I__10104 (
            .O(N__51634),
            .I(N__51631));
    InMux I__10103 (
            .O(N__51631),
            .I(N__51628));
    LocalMux I__10102 (
            .O(N__51628),
            .I(N__51625));
    Odrv4 I__10101 (
            .O(N__51625),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n602 ));
    InMux I__10100 (
            .O(N__51622),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18229 ));
    CascadeMux I__10099 (
            .O(N__51619),
            .I(N__51616));
    InMux I__10098 (
            .O(N__51616),
            .I(N__51613));
    LocalMux I__10097 (
            .O(N__51613),
            .I(N__51610));
    Span4Mux_h I__10096 (
            .O(N__51610),
            .I(N__51607));
    Odrv4 I__10095 (
            .O(N__51607),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n651 ));
    InMux I__10094 (
            .O(N__51604),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18230 ));
    CascadeMux I__10093 (
            .O(N__51601),
            .I(N__51598));
    InMux I__10092 (
            .O(N__51598),
            .I(N__51595));
    LocalMux I__10091 (
            .O(N__51595),
            .I(N__51592));
    Odrv4 I__10090 (
            .O(N__51592),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n700 ));
    InMux I__10089 (
            .O(N__51589),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18231 ));
    InMux I__10088 (
            .O(N__51586),
            .I(N__51583));
    LocalMux I__10087 (
            .O(N__51583),
            .I(N__51580));
    Span4Mux_v I__10086 (
            .O(N__51580),
            .I(N__51577));
    Odrv4 I__10085 (
            .O(N__51577),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n754 ));
    InMux I__10084 (
            .O(N__51574),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18232 ));
    InMux I__10083 (
            .O(N__51571),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755 ));
    CascadeMux I__10082 (
            .O(N__51568),
            .I(N__51565));
    InMux I__10081 (
            .O(N__51565),
            .I(N__51562));
    LocalMux I__10080 (
            .O(N__51562),
            .I(N__51559));
    Span4Mux_v I__10079 (
            .O(N__51559),
            .I(N__51556));
    Odrv4 I__10078 (
            .O(N__51556),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO ));
    CascadeMux I__10077 (
            .O(N__51553),
            .I(N__51550));
    InMux I__10076 (
            .O(N__51550),
            .I(N__51547));
    LocalMux I__10075 (
            .O(N__51547),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n66 ));
    InMux I__10074 (
            .O(N__51544),
            .I(N__51541));
    LocalMux I__10073 (
            .O(N__51541),
            .I(N__51538));
    Odrv4 I__10072 (
            .O(N__51538),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n112 ));
    InMux I__10071 (
            .O(N__51535),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18219 ));
    InMux I__10070 (
            .O(N__51532),
            .I(N__51529));
    LocalMux I__10069 (
            .O(N__51529),
            .I(N__51526));
    Odrv4 I__10068 (
            .O(N__51526),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n161 ));
    InMux I__10067 (
            .O(N__51523),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18220 ));
    InMux I__10066 (
            .O(N__51520),
            .I(N__51517));
    LocalMux I__10065 (
            .O(N__51517),
            .I(N__51514));
    Odrv4 I__10064 (
            .O(N__51514),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n210 ));
    InMux I__10063 (
            .O(N__51511),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18221 ));
    InMux I__10062 (
            .O(N__51508),
            .I(N__51505));
    LocalMux I__10061 (
            .O(N__51505),
            .I(N__51502));
    Odrv4 I__10060 (
            .O(N__51502),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n259 ));
    InMux I__10059 (
            .O(N__51499),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18222 ));
    CascadeMux I__10058 (
            .O(N__51496),
            .I(N__51493));
    InMux I__10057 (
            .O(N__51493),
            .I(N__51490));
    LocalMux I__10056 (
            .O(N__51490),
            .I(N__51487));
    Odrv4 I__10055 (
            .O(N__51487),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n308 ));
    InMux I__10054 (
            .O(N__51484),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18223 ));
    CascadeMux I__10053 (
            .O(N__51481),
            .I(N__51478));
    InMux I__10052 (
            .O(N__51478),
            .I(N__51475));
    LocalMux I__10051 (
            .O(N__51475),
            .I(N__51472));
    Odrv12 I__10050 (
            .O(N__51472),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n357 ));
    InMux I__10049 (
            .O(N__51469),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18224 ));
    InMux I__10048 (
            .O(N__51466),
            .I(N__51463));
    LocalMux I__10047 (
            .O(N__51463),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n406 ));
    InMux I__10046 (
            .O(N__51460),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18225 ));
    InMux I__10045 (
            .O(N__51457),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18210 ));
    InMux I__10044 (
            .O(N__51454),
            .I(N__51451));
    LocalMux I__10043 (
            .O(N__51451),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n452 ));
    InMux I__10042 (
            .O(N__51448),
            .I(bfn_20_24_0_));
    InMux I__10041 (
            .O(N__51445),
            .I(N__51442));
    LocalMux I__10040 (
            .O(N__51442),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n501 ));
    InMux I__10039 (
            .O(N__51439),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18212 ));
    InMux I__10038 (
            .O(N__51436),
            .I(N__51433));
    LocalMux I__10037 (
            .O(N__51433),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n550 ));
    InMux I__10036 (
            .O(N__51430),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18213 ));
    InMux I__10035 (
            .O(N__51427),
            .I(N__51424));
    LocalMux I__10034 (
            .O(N__51424),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n599 ));
    InMux I__10033 (
            .O(N__51421),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18214 ));
    CascadeMux I__10032 (
            .O(N__51418),
            .I(N__51415));
    InMux I__10031 (
            .O(N__51415),
            .I(N__51412));
    LocalMux I__10030 (
            .O(N__51412),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n648 ));
    InMux I__10029 (
            .O(N__51409),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18215 ));
    CascadeMux I__10028 (
            .O(N__51406),
            .I(N__51403));
    InMux I__10027 (
            .O(N__51403),
            .I(N__51400));
    LocalMux I__10026 (
            .O(N__51400),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n697 ));
    InMux I__10025 (
            .O(N__51397),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18216 ));
    InMux I__10024 (
            .O(N__51394),
            .I(N__51391));
    LocalMux I__10023 (
            .O(N__51391),
            .I(N__51388));
    Span4Mux_v I__10022 (
            .O(N__51388),
            .I(N__51385));
    Odrv4 I__10021 (
            .O(N__51385),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n750 ));
    InMux I__10020 (
            .O(N__51382),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18217 ));
    InMux I__10019 (
            .O(N__51379),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751 ));
    CascadeMux I__10018 (
            .O(N__51376),
            .I(N__51373));
    InMux I__10017 (
            .O(N__51373),
            .I(N__51370));
    LocalMux I__10016 (
            .O(N__51370),
            .I(N__51367));
    Span4Mux_v I__10015 (
            .O(N__51367),
            .I(N__51364));
    Odrv4 I__10014 (
            .O(N__51364),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO ));
    CascadeMux I__10013 (
            .O(N__51361),
            .I(N__51358));
    InMux I__10012 (
            .O(N__51358),
            .I(N__51355));
    LocalMux I__10011 (
            .O(N__51355),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n63 ));
    CascadeMux I__10010 (
            .O(N__51352),
            .I(N__51349));
    InMux I__10009 (
            .O(N__51349),
            .I(N__51346));
    LocalMux I__10008 (
            .O(N__51346),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n109 ));
    InMux I__10007 (
            .O(N__51343),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18204 ));
    InMux I__10006 (
            .O(N__51340),
            .I(N__51337));
    LocalMux I__10005 (
            .O(N__51337),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n158 ));
    InMux I__10004 (
            .O(N__51334),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18205 ));
    InMux I__10003 (
            .O(N__51331),
            .I(N__51328));
    LocalMux I__10002 (
            .O(N__51328),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n207 ));
    InMux I__10001 (
            .O(N__51325),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18206 ));
    InMux I__10000 (
            .O(N__51322),
            .I(N__51319));
    LocalMux I__9999 (
            .O(N__51319),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n256 ));
    InMux I__9998 (
            .O(N__51316),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18207 ));
    InMux I__9997 (
            .O(N__51313),
            .I(N__51310));
    LocalMux I__9996 (
            .O(N__51310),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n305 ));
    InMux I__9995 (
            .O(N__51307),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18208 ));
    InMux I__9994 (
            .O(N__51304),
            .I(N__51301));
    LocalMux I__9993 (
            .O(N__51301),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n354 ));
    InMux I__9992 (
            .O(N__51298),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18209 ));
    InMux I__9991 (
            .O(N__51295),
            .I(N__51292));
    LocalMux I__9990 (
            .O(N__51292),
            .I(N__51289));
    Odrv4 I__9989 (
            .O(N__51289),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n403 ));
    CascadeMux I__9988 (
            .O(N__51286),
            .I(Saturate_out1_31__N_267_adj_2418_cascade_));
    CascadeMux I__9987 (
            .O(N__51283),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_ ));
    CascadeMux I__9986 (
            .O(N__51280),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_ ));
    CascadeMux I__9985 (
            .O(N__51277),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_ ));
    InMux I__9984 (
            .O(N__51274),
            .I(N__51271));
    LocalMux I__9983 (
            .O(N__51271),
            .I(N__51268));
    Odrv4 I__9982 (
            .O(N__51268),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20676 ));
    CascadeMux I__9981 (
            .O(N__51265),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_ ));
    CascadeMux I__9980 (
            .O(N__51262),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_ ));
    CascadeMux I__9979 (
            .O(N__51259),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_ ));
    CascadeMux I__9978 (
            .O(N__51256),
            .I(Saturate_out1_31__N_266_adj_2417_cascade_));
    InMux I__9977 (
            .O(N__51253),
            .I(N__51250));
    LocalMux I__9976 (
            .O(N__51250),
            .I(N__51247));
    Odrv4 I__9975 (
            .O(N__51247),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20620 ));
    InMux I__9974 (
            .O(N__51244),
            .I(N__51241));
    LocalMux I__9973 (
            .O(N__51241),
            .I(N__51238));
    Odrv12 I__9972 (
            .O(N__51238),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20608 ));
    InMux I__9971 (
            .O(N__51235),
            .I(N__51232));
    LocalMux I__9970 (
            .O(N__51232),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18 ));
    InMux I__9969 (
            .O(N__51229),
            .I(N__51226));
    LocalMux I__9968 (
            .O(N__51226),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n27 ));
    CascadeMux I__9967 (
            .O(N__51223),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_ ));
    InMux I__9966 (
            .O(N__51220),
            .I(N__51217));
    LocalMux I__9965 (
            .O(N__51217),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20590 ));
    InMux I__9964 (
            .O(N__51214),
            .I(N__51211));
    LocalMux I__9963 (
            .O(N__51211),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20614 ));
    InMux I__9962 (
            .O(N__51208),
            .I(N__51205));
    LocalMux I__9961 (
            .O(N__51205),
            .I(N__51201));
    InMux I__9960 (
            .O(N__51204),
            .I(N__51198));
    Span4Mux_h I__9959 (
            .O(N__51201),
            .I(N__51194));
    LocalMux I__9958 (
            .O(N__51198),
            .I(N__51191));
    CascadeMux I__9957 (
            .O(N__51197),
            .I(N__51187));
    Sp12to4 I__9956 (
            .O(N__51194),
            .I(N__51182));
    Span12Mux_h I__9955 (
            .O(N__51191),
            .I(N__51182));
    InMux I__9954 (
            .O(N__51190),
            .I(N__51179));
    InMux I__9953 (
            .O(N__51187),
            .I(N__51176));
    Odrv12 I__9952 (
            .O(N__51182),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16 ));
    LocalMux I__9951 (
            .O(N__51179),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16 ));
    LocalMux I__9950 (
            .O(N__51176),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16 ));
    CascadeMux I__9949 (
            .O(N__51169),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_ ));
    InMux I__9948 (
            .O(N__51166),
            .I(N__51163));
    LocalMux I__9947 (
            .O(N__51163),
            .I(\foc.qVoltage_7 ));
    InMux I__9946 (
            .O(N__51160),
            .I(N__51153));
    InMux I__9945 (
            .O(N__51159),
            .I(N__51153));
    CascadeMux I__9944 (
            .O(N__51158),
            .I(N__51150));
    LocalMux I__9943 (
            .O(N__51153),
            .I(N__51146));
    InMux I__9942 (
            .O(N__51150),
            .I(N__51143));
    InMux I__9941 (
            .O(N__51149),
            .I(N__51140));
    Span4Mux_v I__9940 (
            .O(N__51146),
            .I(N__51132));
    LocalMux I__9939 (
            .O(N__51143),
            .I(N__51132));
    LocalMux I__9938 (
            .O(N__51140),
            .I(N__51132));
    InMux I__9937 (
            .O(N__51139),
            .I(N__51129));
    Span4Mux_v I__9936 (
            .O(N__51132),
            .I(N__51122));
    LocalMux I__9935 (
            .O(N__51129),
            .I(N__51122));
    InMux I__9934 (
            .O(N__51128),
            .I(N__51119));
    InMux I__9933 (
            .O(N__51127),
            .I(N__51116));
    Span4Mux_v I__9932 (
            .O(N__51122),
            .I(N__51113));
    LocalMux I__9931 (
            .O(N__51119),
            .I(N__51108));
    LocalMux I__9930 (
            .O(N__51116),
            .I(N__51108));
    Span4Mux_h I__9929 (
            .O(N__51113),
            .I(N__51105));
    Span4Mux_v I__9928 (
            .O(N__51108),
            .I(N__51102));
    Odrv4 I__9927 (
            .O(N__51105),
            .I(Error_sub_temp_31));
    Odrv4 I__9926 (
            .O(N__51102),
            .I(Error_sub_temp_31));
    CascadeMux I__9925 (
            .O(N__51097),
            .I(N__51094));
    InMux I__9924 (
            .O(N__51094),
            .I(N__51090));
    InMux I__9923 (
            .O(N__51093),
            .I(N__51087));
    LocalMux I__9922 (
            .O(N__51090),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424 ));
    LocalMux I__9921 (
            .O(N__51087),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424 ));
    InMux I__9920 (
            .O(N__51082),
            .I(N__51079));
    LocalMux I__9919 (
            .O(N__51079),
            .I(N__51075));
    InMux I__9918 (
            .O(N__51078),
            .I(N__51072));
    Span4Mux_v I__9917 (
            .O(N__51075),
            .I(N__51069));
    LocalMux I__9916 (
            .O(N__51072),
            .I(N__51066));
    Odrv4 I__9915 (
            .O(N__51069),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17 ));
    Odrv12 I__9914 (
            .O(N__51066),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17 ));
    InMux I__9913 (
            .O(N__51061),
            .I(N__51058));
    LocalMux I__9912 (
            .O(N__51058),
            .I(\foc.qVoltage_3 ));
    InMux I__9911 (
            .O(N__51055),
            .I(N__51049));
    InMux I__9910 (
            .O(N__51054),
            .I(N__51049));
    LocalMux I__9909 (
            .O(N__51049),
            .I(N__51046));
    Span4Mux_h I__9908 (
            .O(N__51046),
            .I(N__51043));
    Span4Mux_v I__9907 (
            .O(N__51043),
            .I(N__51038));
    InMux I__9906 (
            .O(N__51042),
            .I(N__51035));
    InMux I__9905 (
            .O(N__51041),
            .I(N__51032));
    Odrv4 I__9904 (
            .O(N__51038),
            .I(\foc.preSatVoltage_13 ));
    LocalMux I__9903 (
            .O(N__51035),
            .I(\foc.preSatVoltage_13 ));
    LocalMux I__9902 (
            .O(N__51032),
            .I(\foc.preSatVoltage_13 ));
    CascadeMux I__9901 (
            .O(N__51025),
            .I(\foc.qVoltage_4_cascade_ ));
    InMux I__9900 (
            .O(N__51022),
            .I(N__51018));
    InMux I__9899 (
            .O(N__51021),
            .I(N__51015));
    LocalMux I__9898 (
            .O(N__51018),
            .I(N__51010));
    LocalMux I__9897 (
            .O(N__51015),
            .I(N__51010));
    Span4Mux_v I__9896 (
            .O(N__51010),
            .I(N__51005));
    CascadeMux I__9895 (
            .O(N__51009),
            .I(N__51002));
    CascadeMux I__9894 (
            .O(N__51008),
            .I(N__50999));
    Span4Mux_v I__9893 (
            .O(N__51005),
            .I(N__50996));
    InMux I__9892 (
            .O(N__51002),
            .I(N__50993));
    InMux I__9891 (
            .O(N__50999),
            .I(N__50990));
    Odrv4 I__9890 (
            .O(N__50996),
            .I(\foc.preSatVoltage_12 ));
    LocalMux I__9889 (
            .O(N__50993),
            .I(\foc.preSatVoltage_12 ));
    LocalMux I__9888 (
            .O(N__50990),
            .I(\foc.preSatVoltage_12 ));
    InMux I__9887 (
            .O(N__50983),
            .I(N__50980));
    LocalMux I__9886 (
            .O(N__50980),
            .I(N__50977));
    Span4Mux_h I__9885 (
            .O(N__50977),
            .I(N__50972));
    InMux I__9884 (
            .O(N__50976),
            .I(N__50967));
    InMux I__9883 (
            .O(N__50975),
            .I(N__50967));
    Sp12to4 I__9882 (
            .O(N__50972),
            .I(N__50962));
    LocalMux I__9881 (
            .O(N__50967),
            .I(N__50962));
    Odrv12 I__9880 (
            .O(N__50962),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26 ));
    CascadeMux I__9879 (
            .O(N__50959),
            .I(N__50956));
    InMux I__9878 (
            .O(N__50956),
            .I(N__50953));
    LocalMux I__9877 (
            .O(N__50953),
            .I(N__50950));
    Span4Mux_h I__9876 (
            .O(N__50950),
            .I(N__50945));
    InMux I__9875 (
            .O(N__50949),
            .I(N__50940));
    InMux I__9874 (
            .O(N__50948),
            .I(N__50940));
    Sp12to4 I__9873 (
            .O(N__50945),
            .I(N__50935));
    LocalMux I__9872 (
            .O(N__50940),
            .I(N__50935));
    Odrv12 I__9871 (
            .O(N__50935),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28 ));
    InMux I__9870 (
            .O(N__50932),
            .I(N__50926));
    InMux I__9869 (
            .O(N__50931),
            .I(N__50926));
    LocalMux I__9868 (
            .O(N__50926),
            .I(N__50923));
    Span4Mux_h I__9867 (
            .O(N__50923),
            .I(N__50919));
    InMux I__9866 (
            .O(N__50922),
            .I(N__50916));
    Span4Mux_v I__9865 (
            .O(N__50919),
            .I(N__50912));
    LocalMux I__9864 (
            .O(N__50916),
            .I(N__50909));
    InMux I__9863 (
            .O(N__50915),
            .I(N__50906));
    Odrv4 I__9862 (
            .O(N__50912),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17 ));
    Odrv4 I__9861 (
            .O(N__50909),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17 ));
    LocalMux I__9860 (
            .O(N__50906),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17 ));
    CascadeMux I__9859 (
            .O(N__50899),
            .I(\foc.qVoltage_8_cascade_ ));
    InMux I__9858 (
            .O(N__50896),
            .I(N__50893));
    LocalMux I__9857 (
            .O(N__50893),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n8265 ));
    InMux I__9856 (
            .O(N__50890),
            .I(N__50887));
    LocalMux I__9855 (
            .O(N__50887),
            .I(N__50884));
    Odrv4 I__9854 (
            .O(N__50884),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19884 ));
    InMux I__9853 (
            .O(N__50881),
            .I(N__50878));
    LocalMux I__9852 (
            .O(N__50878),
            .I(N__50874));
    CascadeMux I__9851 (
            .O(N__50877),
            .I(N__50870));
    Span4Mux_h I__9850 (
            .O(N__50874),
            .I(N__50867));
    InMux I__9849 (
            .O(N__50873),
            .I(N__50862));
    InMux I__9848 (
            .O(N__50870),
            .I(N__50862));
    Span4Mux_v I__9847 (
            .O(N__50867),
            .I(N__50859));
    LocalMux I__9846 (
            .O(N__50862),
            .I(N__50856));
    Odrv4 I__9845 (
            .O(N__50859),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27 ));
    Odrv12 I__9844 (
            .O(N__50856),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27 ));
    CascadeMux I__9843 (
            .O(N__50851),
            .I(N__50848));
    InMux I__9842 (
            .O(N__50848),
            .I(N__50845));
    LocalMux I__9841 (
            .O(N__50845),
            .I(N__50842));
    Span4Mux_v I__9840 (
            .O(N__50842),
            .I(N__50839));
    Span4Mux_v I__9839 (
            .O(N__50839),
            .I(N__50836));
    Span4Mux_v I__9838 (
            .O(N__50836),
            .I(N__50833));
    Odrv4 I__9837 (
            .O(N__50833),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO ));
    InMux I__9836 (
            .O(N__50830),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17516 ));
    InMux I__9835 (
            .O(N__50827),
            .I(N__50824));
    LocalMux I__9834 (
            .O(N__50824),
            .I(N__50821));
    Span4Mux_v I__9833 (
            .O(N__50821),
            .I(N__50818));
    Span4Mux_v I__9832 (
            .O(N__50818),
            .I(N__50815));
    Odrv4 I__9831 (
            .O(N__50815),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348 ));
    CascadeMux I__9830 (
            .O(N__50812),
            .I(N__50809));
    InMux I__9829 (
            .O(N__50809),
            .I(N__50806));
    LocalMux I__9828 (
            .O(N__50806),
            .I(N__50803));
    Span12Mux_h I__9827 (
            .O(N__50803),
            .I(N__50800));
    Odrv12 I__9826 (
            .O(N__50800),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO ));
    InMux I__9825 (
            .O(N__50797),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17517 ));
    InMux I__9824 (
            .O(N__50794),
            .I(N__50791));
    LocalMux I__9823 (
            .O(N__50791),
            .I(N__50788));
    Span4Mux_v I__9822 (
            .O(N__50788),
            .I(N__50785));
    Odrv4 I__9821 (
            .O(N__50785),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n790 ));
    CascadeMux I__9820 (
            .O(N__50782),
            .I(N__50779));
    InMux I__9819 (
            .O(N__50779),
            .I(N__50776));
    LocalMux I__9818 (
            .O(N__50776),
            .I(N__50773));
    Span4Mux_v I__9817 (
            .O(N__50773),
            .I(N__50770));
    Span4Mux_v I__9816 (
            .O(N__50770),
            .I(N__50767));
    Odrv4 I__9815 (
            .O(N__50767),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO ));
    InMux I__9814 (
            .O(N__50764),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17518 ));
    InMux I__9813 (
            .O(N__50761),
            .I(N__50758));
    LocalMux I__9812 (
            .O(N__50758),
            .I(N__50755));
    Odrv4 I__9811 (
            .O(N__50755),
            .I(n794_adj_2420));
    CascadeMux I__9810 (
            .O(N__50752),
            .I(N__50749));
    InMux I__9809 (
            .O(N__50749),
            .I(N__50746));
    LocalMux I__9808 (
            .O(N__50746),
            .I(N__50743));
    Span4Mux_v I__9807 (
            .O(N__50743),
            .I(N__50740));
    Odrv4 I__9806 (
            .O(N__50740),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n791 ));
    InMux I__9805 (
            .O(N__50737),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17519 ));
    InMux I__9804 (
            .O(N__50734),
            .I(N__50731));
    LocalMux I__9803 (
            .O(N__50731),
            .I(N__50727));
    InMux I__9802 (
            .O(N__50730),
            .I(N__50724));
    Span4Mux_v I__9801 (
            .O(N__50727),
            .I(N__50719));
    LocalMux I__9800 (
            .O(N__50724),
            .I(N__50719));
    Odrv4 I__9799 (
            .O(N__50719),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n796 ));
    InMux I__9798 (
            .O(N__50716),
            .I(bfn_20_16_0_));
    CascadeMux I__9797 (
            .O(N__50713),
            .I(N__50709));
    InMux I__9796 (
            .O(N__50712),
            .I(N__50703));
    InMux I__9795 (
            .O(N__50709),
            .I(N__50703));
    CascadeMux I__9794 (
            .O(N__50708),
            .I(N__50700));
    LocalMux I__9793 (
            .O(N__50703),
            .I(N__50697));
    InMux I__9792 (
            .O(N__50700),
            .I(N__50694));
    Span4Mux_h I__9791 (
            .O(N__50697),
            .I(N__50690));
    LocalMux I__9790 (
            .O(N__50694),
            .I(N__50687));
    InMux I__9789 (
            .O(N__50693),
            .I(N__50684));
    Span4Mux_v I__9788 (
            .O(N__50690),
            .I(N__50681));
    Span4Mux_h I__9787 (
            .O(N__50687),
            .I(N__50676));
    LocalMux I__9786 (
            .O(N__50684),
            .I(N__50676));
    Odrv4 I__9785 (
            .O(N__50681),
            .I(\foc.preSatVoltage_19 ));
    Odrv4 I__9784 (
            .O(N__50676),
            .I(\foc.preSatVoltage_19 ));
    InMux I__9783 (
            .O(N__50671),
            .I(N__50668));
    LocalMux I__9782 (
            .O(N__50668),
            .I(\foc.qVoltage_10 ));
    InMux I__9781 (
            .O(N__50665),
            .I(N__50659));
    InMux I__9780 (
            .O(N__50664),
            .I(N__50659));
    LocalMux I__9779 (
            .O(N__50659),
            .I(N__50656));
    Span4Mux_v I__9778 (
            .O(N__50656),
            .I(N__50651));
    CascadeMux I__9777 (
            .O(N__50655),
            .I(N__50648));
    CascadeMux I__9776 (
            .O(N__50654),
            .I(N__50645));
    Sp12to4 I__9775 (
            .O(N__50651),
            .I(N__50642));
    InMux I__9774 (
            .O(N__50648),
            .I(N__50639));
    InMux I__9773 (
            .O(N__50645),
            .I(N__50636));
    Span12Mux_h I__9772 (
            .O(N__50642),
            .I(N__50629));
    LocalMux I__9771 (
            .O(N__50639),
            .I(N__50629));
    LocalMux I__9770 (
            .O(N__50636),
            .I(N__50629));
    Odrv12 I__9769 (
            .O(N__50629),
            .I(\foc.preSatVoltage_22 ));
    InMux I__9768 (
            .O(N__50626),
            .I(N__50623));
    LocalMux I__9767 (
            .O(N__50623),
            .I(\foc.qVoltage_13 ));
    InMux I__9766 (
            .O(N__50620),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17508 ));
    InMux I__9765 (
            .O(N__50617),
            .I(N__50614));
    LocalMux I__9764 (
            .O(N__50614),
            .I(N__50611));
    Odrv12 I__9763 (
            .O(N__50611),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405 ));
    InMux I__9762 (
            .O(N__50608),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17509 ));
    CascadeMux I__9761 (
            .O(N__50605),
            .I(N__50602));
    InMux I__9760 (
            .O(N__50602),
            .I(N__50599));
    LocalMux I__9759 (
            .O(N__50599),
            .I(N__50596));
    Odrv12 I__9758 (
            .O(N__50596),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO ));
    InMux I__9757 (
            .O(N__50593),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17510 ));
    InMux I__9756 (
            .O(N__50590),
            .I(N__50587));
    LocalMux I__9755 (
            .O(N__50587),
            .I(N__50584));
    Odrv12 I__9754 (
            .O(N__50584),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402 ));
    InMux I__9753 (
            .O(N__50581),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17511 ));
    InMux I__9752 (
            .O(N__50578),
            .I(N__50575));
    LocalMux I__9751 (
            .O(N__50575),
            .I(N__50572));
    Span4Mux_v I__9750 (
            .O(N__50572),
            .I(N__50569));
    Odrv4 I__9749 (
            .O(N__50569),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385 ));
    CascadeMux I__9748 (
            .O(N__50566),
            .I(N__50563));
    InMux I__9747 (
            .O(N__50563),
            .I(N__50560));
    LocalMux I__9746 (
            .O(N__50560),
            .I(N__50557));
    Odrv12 I__9745 (
            .O(N__50557),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO ));
    InMux I__9744 (
            .O(N__50554),
            .I(bfn_20_15_0_));
    InMux I__9743 (
            .O(N__50551),
            .I(N__50548));
    LocalMux I__9742 (
            .O(N__50548),
            .I(N__50545));
    Span4Mux_v I__9741 (
            .O(N__50545),
            .I(N__50542));
    Span4Mux_v I__9740 (
            .O(N__50542),
            .I(N__50539));
    Odrv4 I__9739 (
            .O(N__50539),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381 ));
    CascadeMux I__9738 (
            .O(N__50536),
            .I(N__50533));
    InMux I__9737 (
            .O(N__50533),
            .I(N__50530));
    LocalMux I__9736 (
            .O(N__50530),
            .I(N__50527));
    Span12Mux_v I__9735 (
            .O(N__50527),
            .I(N__50524));
    Odrv12 I__9734 (
            .O(N__50524),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO ));
    InMux I__9733 (
            .O(N__50521),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17513 ));
    InMux I__9732 (
            .O(N__50518),
            .I(N__50515));
    LocalMux I__9731 (
            .O(N__50515),
            .I(N__50512));
    Span12Mux_v I__9730 (
            .O(N__50512),
            .I(N__50509));
    Odrv12 I__9729 (
            .O(N__50509),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374 ));
    CascadeMux I__9728 (
            .O(N__50506),
            .I(N__50503));
    InMux I__9727 (
            .O(N__50503),
            .I(N__50500));
    LocalMux I__9726 (
            .O(N__50500),
            .I(N__50497));
    Span12Mux_v I__9725 (
            .O(N__50497),
            .I(N__50494));
    Odrv12 I__9724 (
            .O(N__50494),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO ));
    InMux I__9723 (
            .O(N__50491),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17514 ));
    InMux I__9722 (
            .O(N__50488),
            .I(N__50485));
    LocalMux I__9721 (
            .O(N__50485),
            .I(N__50482));
    Span4Mux_h I__9720 (
            .O(N__50482),
            .I(N__50479));
    Span4Mux_v I__9719 (
            .O(N__50479),
            .I(N__50476));
    Span4Mux_v I__9718 (
            .O(N__50476),
            .I(N__50473));
    Odrv4 I__9717 (
            .O(N__50473),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356 ));
    CascadeMux I__9716 (
            .O(N__50470),
            .I(N__50467));
    InMux I__9715 (
            .O(N__50467),
            .I(N__50464));
    LocalMux I__9714 (
            .O(N__50464),
            .I(N__50461));
    Span12Mux_v I__9713 (
            .O(N__50461),
            .I(N__50458));
    Odrv12 I__9712 (
            .O(N__50458),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO ));
    InMux I__9711 (
            .O(N__50455),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17515 ));
    InMux I__9710 (
            .O(N__50452),
            .I(N__50449));
    LocalMux I__9709 (
            .O(N__50449),
            .I(N__50446));
    Span4Mux_v I__9708 (
            .O(N__50446),
            .I(N__50443));
    Span4Mux_v I__9707 (
            .O(N__50443),
            .I(N__50440));
    Span4Mux_v I__9706 (
            .O(N__50440),
            .I(N__50437));
    Odrv4 I__9705 (
            .O(N__50437),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351 ));
    CascadeMux I__9704 (
            .O(N__50434),
            .I(N__50431));
    InMux I__9703 (
            .O(N__50431),
            .I(N__50428));
    LocalMux I__9702 (
            .O(N__50428),
            .I(N__50425));
    Sp12to4 I__9701 (
            .O(N__50425),
            .I(N__50422));
    Span12Mux_s11_v I__9700 (
            .O(N__50422),
            .I(N__50419));
    Odrv12 I__9699 (
            .O(N__50419),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n721 ));
    InMux I__9698 (
            .O(N__50416),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17909 ));
    CascadeMux I__9697 (
            .O(N__50413),
            .I(N__50410));
    InMux I__9696 (
            .O(N__50410),
            .I(N__50407));
    LocalMux I__9695 (
            .O(N__50407),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n724 ));
    InMux I__9694 (
            .O(N__50404),
            .I(N__50401));
    LocalMux I__9693 (
            .O(N__50401),
            .I(N__50398));
    Span4Mux_v I__9692 (
            .O(N__50398),
            .I(N__50395));
    Odrv4 I__9691 (
            .O(N__50395),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n782 ));
    InMux I__9690 (
            .O(N__50392),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17910 ));
    InMux I__9689 (
            .O(N__50389),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n783 ));
    CascadeMux I__9688 (
            .O(N__50386),
            .I(N__50383));
    InMux I__9687 (
            .O(N__50383),
            .I(N__50380));
    LocalMux I__9686 (
            .O(N__50380),
            .I(N__50377));
    Span4Mux_v I__9685 (
            .O(N__50377),
            .I(N__50374));
    Odrv4 I__9684 (
            .O(N__50374),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO ));
    InMux I__9683 (
            .O(N__50371),
            .I(N__50368));
    LocalMux I__9682 (
            .O(N__50368),
            .I(N__50365));
    Span4Mux_v I__9681 (
            .O(N__50365),
            .I(N__50359));
    InMux I__9680 (
            .O(N__50364),
            .I(N__50354));
    InMux I__9679 (
            .O(N__50363),
            .I(N__50354));
    InMux I__9678 (
            .O(N__50362),
            .I(N__50351));
    Span4Mux_h I__9677 (
            .O(N__50359),
            .I(N__50344));
    LocalMux I__9676 (
            .O(N__50354),
            .I(N__50344));
    LocalMux I__9675 (
            .O(N__50351),
            .I(N__50344));
    Span4Mux_v I__9674 (
            .O(N__50344),
            .I(N__50339));
    InMux I__9673 (
            .O(N__50343),
            .I(N__50336));
    InMux I__9672 (
            .O(N__50342),
            .I(N__50333));
    Odrv4 I__9671 (
            .O(N__50339),
            .I(Error_sub_temp_30));
    LocalMux I__9670 (
            .O(N__50336),
            .I(Error_sub_temp_30));
    LocalMux I__9669 (
            .O(N__50333),
            .I(Error_sub_temp_30));
    InMux I__9668 (
            .O(N__50326),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17505 ));
    InMux I__9667 (
            .O(N__50323),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17506 ));
    InMux I__9666 (
            .O(N__50320),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17507 ));
    InMux I__9665 (
            .O(N__50317),
            .I(N__50314));
    LocalMux I__9664 (
            .O(N__50314),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513 ));
    InMux I__9663 (
            .O(N__50311),
            .I(N__50308));
    LocalMux I__9662 (
            .O(N__50308),
            .I(N__50305));
    Span4Mux_v I__9661 (
            .O(N__50305),
            .I(N__50302));
    Odrv4 I__9660 (
            .O(N__50302),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436 ));
    InMux I__9659 (
            .O(N__50299),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17902 ));
    InMux I__9658 (
            .O(N__50296),
            .I(N__50293));
    LocalMux I__9657 (
            .O(N__50293),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n381 ));
    InMux I__9656 (
            .O(N__50290),
            .I(N__50287));
    LocalMux I__9655 (
            .O(N__50287),
            .I(N__50284));
    Odrv4 I__9654 (
            .O(N__50284),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432 ));
    InMux I__9653 (
            .O(N__50281),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17903 ));
    InMux I__9652 (
            .O(N__50278),
            .I(N__50275));
    LocalMux I__9651 (
            .O(N__50275),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n430 ));
    InMux I__9650 (
            .O(N__50272),
            .I(N__50269));
    LocalMux I__9649 (
            .O(N__50269),
            .I(N__50266));
    Span4Mux_v I__9648 (
            .O(N__50266),
            .I(N__50263));
    Odrv4 I__9647 (
            .O(N__50263),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n476 ));
    InMux I__9646 (
            .O(N__50260),
            .I(bfn_20_12_0_));
    InMux I__9645 (
            .O(N__50257),
            .I(N__50254));
    LocalMux I__9644 (
            .O(N__50254),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n479 ));
    InMux I__9643 (
            .O(N__50251),
            .I(N__50248));
    LocalMux I__9642 (
            .O(N__50248),
            .I(N__50245));
    Span4Mux_v I__9641 (
            .O(N__50245),
            .I(N__50242));
    Odrv4 I__9640 (
            .O(N__50242),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n525 ));
    InMux I__9639 (
            .O(N__50239),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17905 ));
    InMux I__9638 (
            .O(N__50236),
            .I(N__50233));
    LocalMux I__9637 (
            .O(N__50233),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n528 ));
    InMux I__9636 (
            .O(N__50230),
            .I(N__50227));
    LocalMux I__9635 (
            .O(N__50227),
            .I(N__50224));
    Span4Mux_h I__9634 (
            .O(N__50224),
            .I(N__50221));
    Odrv4 I__9633 (
            .O(N__50221),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n574 ));
    InMux I__9632 (
            .O(N__50218),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17906 ));
    InMux I__9631 (
            .O(N__50215),
            .I(N__50212));
    LocalMux I__9630 (
            .O(N__50212),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n577 ));
    InMux I__9629 (
            .O(N__50209),
            .I(N__50206));
    LocalMux I__9628 (
            .O(N__50206),
            .I(N__50203));
    Span4Mux_v I__9627 (
            .O(N__50203),
            .I(N__50200));
    Odrv4 I__9626 (
            .O(N__50200),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n623 ));
    InMux I__9625 (
            .O(N__50197),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17907 ));
    InMux I__9624 (
            .O(N__50194),
            .I(N__50191));
    LocalMux I__9623 (
            .O(N__50191),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n626 ));
    CascadeMux I__9622 (
            .O(N__50188),
            .I(N__50185));
    InMux I__9621 (
            .O(N__50185),
            .I(N__50182));
    LocalMux I__9620 (
            .O(N__50182),
            .I(N__50179));
    Span4Mux_h I__9619 (
            .O(N__50179),
            .I(N__50176));
    Odrv4 I__9618 (
            .O(N__50176),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n672 ));
    InMux I__9617 (
            .O(N__50173),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17908 ));
    CascadeMux I__9616 (
            .O(N__50170),
            .I(N__50167));
    InMux I__9615 (
            .O(N__50167),
            .I(N__50164));
    LocalMux I__9614 (
            .O(N__50164),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n675 ));
    InMux I__9613 (
            .O(N__50161),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17593 ));
    InMux I__9612 (
            .O(N__50158),
            .I(N__50155));
    LocalMux I__9611 (
            .O(N__50155),
            .I(N__50151));
    InMux I__9610 (
            .O(N__50154),
            .I(N__50148));
    Span4Mux_v I__9609 (
            .O(N__50151),
            .I(N__50143));
    LocalMux I__9608 (
            .O(N__50148),
            .I(N__50143));
    Span4Mux_h I__9607 (
            .O(N__50143),
            .I(N__50140));
    Odrv4 I__9606 (
            .O(N__50140),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n753 ));
    InMux I__9605 (
            .O(N__50137),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17594 ));
    InMux I__9604 (
            .O(N__50134),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404 ));
    InMux I__9603 (
            .O(N__50131),
            .I(N__50128));
    LocalMux I__9602 (
            .O(N__50128),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n87 ));
    InMux I__9601 (
            .O(N__50125),
            .I(N__50122));
    LocalMux I__9600 (
            .O(N__50122),
            .I(N__50119));
    Span4Mux_v I__9599 (
            .O(N__50119),
            .I(N__50116));
    Odrv4 I__9598 (
            .O(N__50116),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388 ));
    InMux I__9597 (
            .O(N__50113),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17897 ));
    InMux I__9596 (
            .O(N__50110),
            .I(N__50107));
    LocalMux I__9595 (
            .O(N__50107),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n136 ));
    InMux I__9594 (
            .O(N__50104),
            .I(N__50101));
    LocalMux I__9593 (
            .O(N__50101),
            .I(N__50098));
    Span4Mux_h I__9592 (
            .O(N__50098),
            .I(N__50095));
    Odrv4 I__9591 (
            .O(N__50095),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451 ));
    InMux I__9590 (
            .O(N__50092),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17898 ));
    InMux I__9589 (
            .O(N__50089),
            .I(N__50086));
    LocalMux I__9588 (
            .O(N__50086),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n185 ));
    InMux I__9587 (
            .O(N__50083),
            .I(N__50080));
    LocalMux I__9586 (
            .O(N__50080),
            .I(N__50077));
    Span12Mux_h I__9585 (
            .O(N__50077),
            .I(N__50074));
    Odrv12 I__9584 (
            .O(N__50074),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387 ));
    InMux I__9583 (
            .O(N__50071),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17899 ));
    InMux I__9582 (
            .O(N__50068),
            .I(N__50065));
    LocalMux I__9581 (
            .O(N__50065),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n234 ));
    InMux I__9580 (
            .O(N__50062),
            .I(N__50059));
    LocalMux I__9579 (
            .O(N__50059),
            .I(N__50056));
    Span4Mux_h I__9578 (
            .O(N__50056),
            .I(N__50053));
    Odrv4 I__9577 (
            .O(N__50053),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379 ));
    InMux I__9576 (
            .O(N__50050),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17900 ));
    CascadeMux I__9575 (
            .O(N__50047),
            .I(N__50044));
    InMux I__9574 (
            .O(N__50044),
            .I(N__50041));
    LocalMux I__9573 (
            .O(N__50041),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514 ));
    InMux I__9572 (
            .O(N__50038),
            .I(N__50035));
    LocalMux I__9571 (
            .O(N__50035),
            .I(N__50032));
    Span4Mux_h I__9570 (
            .O(N__50032),
            .I(N__50029));
    Odrv4 I__9569 (
            .O(N__50029),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439 ));
    InMux I__9568 (
            .O(N__50026),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17901 ));
    InMux I__9567 (
            .O(N__50023),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17584 ));
    InMux I__9566 (
            .O(N__50020),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17585 ));
    InMux I__9565 (
            .O(N__50017),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17586 ));
    InMux I__9564 (
            .O(N__50014),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17587 ));
    InMux I__9563 (
            .O(N__50011),
            .I(bfn_20_10_0_));
    InMux I__9562 (
            .O(N__50008),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17589 ));
    InMux I__9561 (
            .O(N__50005),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17590 ));
    InMux I__9560 (
            .O(N__50002),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17591 ));
    InMux I__9559 (
            .O(N__49999),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17592 ));
    InMux I__9558 (
            .O(N__49996),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17621 ));
    InMux I__9557 (
            .O(N__49993),
            .I(N__49990));
    LocalMux I__9556 (
            .O(N__49990),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n611 ));
    InMux I__9555 (
            .O(N__49987),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17622 ));
    CascadeMux I__9554 (
            .O(N__49984),
            .I(N__49981));
    InMux I__9553 (
            .O(N__49981),
            .I(N__49978));
    LocalMux I__9552 (
            .O(N__49978),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n660 ));
    InMux I__9551 (
            .O(N__49975),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17623 ));
    InMux I__9550 (
            .O(N__49972),
            .I(N__49969));
    LocalMux I__9549 (
            .O(N__49969),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512 ));
    CascadeMux I__9548 (
            .O(N__49966),
            .I(N__49963));
    InMux I__9547 (
            .O(N__49963),
            .I(N__49960));
    LocalMux I__9546 (
            .O(N__49960),
            .I(N__49957));
    Span4Mux_v I__9545 (
            .O(N__49957),
            .I(N__49953));
    InMux I__9544 (
            .O(N__49956),
            .I(N__49950));
    Odrv4 I__9543 (
            .O(N__49953),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n761 ));
    LocalMux I__9542 (
            .O(N__49950),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n761 ));
    InMux I__9541 (
            .O(N__49945),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17624 ));
    InMux I__9540 (
            .O(N__49942),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386 ));
    InMux I__9539 (
            .O(N__49939),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17581 ));
    InMux I__9538 (
            .O(N__49936),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17582 ));
    InMux I__9537 (
            .O(N__49933),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17583 ));
    InMux I__9536 (
            .O(N__49930),
            .I(N__49927));
    LocalMux I__9535 (
            .O(N__49927),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490 ));
    InMux I__9534 (
            .O(N__49924),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17613 ));
    InMux I__9533 (
            .O(N__49921),
            .I(N__49918));
    LocalMux I__9532 (
            .O(N__49918),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472 ));
    InMux I__9531 (
            .O(N__49915),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17614 ));
    InMux I__9530 (
            .O(N__49912),
            .I(N__49909));
    LocalMux I__9529 (
            .O(N__49909),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n268 ));
    InMux I__9528 (
            .O(N__49906),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17615 ));
    InMux I__9527 (
            .O(N__49903),
            .I(N__49900));
    LocalMux I__9526 (
            .O(N__49900),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n317 ));
    InMux I__9525 (
            .O(N__49897),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17616 ));
    InMux I__9524 (
            .O(N__49894),
            .I(N__49891));
    LocalMux I__9523 (
            .O(N__49891),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n366 ));
    InMux I__9522 (
            .O(N__49888),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17617 ));
    InMux I__9521 (
            .O(N__49885),
            .I(N__49882));
    LocalMux I__9520 (
            .O(N__49882),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449 ));
    InMux I__9519 (
            .O(N__49879),
            .I(bfn_20_8_0_));
    CascadeMux I__9518 (
            .O(N__49876),
            .I(N__49873));
    InMux I__9517 (
            .O(N__49873),
            .I(N__49870));
    LocalMux I__9516 (
            .O(N__49870),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n464 ));
    InMux I__9515 (
            .O(N__49867),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17619 ));
    InMux I__9514 (
            .O(N__49864),
            .I(N__49861));
    LocalMux I__9513 (
            .O(N__49861),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n513 ));
    InMux I__9512 (
            .O(N__49858),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17620 ));
    CascadeMux I__9511 (
            .O(N__49855),
            .I(N__49852));
    InMux I__9510 (
            .O(N__49852),
            .I(N__49849));
    LocalMux I__9509 (
            .O(N__49849),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n562 ));
    InMux I__9508 (
            .O(N__49846),
            .I(N__49843));
    LocalMux I__9507 (
            .O(N__49843),
            .I(N__49840));
    Odrv4 I__9506 (
            .O(N__49840),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n473 ));
    CascadeMux I__9505 (
            .O(N__49837),
            .I(N__49834));
    InMux I__9504 (
            .O(N__49834),
            .I(N__49831));
    LocalMux I__9503 (
            .O(N__49831),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n519 ));
    InMux I__9502 (
            .O(N__49828),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18130 ));
    InMux I__9501 (
            .O(N__49825),
            .I(N__49822));
    LocalMux I__9500 (
            .O(N__49822),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n568 ));
    InMux I__9499 (
            .O(N__49819),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18131 ));
    CascadeMux I__9498 (
            .O(N__49816),
            .I(N__49811));
    InMux I__9497 (
            .O(N__49815),
            .I(N__49808));
    InMux I__9496 (
            .O(N__49814),
            .I(N__49803));
    InMux I__9495 (
            .O(N__49811),
            .I(N__49803));
    LocalMux I__9494 (
            .O(N__49808),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n617 ));
    LocalMux I__9493 (
            .O(N__49803),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n617 ));
    InMux I__9492 (
            .O(N__49798),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18132 ));
    InMux I__9491 (
            .O(N__49795),
            .I(N__49791));
    InMux I__9490 (
            .O(N__49794),
            .I(N__49788));
    LocalMux I__9489 (
            .O(N__49791),
            .I(N__49785));
    LocalMux I__9488 (
            .O(N__49788),
            .I(N__49782));
    Span4Mux_h I__9487 (
            .O(N__49785),
            .I(N__49779));
    Span4Mux_v I__9486 (
            .O(N__49782),
            .I(N__49776));
    Odrv4 I__9485 (
            .O(N__49779),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n773 ));
    Odrv4 I__9484 (
            .O(N__49776),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n773 ));
    CascadeMux I__9483 (
            .O(N__49771),
            .I(N__49767));
    CascadeMux I__9482 (
            .O(N__49770),
            .I(N__49764));
    InMux I__9481 (
            .O(N__49767),
            .I(N__49760));
    InMux I__9480 (
            .O(N__49764),
            .I(N__49755));
    InMux I__9479 (
            .O(N__49763),
            .I(N__49755));
    LocalMux I__9478 (
            .O(N__49760),
            .I(N__49750));
    LocalMux I__9477 (
            .O(N__49755),
            .I(N__49750));
    Odrv4 I__9476 (
            .O(N__49750),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n522 ));
    InMux I__9475 (
            .O(N__49747),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18133 ));
    InMux I__9474 (
            .O(N__49744),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357 ));
    InMux I__9473 (
            .O(N__49741),
            .I(N__49738));
    LocalMux I__9472 (
            .O(N__49738),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508 ));
    InMux I__9471 (
            .O(N__49735),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17611 ));
    CascadeMux I__9470 (
            .O(N__49732),
            .I(N__49729));
    InMux I__9469 (
            .O(N__49729),
            .I(N__49726));
    LocalMux I__9468 (
            .O(N__49726),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504 ));
    InMux I__9467 (
            .O(N__49723),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17612 ));
    CascadeMux I__9466 (
            .O(N__49720),
            .I(N__49717));
    InMux I__9465 (
            .O(N__49717),
            .I(N__49714));
    LocalMux I__9464 (
            .O(N__49714),
            .I(N__49711));
    Odrv12 I__9463 (
            .O(N__49711),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n81 ));
    InMux I__9462 (
            .O(N__49708),
            .I(N__49705));
    LocalMux I__9461 (
            .O(N__49705),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n127 ));
    InMux I__9460 (
            .O(N__49702),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18122 ));
    InMux I__9459 (
            .O(N__49699),
            .I(N__49696));
    LocalMux I__9458 (
            .O(N__49696),
            .I(N__49693));
    Odrv4 I__9457 (
            .O(N__49693),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n130 ));
    CascadeMux I__9456 (
            .O(N__49690),
            .I(N__49687));
    InMux I__9455 (
            .O(N__49687),
            .I(N__49684));
    LocalMux I__9454 (
            .O(N__49684),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n176 ));
    InMux I__9453 (
            .O(N__49681),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18123 ));
    CascadeMux I__9452 (
            .O(N__49678),
            .I(N__49675));
    InMux I__9451 (
            .O(N__49675),
            .I(N__49672));
    LocalMux I__9450 (
            .O(N__49672),
            .I(N__49669));
    Odrv12 I__9449 (
            .O(N__49669),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n179 ));
    InMux I__9448 (
            .O(N__49666),
            .I(N__49663));
    LocalMux I__9447 (
            .O(N__49663),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n225 ));
    InMux I__9446 (
            .O(N__49660),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18124 ));
    InMux I__9445 (
            .O(N__49657),
            .I(N__49654));
    LocalMux I__9444 (
            .O(N__49654),
            .I(N__49651));
    Odrv12 I__9443 (
            .O(N__49651),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n228 ));
    InMux I__9442 (
            .O(N__49648),
            .I(N__49645));
    LocalMux I__9441 (
            .O(N__49645),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n274 ));
    InMux I__9440 (
            .O(N__49642),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18125 ));
    CascadeMux I__9439 (
            .O(N__49639),
            .I(N__49636));
    InMux I__9438 (
            .O(N__49636),
            .I(N__49633));
    LocalMux I__9437 (
            .O(N__49633),
            .I(N__49630));
    Odrv4 I__9436 (
            .O(N__49630),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n277 ));
    InMux I__9435 (
            .O(N__49627),
            .I(N__49624));
    LocalMux I__9434 (
            .O(N__49624),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n323 ));
    InMux I__9433 (
            .O(N__49621),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18126 ));
    CascadeMux I__9432 (
            .O(N__49618),
            .I(N__49615));
    InMux I__9431 (
            .O(N__49615),
            .I(N__49612));
    LocalMux I__9430 (
            .O(N__49612),
            .I(N__49609));
    Odrv12 I__9429 (
            .O(N__49609),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n326 ));
    CascadeMux I__9428 (
            .O(N__49606),
            .I(N__49603));
    InMux I__9427 (
            .O(N__49603),
            .I(N__49600));
    LocalMux I__9426 (
            .O(N__49600),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n372 ));
    InMux I__9425 (
            .O(N__49597),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18127 ));
    InMux I__9424 (
            .O(N__49594),
            .I(N__49591));
    LocalMux I__9423 (
            .O(N__49591),
            .I(N__49588));
    Odrv12 I__9422 (
            .O(N__49588),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n375 ));
    CascadeMux I__9421 (
            .O(N__49585),
            .I(N__49582));
    InMux I__9420 (
            .O(N__49582),
            .I(N__49579));
    LocalMux I__9419 (
            .O(N__49579),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n421 ));
    InMux I__9418 (
            .O(N__49576),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18128 ));
    InMux I__9417 (
            .O(N__49573),
            .I(N__49570));
    LocalMux I__9416 (
            .O(N__49570),
            .I(N__49567));
    Span4Mux_h I__9415 (
            .O(N__49567),
            .I(N__49564));
    Odrv4 I__9414 (
            .O(N__49564),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n424 ));
    InMux I__9413 (
            .O(N__49561),
            .I(N__49558));
    LocalMux I__9412 (
            .O(N__49558),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n470 ));
    InMux I__9411 (
            .O(N__49555),
            .I(bfn_20_6_0_));
    InMux I__9410 (
            .O(N__49552),
            .I(bfn_19_29_0_));
    InMux I__9409 (
            .O(N__49549),
            .I(N__49546));
    LocalMux I__9408 (
            .O(N__49546),
            .I(N__49543));
    Odrv4 I__9407 (
            .O(N__49543),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n479 ));
    InMux I__9406 (
            .O(N__49540),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18332 ));
    InMux I__9405 (
            .O(N__49537),
            .I(N__49534));
    LocalMux I__9404 (
            .O(N__49534),
            .I(N__49531));
    Odrv4 I__9403 (
            .O(N__49531),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n528 ));
    InMux I__9402 (
            .O(N__49528),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18333 ));
    InMux I__9401 (
            .O(N__49525),
            .I(N__49522));
    LocalMux I__9400 (
            .O(N__49522),
            .I(N__49519));
    Odrv12 I__9399 (
            .O(N__49519),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n577 ));
    InMux I__9398 (
            .O(N__49516),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18334 ));
    InMux I__9397 (
            .O(N__49513),
            .I(N__49510));
    LocalMux I__9396 (
            .O(N__49510),
            .I(N__49507));
    Odrv12 I__9395 (
            .O(N__49507),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n626 ));
    InMux I__9394 (
            .O(N__49504),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18335 ));
    CascadeMux I__9393 (
            .O(N__49501),
            .I(N__49498));
    InMux I__9392 (
            .O(N__49498),
            .I(N__49495));
    LocalMux I__9391 (
            .O(N__49495),
            .I(N__49492));
    Span4Mux_v I__9390 (
            .O(N__49492),
            .I(N__49489));
    Odrv4 I__9389 (
            .O(N__49489),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n675 ));
    InMux I__9388 (
            .O(N__49486),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18336 ));
    InMux I__9387 (
            .O(N__49483),
            .I(N__49480));
    LocalMux I__9386 (
            .O(N__49480),
            .I(N__49477));
    Odrv4 I__9385 (
            .O(N__49477),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n724 ));
    InMux I__9384 (
            .O(N__49474),
            .I(N__49471));
    LocalMux I__9383 (
            .O(N__49471),
            .I(N__49468));
    Span12Mux_v I__9382 (
            .O(N__49468),
            .I(N__49465));
    Odrv12 I__9381 (
            .O(N__49465),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n782 ));
    InMux I__9380 (
            .O(N__49462),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18337 ));
    InMux I__9379 (
            .O(N__49459),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783 ));
    CascadeMux I__9378 (
            .O(N__49456),
            .I(N__49453));
    InMux I__9377 (
            .O(N__49453),
            .I(N__49450));
    LocalMux I__9376 (
            .O(N__49450),
            .I(N__49447));
    Span12Mux_v I__9375 (
            .O(N__49447),
            .I(N__49444));
    Odrv12 I__9374 (
            .O(N__49444),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO ));
    CascadeMux I__9373 (
            .O(N__49441),
            .I(N__49438));
    InMux I__9372 (
            .O(N__49438),
            .I(N__49435));
    LocalMux I__9371 (
            .O(N__49435),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n78 ));
    CascadeMux I__9370 (
            .O(N__49432),
            .I(N__49429));
    InMux I__9369 (
            .O(N__49429),
            .I(N__49426));
    LocalMux I__9368 (
            .O(N__49426),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n87 ));
    InMux I__9367 (
            .O(N__49423),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18324 ));
    InMux I__9366 (
            .O(N__49420),
            .I(N__49417));
    LocalMux I__9365 (
            .O(N__49417),
            .I(N__49414));
    Odrv4 I__9364 (
            .O(N__49414),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n136 ));
    InMux I__9363 (
            .O(N__49411),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18325 ));
    CascadeMux I__9362 (
            .O(N__49408),
            .I(N__49405));
    InMux I__9361 (
            .O(N__49405),
            .I(N__49402));
    LocalMux I__9360 (
            .O(N__49402),
            .I(N__49399));
    Odrv4 I__9359 (
            .O(N__49399),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n185 ));
    InMux I__9358 (
            .O(N__49396),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18326 ));
    InMux I__9357 (
            .O(N__49393),
            .I(N__49390));
    LocalMux I__9356 (
            .O(N__49390),
            .I(N__49387));
    Odrv4 I__9355 (
            .O(N__49387),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n234 ));
    InMux I__9354 (
            .O(N__49384),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18327 ));
    InMux I__9353 (
            .O(N__49381),
            .I(N__49378));
    LocalMux I__9352 (
            .O(N__49378),
            .I(N__49375));
    Odrv4 I__9351 (
            .O(N__49375),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n283 ));
    InMux I__9350 (
            .O(N__49372),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18328 ));
    InMux I__9349 (
            .O(N__49369),
            .I(N__49366));
    LocalMux I__9348 (
            .O(N__49366),
            .I(N__49363));
    Odrv4 I__9347 (
            .O(N__49363),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n332 ));
    InMux I__9346 (
            .O(N__49360),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18329 ));
    InMux I__9345 (
            .O(N__49357),
            .I(N__49354));
    LocalMux I__9344 (
            .O(N__49354),
            .I(N__49351));
    Odrv4 I__9343 (
            .O(N__49351),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n381 ));
    InMux I__9342 (
            .O(N__49348),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18330 ));
    InMux I__9341 (
            .O(N__49345),
            .I(N__49342));
    LocalMux I__9340 (
            .O(N__49342),
            .I(N__49339));
    Odrv12 I__9339 (
            .O(N__49339),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n430 ));
    CascadeMux I__9338 (
            .O(N__49336),
            .I(N__49333));
    InMux I__9337 (
            .O(N__49333),
            .I(N__49330));
    LocalMux I__9336 (
            .O(N__49330),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n433 ));
    InMux I__9335 (
            .O(N__49327),
            .I(bfn_19_27_0_));
    InMux I__9334 (
            .O(N__49324),
            .I(N__49321));
    LocalMux I__9333 (
            .O(N__49321),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n482 ));
    InMux I__9332 (
            .O(N__49318),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18347 ));
    CascadeMux I__9331 (
            .O(N__49315),
            .I(N__49312));
    InMux I__9330 (
            .O(N__49312),
            .I(N__49309));
    LocalMux I__9329 (
            .O(N__49309),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n531 ));
    InMux I__9328 (
            .O(N__49306),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18348 ));
    InMux I__9327 (
            .O(N__49303),
            .I(N__49300));
    LocalMux I__9326 (
            .O(N__49300),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n580 ));
    InMux I__9325 (
            .O(N__49297),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18349 ));
    InMux I__9324 (
            .O(N__49294),
            .I(N__49291));
    LocalMux I__9323 (
            .O(N__49291),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n629 ));
    InMux I__9322 (
            .O(N__49288),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18350 ));
    InMux I__9321 (
            .O(N__49285),
            .I(N__49282));
    LocalMux I__9320 (
            .O(N__49282),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n678 ));
    InMux I__9319 (
            .O(N__49279),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18351 ));
    CascadeMux I__9318 (
            .O(N__49276),
            .I(N__49273));
    InMux I__9317 (
            .O(N__49273),
            .I(N__49270));
    LocalMux I__9316 (
            .O(N__49270),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n727 ));
    InMux I__9315 (
            .O(N__49267),
            .I(N__49264));
    LocalMux I__9314 (
            .O(N__49264),
            .I(N__49261));
    Odrv12 I__9313 (
            .O(N__49261),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n786 ));
    InMux I__9312 (
            .O(N__49258),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18352 ));
    InMux I__9311 (
            .O(N__49255),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787 ));
    CascadeMux I__9310 (
            .O(N__49252),
            .I(N__49249));
    InMux I__9309 (
            .O(N__49249),
            .I(N__49246));
    LocalMux I__9308 (
            .O(N__49246),
            .I(N__49243));
    Span4Mux_v I__9307 (
            .O(N__49243),
            .I(N__49240));
    Odrv4 I__9306 (
            .O(N__49240),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO ));
    InMux I__9305 (
            .O(N__49237),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747 ));
    CascadeMux I__9304 (
            .O(N__49234),
            .I(N__49231));
    InMux I__9303 (
            .O(N__49231),
            .I(N__49228));
    LocalMux I__9302 (
            .O(N__49228),
            .I(N__49225));
    Odrv12 I__9301 (
            .O(N__49225),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO ));
    InMux I__9300 (
            .O(N__49222),
            .I(N__49219));
    LocalMux I__9299 (
            .O(N__49219),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n90 ));
    InMux I__9298 (
            .O(N__49216),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18339 ));
    CascadeMux I__9297 (
            .O(N__49213),
            .I(N__49210));
    InMux I__9296 (
            .O(N__49210),
            .I(N__49207));
    LocalMux I__9295 (
            .O(N__49207),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n139 ));
    InMux I__9294 (
            .O(N__49204),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18340 ));
    InMux I__9293 (
            .O(N__49201),
            .I(N__49198));
    LocalMux I__9292 (
            .O(N__49198),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n188 ));
    InMux I__9291 (
            .O(N__49195),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18341 ));
    InMux I__9290 (
            .O(N__49192),
            .I(N__49189));
    LocalMux I__9289 (
            .O(N__49189),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n237 ));
    InMux I__9288 (
            .O(N__49186),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18342 ));
    InMux I__9287 (
            .O(N__49183),
            .I(N__49180));
    LocalMux I__9286 (
            .O(N__49180),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n286 ));
    InMux I__9285 (
            .O(N__49177),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18343 ));
    InMux I__9284 (
            .O(N__49174),
            .I(N__49171));
    LocalMux I__9283 (
            .O(N__49171),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n335 ));
    InMux I__9282 (
            .O(N__49168),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18344 ));
    InMux I__9281 (
            .O(N__49165),
            .I(N__49162));
    LocalMux I__9280 (
            .O(N__49162),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n384 ));
    InMux I__9279 (
            .O(N__49159),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18345 ));
    InMux I__9278 (
            .O(N__49156),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18194 ));
    InMux I__9277 (
            .O(N__49153),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18195 ));
    InMux I__9276 (
            .O(N__49150),
            .I(bfn_19_25_0_));
    InMux I__9275 (
            .O(N__49147),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18197 ));
    InMux I__9274 (
            .O(N__49144),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18198 ));
    InMux I__9273 (
            .O(N__49141),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18199 ));
    InMux I__9272 (
            .O(N__49138),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18200 ));
    InMux I__9271 (
            .O(N__49135),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18201 ));
    InMux I__9270 (
            .O(N__49132),
            .I(N__49129));
    LocalMux I__9269 (
            .O(N__49129),
            .I(N__49126));
    Odrv12 I__9268 (
            .O(N__49126),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n746 ));
    InMux I__9267 (
            .O(N__49123),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18202 ));
    InMux I__9266 (
            .O(N__49120),
            .I(N__49117));
    LocalMux I__9265 (
            .O(N__49117),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n60 ));
    InMux I__9264 (
            .O(N__49114),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18189 ));
    InMux I__9263 (
            .O(N__49111),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18190 ));
    InMux I__9262 (
            .O(N__49108),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18191 ));
    InMux I__9261 (
            .O(N__49105),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18192 ));
    InMux I__9260 (
            .O(N__49102),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18193 ));
    InMux I__9259 (
            .O(N__49099),
            .I(bfn_19_22_0_));
    InMux I__9258 (
            .O(N__49096),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18152 ));
    InMux I__9257 (
            .O(N__49093),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18153 ));
    InMux I__9256 (
            .O(N__49090),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18154 ));
    InMux I__9255 (
            .O(N__49087),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18155 ));
    InMux I__9254 (
            .O(N__49084),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18156 ));
    InMux I__9253 (
            .O(N__49081),
            .I(N__49078));
    LocalMux I__9252 (
            .O(N__49078),
            .I(N__49075));
    Span4Mux_v I__9251 (
            .O(N__49075),
            .I(N__49072));
    Odrv4 I__9250 (
            .O(N__49072),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n790 ));
    InMux I__9249 (
            .O(N__49069),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18157 ));
    InMux I__9248 (
            .O(N__49066),
            .I(N__49063));
    LocalMux I__9247 (
            .O(N__49063),
            .I(N__49060));
    Span4Mux_h I__9246 (
            .O(N__49060),
            .I(N__49057));
    Span4Mux_v I__9245 (
            .O(N__49057),
            .I(N__49054));
    Odrv4 I__9244 (
            .O(N__49054),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n794 ));
    CascadeMux I__9243 (
            .O(N__49051),
            .I(N__49048));
    InMux I__9242 (
            .O(N__49048),
            .I(N__49045));
    LocalMux I__9241 (
            .O(N__49045),
            .I(N__49042));
    Span12Mux_h I__9240 (
            .O(N__49042),
            .I(N__49039));
    Odrv12 I__9239 (
            .O(N__49039),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO ));
    InMux I__9238 (
            .O(N__49036),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18158 ));
    InMux I__9237 (
            .O(N__49033),
            .I(N__49030));
    LocalMux I__9236 (
            .O(N__49030),
            .I(N__49027));
    Span4Mux_h I__9235 (
            .O(N__49027),
            .I(N__49024));
    Odrv4 I__9234 (
            .O(N__49024),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO ));
    CascadeMux I__9233 (
            .O(N__49021),
            .I(N__49018));
    InMux I__9232 (
            .O(N__49018),
            .I(N__49015));
    LocalMux I__9231 (
            .O(N__49015),
            .I(N__49012));
    Span4Mux_v I__9230 (
            .O(N__49012),
            .I(N__49008));
    InMux I__9229 (
            .O(N__49011),
            .I(N__49005));
    Span4Mux_h I__9228 (
            .O(N__49008),
            .I(N__49002));
    LocalMux I__9227 (
            .O(N__49005),
            .I(N__48999));
    Odrv4 I__9226 (
            .O(N__49002),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n796 ));
    Odrv4 I__9225 (
            .O(N__48999),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n796 ));
    InMux I__9224 (
            .O(N__48994),
            .I(bfn_19_23_0_));
    CascadeMux I__9223 (
            .O(N__48991),
            .I(N__48988));
    InMux I__9222 (
            .O(N__48988),
            .I(N__48984));
    InMux I__9221 (
            .O(N__48987),
            .I(N__48981));
    LocalMux I__9220 (
            .O(N__48984),
            .I(N__48976));
    LocalMux I__9219 (
            .O(N__48981),
            .I(N__48976));
    Odrv4 I__9218 (
            .O(N__48976),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n738 ));
    CascadeMux I__9217 (
            .O(N__48973),
            .I(N__48970));
    InMux I__9216 (
            .O(N__48970),
            .I(N__48962));
    InMux I__9215 (
            .O(N__48969),
            .I(N__48962));
    InMux I__9214 (
            .O(N__48968),
            .I(N__48959));
    InMux I__9213 (
            .O(N__48967),
            .I(N__48956));
    LocalMux I__9212 (
            .O(N__48962),
            .I(N__48953));
    LocalMux I__9211 (
            .O(N__48959),
            .I(N__48947));
    LocalMux I__9210 (
            .O(N__48956),
            .I(N__48947));
    Sp12to4 I__9209 (
            .O(N__48953),
            .I(N__48944));
    InMux I__9208 (
            .O(N__48952),
            .I(N__48941));
    Span4Mux_v I__9207 (
            .O(N__48947),
            .I(N__48936));
    Span12Mux_v I__9206 (
            .O(N__48944),
            .I(N__48931));
    LocalMux I__9205 (
            .O(N__48941),
            .I(N__48931));
    InMux I__9204 (
            .O(N__48940),
            .I(N__48926));
    InMux I__9203 (
            .O(N__48939),
            .I(N__48926));
    Odrv4 I__9202 (
            .O(N__48936),
            .I(Error_sub_temp_31_adj_2384));
    Odrv12 I__9201 (
            .O(N__48931),
            .I(Error_sub_temp_31_adj_2384));
    LocalMux I__9200 (
            .O(N__48926),
            .I(Error_sub_temp_31_adj_2384));
    InMux I__9199 (
            .O(N__48919),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18144 ));
    InMux I__9198 (
            .O(N__48916),
            .I(N__48913));
    LocalMux I__9197 (
            .O(N__48913),
            .I(N__48910));
    Odrv4 I__9196 (
            .O(N__48910),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n8356 ));
    InMux I__9195 (
            .O(N__48907),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18145 ));
    InMux I__9194 (
            .O(N__48904),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18146 ));
    InMux I__9193 (
            .O(N__48901),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18147 ));
    InMux I__9192 (
            .O(N__48898),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18148 ));
    InMux I__9191 (
            .O(N__48895),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18149 ));
    InMux I__9190 (
            .O(N__48892),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18150 ));
    InMux I__9189 (
            .O(N__48889),
            .I(N__48886));
    LocalMux I__9188 (
            .O(N__48886),
            .I(N__48883));
    Span4Mux_v I__9187 (
            .O(N__48883),
            .I(N__48880));
    Span4Mux_v I__9186 (
            .O(N__48880),
            .I(N__48877));
    Odrv4 I__9185 (
            .O(N__48877),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO ));
    InMux I__9184 (
            .O(N__48874),
            .I(bfn_19_19_0_));
    InMux I__9183 (
            .O(N__48871),
            .I(N__48868));
    LocalMux I__9182 (
            .O(N__48868),
            .I(N__48864));
    InMux I__9181 (
            .O(N__48867),
            .I(N__48861));
    Odrv4 I__9180 (
            .O(N__48864),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8 ));
    LocalMux I__9179 (
            .O(N__48861),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8 ));
    InMux I__9178 (
            .O(N__48856),
            .I(N__48853));
    LocalMux I__9177 (
            .O(N__48853),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20870 ));
    CascadeMux I__9176 (
            .O(N__48850),
            .I(N__48847));
    InMux I__9175 (
            .O(N__48847),
            .I(N__48844));
    LocalMux I__9174 (
            .O(N__48844),
            .I(N__48841));
    Span12Mux_h I__9173 (
            .O(N__48841),
            .I(N__48836));
    InMux I__9172 (
            .O(N__48840),
            .I(N__48833));
    InMux I__9171 (
            .O(N__48839),
            .I(N__48830));
    Odrv12 I__9170 (
            .O(N__48836),
            .I(\foc.preSatVoltage_10 ));
    LocalMux I__9169 (
            .O(N__48833),
            .I(\foc.preSatVoltage_10 ));
    LocalMux I__9168 (
            .O(N__48830),
            .I(\foc.preSatVoltage_10 ));
    InMux I__9167 (
            .O(N__48823),
            .I(N__48820));
    LocalMux I__9166 (
            .O(N__48820),
            .I(N__48816));
    InMux I__9165 (
            .O(N__48819),
            .I(N__48813));
    Odrv4 I__9164 (
            .O(N__48816),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9 ));
    LocalMux I__9163 (
            .O(N__48813),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9 ));
    InMux I__9162 (
            .O(N__48808),
            .I(N__48805));
    LocalMux I__9161 (
            .O(N__48805),
            .I(N__48802));
    Odrv12 I__9160 (
            .O(N__48802),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO ));
    CascadeMux I__9159 (
            .O(N__48799),
            .I(N__48796));
    InMux I__9158 (
            .O(N__48796),
            .I(N__48793));
    LocalMux I__9157 (
            .O(N__48793),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n766 ));
    InMux I__9156 (
            .O(N__48790),
            .I(bfn_19_18_0_));
    InMux I__9155 (
            .O(N__48787),
            .I(N__48784));
    LocalMux I__9154 (
            .O(N__48784),
            .I(N__48781));
    Odrv4 I__9153 (
            .O(N__48781),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n770 ));
    CascadeMux I__9152 (
            .O(N__48778),
            .I(N__48775));
    InMux I__9151 (
            .O(N__48775),
            .I(N__48772));
    LocalMux I__9150 (
            .O(N__48772),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO ));
    InMux I__9149 (
            .O(N__48769),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17719 ));
    InMux I__9148 (
            .O(N__48766),
            .I(N__48763));
    LocalMux I__9147 (
            .O(N__48763),
            .I(N__48760));
    Span4Mux_v I__9146 (
            .O(N__48760),
            .I(N__48757));
    Odrv4 I__9145 (
            .O(N__48757),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n774 ));
    CascadeMux I__9144 (
            .O(N__48754),
            .I(N__48751));
    InMux I__9143 (
            .O(N__48751),
            .I(N__48748));
    LocalMux I__9142 (
            .O(N__48748),
            .I(N__48745));
    Span4Mux_v I__9141 (
            .O(N__48745),
            .I(N__48742));
    Odrv4 I__9140 (
            .O(N__48742),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO ));
    InMux I__9139 (
            .O(N__48739),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17720 ));
    InMux I__9138 (
            .O(N__48736),
            .I(N__48733));
    LocalMux I__9137 (
            .O(N__48733),
            .I(N__48730));
    Sp12to4 I__9136 (
            .O(N__48730),
            .I(N__48727));
    Span12Mux_v I__9135 (
            .O(N__48727),
            .I(N__48724));
    Odrv12 I__9134 (
            .O(N__48724),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n778 ));
    CascadeMux I__9133 (
            .O(N__48721),
            .I(N__48718));
    InMux I__9132 (
            .O(N__48718),
            .I(N__48715));
    LocalMux I__9131 (
            .O(N__48715),
            .I(N__48712));
    Span4Mux_v I__9130 (
            .O(N__48712),
            .I(N__48709));
    Odrv4 I__9129 (
            .O(N__48709),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO ));
    InMux I__9128 (
            .O(N__48706),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17721 ));
    CascadeMux I__9127 (
            .O(N__48703),
            .I(N__48700));
    InMux I__9126 (
            .O(N__48700),
            .I(N__48697));
    LocalMux I__9125 (
            .O(N__48697),
            .I(N__48694));
    Span12Mux_v I__9124 (
            .O(N__48694),
            .I(N__48691));
    Odrv12 I__9123 (
            .O(N__48691),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO ));
    InMux I__9122 (
            .O(N__48688),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17722 ));
    InMux I__9121 (
            .O(N__48685),
            .I(N__48682));
    LocalMux I__9120 (
            .O(N__48682),
            .I(N__48679));
    Odrv12 I__9119 (
            .O(N__48679),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n786 ));
    InMux I__9118 (
            .O(N__48676),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17723 ));
    InMux I__9117 (
            .O(N__48673),
            .I(N__48670));
    LocalMux I__9116 (
            .O(N__48670),
            .I(N__48667));
    Span12Mux_v I__9115 (
            .O(N__48667),
            .I(N__48664));
    Odrv12 I__9114 (
            .O(N__48664),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415 ));
    CascadeMux I__9113 (
            .O(N__48661),
            .I(N__48658));
    InMux I__9112 (
            .O(N__48658),
            .I(N__48655));
    LocalMux I__9111 (
            .O(N__48655),
            .I(N__48652));
    Span4Mux_v I__9110 (
            .O(N__48652),
            .I(N__48649));
    Odrv4 I__9109 (
            .O(N__48649),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO ));
    InMux I__9108 (
            .O(N__48646),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17724 ));
    InMux I__9107 (
            .O(N__48643),
            .I(N__48640));
    LocalMux I__9106 (
            .O(N__48640),
            .I(N__48637));
    Span4Mux_v I__9105 (
            .O(N__48637),
            .I(N__48634));
    Span4Mux_v I__9104 (
            .O(N__48634),
            .I(N__48631));
    Odrv4 I__9103 (
            .O(N__48631),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413 ));
    CascadeMux I__9102 (
            .O(N__48628),
            .I(N__48625));
    InMux I__9101 (
            .O(N__48625),
            .I(N__48622));
    LocalMux I__9100 (
            .O(N__48622),
            .I(N__48619));
    Sp12to4 I__9099 (
            .O(N__48619),
            .I(N__48616));
    Odrv12 I__9098 (
            .O(N__48616),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO ));
    InMux I__9097 (
            .O(N__48613),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17725 ));
    InMux I__9096 (
            .O(N__48610),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17711 ));
    InMux I__9095 (
            .O(N__48607),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17712 ));
    InMux I__9094 (
            .O(N__48604),
            .I(N__48601));
    LocalMux I__9093 (
            .O(N__48601),
            .I(N__48598));
    Odrv4 I__9092 (
            .O(N__48598),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n746 ));
    InMux I__9091 (
            .O(N__48595),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17713 ));
    InMux I__9090 (
            .O(N__48592),
            .I(N__48589));
    LocalMux I__9089 (
            .O(N__48589),
            .I(N__48586));
    Span4Mux_v I__9088 (
            .O(N__48586),
            .I(N__48583));
    Odrv4 I__9087 (
            .O(N__48583),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n750 ));
    CascadeMux I__9086 (
            .O(N__48580),
            .I(N__48577));
    InMux I__9085 (
            .O(N__48577),
            .I(N__48574));
    LocalMux I__9084 (
            .O(N__48574),
            .I(N__48571));
    Span4Mux_v I__9083 (
            .O(N__48571),
            .I(N__48568));
    Odrv4 I__9082 (
            .O(N__48568),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO ));
    InMux I__9081 (
            .O(N__48565),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17714 ));
    InMux I__9080 (
            .O(N__48562),
            .I(N__48559));
    LocalMux I__9079 (
            .O(N__48559),
            .I(N__48556));
    Span4Mux_v I__9078 (
            .O(N__48556),
            .I(N__48553));
    Span4Mux_h I__9077 (
            .O(N__48553),
            .I(N__48550));
    Odrv4 I__9076 (
            .O(N__48550),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n754 ));
    CascadeMux I__9075 (
            .O(N__48547),
            .I(N__48544));
    InMux I__9074 (
            .O(N__48544),
            .I(N__48541));
    LocalMux I__9073 (
            .O(N__48541),
            .I(N__48538));
    Span4Mux_v I__9072 (
            .O(N__48538),
            .I(N__48535));
    Odrv4 I__9071 (
            .O(N__48535),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO ));
    InMux I__9070 (
            .O(N__48532),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17715 ));
    InMux I__9069 (
            .O(N__48529),
            .I(N__48526));
    LocalMux I__9068 (
            .O(N__48526),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n758 ));
    CascadeMux I__9067 (
            .O(N__48523),
            .I(N__48520));
    InMux I__9066 (
            .O(N__48520),
            .I(N__48517));
    LocalMux I__9065 (
            .O(N__48517),
            .I(N__48514));
    Span4Mux_h I__9064 (
            .O(N__48514),
            .I(N__48511));
    Odrv4 I__9063 (
            .O(N__48511),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO ));
    InMux I__9062 (
            .O(N__48508),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17716 ));
    InMux I__9061 (
            .O(N__48505),
            .I(N__48502));
    LocalMux I__9060 (
            .O(N__48502),
            .I(N__48499));
    Odrv4 I__9059 (
            .O(N__48499),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n762 ));
    CascadeMux I__9058 (
            .O(N__48496),
            .I(N__48493));
    InMux I__9057 (
            .O(N__48493),
            .I(N__48490));
    LocalMux I__9056 (
            .O(N__48490),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO ));
    InMux I__9055 (
            .O(N__48487),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17717 ));
    CascadeMux I__9054 (
            .O(N__48484),
            .I(N__48481));
    InMux I__9053 (
            .O(N__48481),
            .I(N__48478));
    LocalMux I__9052 (
            .O(N__48478),
            .I(N__48475));
    Odrv4 I__9051 (
            .O(N__48475),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n412 ));
    InMux I__9050 (
            .O(N__48472),
            .I(N__48469));
    LocalMux I__9049 (
            .O(N__48469),
            .I(N__48466));
    Odrv4 I__9048 (
            .O(N__48466),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n458 ));
    InMux I__9047 (
            .O(N__48463),
            .I(bfn_19_16_0_));
    InMux I__9046 (
            .O(N__48460),
            .I(N__48457));
    LocalMux I__9045 (
            .O(N__48457),
            .I(N__48454));
    Odrv12 I__9044 (
            .O(N__48454),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n461 ));
    InMux I__9043 (
            .O(N__48451),
            .I(N__48448));
    LocalMux I__9042 (
            .O(N__48448),
            .I(N__48445));
    Odrv12 I__9041 (
            .O(N__48445),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n507 ));
    InMux I__9040 (
            .O(N__48442),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17804 ));
    InMux I__9039 (
            .O(N__48439),
            .I(N__48436));
    LocalMux I__9038 (
            .O(N__48436),
            .I(N__48433));
    Odrv4 I__9037 (
            .O(N__48433),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n510 ));
    InMux I__9036 (
            .O(N__48430),
            .I(N__48427));
    LocalMux I__9035 (
            .O(N__48427),
            .I(N__48424));
    Odrv4 I__9034 (
            .O(N__48424),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370 ));
    InMux I__9033 (
            .O(N__48421),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17805 ));
    InMux I__9032 (
            .O(N__48418),
            .I(N__48415));
    LocalMux I__9031 (
            .O(N__48415),
            .I(N__48412));
    Odrv12 I__9030 (
            .O(N__48412),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358 ));
    InMux I__9029 (
            .O(N__48409),
            .I(N__48406));
    LocalMux I__9028 (
            .O(N__48406),
            .I(N__48403));
    Odrv12 I__9027 (
            .O(N__48403),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462 ));
    InMux I__9026 (
            .O(N__48400),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17806 ));
    InMux I__9025 (
            .O(N__48397),
            .I(N__48394));
    LocalMux I__9024 (
            .O(N__48394),
            .I(N__48391));
    Odrv4 I__9023 (
            .O(N__48391),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377 ));
    CascadeMux I__9022 (
            .O(N__48388),
            .I(N__48385));
    InMux I__9021 (
            .O(N__48385),
            .I(N__48382));
    LocalMux I__9020 (
            .O(N__48382),
            .I(N__48379));
    Odrv4 I__9019 (
            .O(N__48379),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456 ));
    InMux I__9018 (
            .O(N__48376),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17807 ));
    CascadeMux I__9017 (
            .O(N__48373),
            .I(N__48370));
    InMux I__9016 (
            .O(N__48370),
            .I(N__48367));
    LocalMux I__9015 (
            .O(N__48367),
            .I(N__48364));
    Odrv4 I__9014 (
            .O(N__48364),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360 ));
    CascadeMux I__9013 (
            .O(N__48361),
            .I(N__48358));
    InMux I__9012 (
            .O(N__48358),
            .I(N__48355));
    LocalMux I__9011 (
            .O(N__48355),
            .I(N__48352));
    Odrv12 I__9010 (
            .O(N__48352),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359 ));
    InMux I__9009 (
            .O(N__48349),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17808 ));
    CascadeMux I__9008 (
            .O(N__48346),
            .I(N__48343));
    InMux I__9007 (
            .O(N__48343),
            .I(N__48340));
    LocalMux I__9006 (
            .O(N__48340),
            .I(N__48337));
    Odrv12 I__9005 (
            .O(N__48337),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371 ));
    InMux I__9004 (
            .O(N__48334),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17809 ));
    InMux I__9003 (
            .O(N__48331),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354 ));
    InMux I__9002 (
            .O(N__48328),
            .I(N__48325));
    LocalMux I__9001 (
            .O(N__48325),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n69 ));
    InMux I__9000 (
            .O(N__48322),
            .I(N__48319));
    LocalMux I__8999 (
            .O(N__48319),
            .I(N__48316));
    Odrv12 I__8998 (
            .O(N__48316),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n115 ));
    InMux I__8997 (
            .O(N__48313),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17796 ));
    InMux I__8996 (
            .O(N__48310),
            .I(N__48307));
    LocalMux I__8995 (
            .O(N__48307),
            .I(N__48304));
    Odrv4 I__8994 (
            .O(N__48304),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n118 ));
    InMux I__8993 (
            .O(N__48301),
            .I(N__48298));
    LocalMux I__8992 (
            .O(N__48298),
            .I(N__48295));
    Odrv4 I__8991 (
            .O(N__48295),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n164 ));
    InMux I__8990 (
            .O(N__48292),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17797 ));
    CascadeMux I__8989 (
            .O(N__48289),
            .I(N__48286));
    InMux I__8988 (
            .O(N__48286),
            .I(N__48283));
    LocalMux I__8987 (
            .O(N__48283),
            .I(N__48280));
    Odrv4 I__8986 (
            .O(N__48280),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n167 ));
    InMux I__8985 (
            .O(N__48277),
            .I(N__48274));
    LocalMux I__8984 (
            .O(N__48274),
            .I(N__48271));
    Odrv12 I__8983 (
            .O(N__48271),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n213 ));
    InMux I__8982 (
            .O(N__48268),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17798 ));
    InMux I__8981 (
            .O(N__48265),
            .I(N__48262));
    LocalMux I__8980 (
            .O(N__48262),
            .I(N__48259));
    Odrv4 I__8979 (
            .O(N__48259),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n216 ));
    InMux I__8978 (
            .O(N__48256),
            .I(N__48253));
    LocalMux I__8977 (
            .O(N__48253),
            .I(N__48250));
    Odrv4 I__8976 (
            .O(N__48250),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425 ));
    InMux I__8975 (
            .O(N__48247),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17799 ));
    InMux I__8974 (
            .O(N__48244),
            .I(N__48241));
    LocalMux I__8973 (
            .O(N__48241),
            .I(N__48238));
    Odrv4 I__8972 (
            .O(N__48238),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n265 ));
    CascadeMux I__8971 (
            .O(N__48235),
            .I(N__48232));
    InMux I__8970 (
            .O(N__48232),
            .I(N__48229));
    LocalMux I__8969 (
            .O(N__48229),
            .I(N__48226));
    Odrv4 I__8968 (
            .O(N__48226),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422 ));
    InMux I__8967 (
            .O(N__48223),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17800 ));
    InMux I__8966 (
            .O(N__48220),
            .I(N__48217));
    LocalMux I__8965 (
            .O(N__48217),
            .I(N__48214));
    Odrv12 I__8964 (
            .O(N__48214),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401 ));
    CascadeMux I__8963 (
            .O(N__48211),
            .I(N__48208));
    InMux I__8962 (
            .O(N__48208),
            .I(N__48205));
    LocalMux I__8961 (
            .O(N__48205),
            .I(N__48202));
    Odrv12 I__8960 (
            .O(N__48202),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n360 ));
    InMux I__8959 (
            .O(N__48199),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17801 ));
    InMux I__8958 (
            .O(N__48196),
            .I(N__48193));
    LocalMux I__8957 (
            .O(N__48193),
            .I(N__48190));
    Odrv4 I__8956 (
            .O(N__48190),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380 ));
    InMux I__8955 (
            .O(N__48187),
            .I(N__48184));
    LocalMux I__8954 (
            .O(N__48184),
            .I(N__48181));
    Span4Mux_v I__8953 (
            .O(N__48181),
            .I(N__48178));
    Odrv4 I__8952 (
            .O(N__48178),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n409 ));
    InMux I__8951 (
            .O(N__48175),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17802 ));
    InMux I__8950 (
            .O(N__48172),
            .I(N__48169));
    LocalMux I__8949 (
            .O(N__48169),
            .I(N__48166));
    Span4Mux_h I__8948 (
            .O(N__48166),
            .I(N__48163));
    Odrv4 I__8947 (
            .O(N__48163),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426 ));
    InMux I__8946 (
            .O(N__48160),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17817 ));
    CascadeMux I__8945 (
            .O(N__48157),
            .I(N__48154));
    InMux I__8944 (
            .O(N__48154),
            .I(N__48151));
    LocalMux I__8943 (
            .O(N__48151),
            .I(N__48148));
    Odrv4 I__8942 (
            .O(N__48148),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n415 ));
    InMux I__8941 (
            .O(N__48145),
            .I(bfn_19_14_0_));
    InMux I__8940 (
            .O(N__48142),
            .I(N__48139));
    LocalMux I__8939 (
            .O(N__48139),
            .I(N__48136));
    Span4Mux_v I__8938 (
            .O(N__48136),
            .I(N__48133));
    Odrv4 I__8937 (
            .O(N__48133),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423 ));
    InMux I__8936 (
            .O(N__48130),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17819 ));
    InMux I__8935 (
            .O(N__48127),
            .I(N__48124));
    LocalMux I__8934 (
            .O(N__48124),
            .I(N__48121));
    Odrv4 I__8933 (
            .O(N__48121),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412 ));
    InMux I__8932 (
            .O(N__48118),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17820 ));
    InMux I__8931 (
            .O(N__48115),
            .I(N__48112));
    LocalMux I__8930 (
            .O(N__48112),
            .I(N__48109));
    Odrv4 I__8929 (
            .O(N__48109),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378 ));
    InMux I__8928 (
            .O(N__48106),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17821 ));
    CascadeMux I__8927 (
            .O(N__48103),
            .I(N__48100));
    InMux I__8926 (
            .O(N__48100),
            .I(N__48097));
    LocalMux I__8925 (
            .O(N__48097),
            .I(N__48094));
    Odrv4 I__8924 (
            .O(N__48094),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373 ));
    InMux I__8923 (
            .O(N__48091),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17822 ));
    InMux I__8922 (
            .O(N__48088),
            .I(N__48085));
    LocalMux I__8921 (
            .O(N__48085),
            .I(N__48082));
    Span4Mux_v I__8920 (
            .O(N__48082),
            .I(N__48079));
    Odrv4 I__8919 (
            .O(N__48079),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372 ));
    InMux I__8918 (
            .O(N__48076),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17823 ));
    CascadeMux I__8917 (
            .O(N__48073),
            .I(N__48070));
    InMux I__8916 (
            .O(N__48070),
            .I(N__48067));
    LocalMux I__8915 (
            .O(N__48067),
            .I(N__48064));
    Odrv4 I__8914 (
            .O(N__48064),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n709 ));
    InMux I__8913 (
            .O(N__48061),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17824 ));
    InMux I__8912 (
            .O(N__48058),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n763 ));
    InMux I__8911 (
            .O(N__48055),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421 ));
    CascadeMux I__8910 (
            .O(N__48052),
            .I(N__48049));
    InMux I__8909 (
            .O(N__48049),
            .I(N__48046));
    LocalMux I__8908 (
            .O(N__48046),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n72 ));
    InMux I__8907 (
            .O(N__48043),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17811 ));
    InMux I__8906 (
            .O(N__48040),
            .I(N__48037));
    LocalMux I__8905 (
            .O(N__48037),
            .I(N__48034));
    Odrv4 I__8904 (
            .O(N__48034),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n121 ));
    InMux I__8903 (
            .O(N__48031),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17812 ));
    InMux I__8902 (
            .O(N__48028),
            .I(N__48025));
    LocalMux I__8901 (
            .O(N__48025),
            .I(N__48022));
    Odrv4 I__8900 (
            .O(N__48022),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n170 ));
    InMux I__8899 (
            .O(N__48019),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17813 ));
    InMux I__8898 (
            .O(N__48016),
            .I(N__48013));
    LocalMux I__8897 (
            .O(N__48013),
            .I(N__48010));
    Odrv4 I__8896 (
            .O(N__48010),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n219 ));
    InMux I__8895 (
            .O(N__48007),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17814 ));
    InMux I__8894 (
            .O(N__48004),
            .I(N__48001));
    LocalMux I__8893 (
            .O(N__48001),
            .I(N__47998));
    Odrv4 I__8892 (
            .O(N__47998),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437 ));
    InMux I__8891 (
            .O(N__47995),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17815 ));
    CascadeMux I__8890 (
            .O(N__47992),
            .I(N__47989));
    InMux I__8889 (
            .O(N__47989),
            .I(N__47986));
    LocalMux I__8888 (
            .O(N__47986),
            .I(N__47983));
    Odrv4 I__8887 (
            .O(N__47983),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428 ));
    InMux I__8886 (
            .O(N__47980),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17816 ));
    InMux I__8885 (
            .O(N__47977),
            .I(N__47974));
    LocalMux I__8884 (
            .O(N__47974),
            .I(N__47971));
    Odrv12 I__8883 (
            .O(N__47971),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n335 ));
    InMux I__8882 (
            .O(N__47968),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17917 ));
    InMux I__8881 (
            .O(N__47965),
            .I(N__47962));
    LocalMux I__8880 (
            .O(N__47962),
            .I(N__47959));
    Odrv4 I__8879 (
            .O(N__47959),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n384 ));
    InMux I__8878 (
            .O(N__47956),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17918 ));
    InMux I__8877 (
            .O(N__47953),
            .I(N__47950));
    LocalMux I__8876 (
            .O(N__47950),
            .I(N__47947));
    Odrv12 I__8875 (
            .O(N__47947),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n433 ));
    InMux I__8874 (
            .O(N__47944),
            .I(bfn_19_12_0_));
    InMux I__8873 (
            .O(N__47941),
            .I(N__47938));
    LocalMux I__8872 (
            .O(N__47938),
            .I(N__47935));
    Odrv4 I__8871 (
            .O(N__47935),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n482 ));
    InMux I__8870 (
            .O(N__47932),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17920 ));
    InMux I__8869 (
            .O(N__47929),
            .I(N__47926));
    LocalMux I__8868 (
            .O(N__47926),
            .I(N__47923));
    Odrv4 I__8867 (
            .O(N__47923),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n531 ));
    InMux I__8866 (
            .O(N__47920),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17921 ));
    InMux I__8865 (
            .O(N__47917),
            .I(N__47914));
    LocalMux I__8864 (
            .O(N__47914),
            .I(N__47911));
    Odrv12 I__8863 (
            .O(N__47911),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n580 ));
    InMux I__8862 (
            .O(N__47908),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17922 ));
    InMux I__8861 (
            .O(N__47905),
            .I(N__47902));
    LocalMux I__8860 (
            .O(N__47902),
            .I(N__47899));
    Odrv4 I__8859 (
            .O(N__47899),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n629 ));
    InMux I__8858 (
            .O(N__47896),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17923 ));
    CascadeMux I__8857 (
            .O(N__47893),
            .I(N__47890));
    InMux I__8856 (
            .O(N__47890),
            .I(N__47887));
    LocalMux I__8855 (
            .O(N__47887),
            .I(N__47884));
    Span4Mux_v I__8854 (
            .O(N__47884),
            .I(N__47881));
    Odrv4 I__8853 (
            .O(N__47881),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n678 ));
    InMux I__8852 (
            .O(N__47878),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17924 ));
    CascadeMux I__8851 (
            .O(N__47875),
            .I(N__47872));
    InMux I__8850 (
            .O(N__47872),
            .I(N__47869));
    LocalMux I__8849 (
            .O(N__47869),
            .I(N__47866));
    Odrv4 I__8848 (
            .O(N__47866),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n727 ));
    InMux I__8847 (
            .O(N__47863),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17925 ));
    CascadeMux I__8846 (
            .O(N__47860),
            .I(N__47857));
    InMux I__8845 (
            .O(N__47857),
            .I(N__47854));
    LocalMux I__8844 (
            .O(N__47854),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n730 ));
    InMux I__8843 (
            .O(N__47851),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17940 ));
    InMux I__8842 (
            .O(N__47848),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416 ));
    CascadeMux I__8841 (
            .O(N__47845),
            .I(N__47842));
    InMux I__8840 (
            .O(N__47842),
            .I(N__47839));
    LocalMux I__8839 (
            .O(N__47839),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420 ));
    InMux I__8838 (
            .O(N__47836),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17912 ));
    InMux I__8837 (
            .O(N__47833),
            .I(N__47830));
    LocalMux I__8836 (
            .O(N__47830),
            .I(N__47827));
    Odrv4 I__8835 (
            .O(N__47827),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419 ));
    InMux I__8834 (
            .O(N__47824),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17913 ));
    InMux I__8833 (
            .O(N__47821),
            .I(N__47818));
    LocalMux I__8832 (
            .O(N__47818),
            .I(N__47815));
    Odrv12 I__8831 (
            .O(N__47815),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418 ));
    InMux I__8830 (
            .O(N__47812),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17914 ));
    InMux I__8829 (
            .O(N__47809),
            .I(N__47806));
    LocalMux I__8828 (
            .O(N__47806),
            .I(N__47803));
    Odrv4 I__8827 (
            .O(N__47803),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417 ));
    InMux I__8826 (
            .O(N__47800),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17915 ));
    InMux I__8825 (
            .O(N__47797),
            .I(N__47794));
    LocalMux I__8824 (
            .O(N__47794),
            .I(N__47791));
    Odrv4 I__8823 (
            .O(N__47791),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n286 ));
    InMux I__8822 (
            .O(N__47788),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17916 ));
    InMux I__8821 (
            .O(N__47785),
            .I(N__47782));
    LocalMux I__8820 (
            .O(N__47782),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n289 ));
    InMux I__8819 (
            .O(N__47779),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17931 ));
    InMux I__8818 (
            .O(N__47776),
            .I(N__47773));
    LocalMux I__8817 (
            .O(N__47773),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n338 ));
    InMux I__8816 (
            .O(N__47770),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17932 ));
    InMux I__8815 (
            .O(N__47767),
            .I(N__47764));
    LocalMux I__8814 (
            .O(N__47764),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n387 ));
    InMux I__8813 (
            .O(N__47761),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17933 ));
    CascadeMux I__8812 (
            .O(N__47758),
            .I(N__47755));
    InMux I__8811 (
            .O(N__47755),
            .I(N__47752));
    LocalMux I__8810 (
            .O(N__47752),
            .I(N__47749));
    Odrv4 I__8809 (
            .O(N__47749),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n436 ));
    InMux I__8808 (
            .O(N__47746),
            .I(bfn_19_10_0_));
    InMux I__8807 (
            .O(N__47743),
            .I(N__47740));
    LocalMux I__8806 (
            .O(N__47740),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n485 ));
    InMux I__8805 (
            .O(N__47737),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17935 ));
    InMux I__8804 (
            .O(N__47734),
            .I(N__47731));
    LocalMux I__8803 (
            .O(N__47731),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n534 ));
    InMux I__8802 (
            .O(N__47728),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17936 ));
    InMux I__8801 (
            .O(N__47725),
            .I(N__47722));
    LocalMux I__8800 (
            .O(N__47722),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n583 ));
    InMux I__8799 (
            .O(N__47719),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17937 ));
    InMux I__8798 (
            .O(N__47716),
            .I(N__47713));
    LocalMux I__8797 (
            .O(N__47713),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n632 ));
    InMux I__8796 (
            .O(N__47710),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17938 ));
    CascadeMux I__8795 (
            .O(N__47707),
            .I(N__47704));
    InMux I__8794 (
            .O(N__47704),
            .I(N__47701));
    LocalMux I__8793 (
            .O(N__47701),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n681 ));
    InMux I__8792 (
            .O(N__47698),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17939 ));
    CascadeMux I__8791 (
            .O(N__47695),
            .I(N__47692));
    InMux I__8790 (
            .O(N__47692),
            .I(N__47689));
    LocalMux I__8789 (
            .O(N__47689),
            .I(N__47686));
    Odrv4 I__8788 (
            .O(N__47686),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n663 ));
    InMux I__8787 (
            .O(N__47683),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17638 ));
    InMux I__8786 (
            .O(N__47680),
            .I(N__47676));
    InMux I__8785 (
            .O(N__47679),
            .I(N__47673));
    LocalMux I__8784 (
            .O(N__47676),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n765 ));
    LocalMux I__8783 (
            .O(N__47673),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n765 ));
    CascadeMux I__8782 (
            .O(N__47668),
            .I(N__47665));
    InMux I__8781 (
            .O(N__47665),
            .I(N__47662));
    LocalMux I__8780 (
            .O(N__47662),
            .I(N__47659));
    Odrv4 I__8779 (
            .O(N__47659),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n712 ));
    InMux I__8778 (
            .O(N__47656),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17639 ));
    InMux I__8777 (
            .O(N__47653),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382 ));
    InMux I__8776 (
            .O(N__47650),
            .I(N__47647));
    LocalMux I__8775 (
            .O(N__47647),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n93 ));
    InMux I__8774 (
            .O(N__47644),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17927 ));
    InMux I__8773 (
            .O(N__47641),
            .I(N__47638));
    LocalMux I__8772 (
            .O(N__47638),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414 ));
    InMux I__8771 (
            .O(N__47635),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17928 ));
    CascadeMux I__8770 (
            .O(N__47632),
            .I(N__47629));
    InMux I__8769 (
            .O(N__47629),
            .I(N__47626));
    LocalMux I__8768 (
            .O(N__47626),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n191 ));
    InMux I__8767 (
            .O(N__47623),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17929 ));
    CascadeMux I__8766 (
            .O(N__47620),
            .I(N__47617));
    InMux I__8765 (
            .O(N__47617),
            .I(N__47614));
    LocalMux I__8764 (
            .O(N__47614),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n240 ));
    InMux I__8763 (
            .O(N__47611),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17930 ));
    InMux I__8762 (
            .O(N__47608),
            .I(N__47605));
    LocalMux I__8761 (
            .O(N__47605),
            .I(N__47602));
    Odrv4 I__8760 (
            .O(N__47602),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n222 ));
    InMux I__8759 (
            .O(N__47599),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17629 ));
    CascadeMux I__8758 (
            .O(N__47596),
            .I(N__47593));
    InMux I__8757 (
            .O(N__47593),
            .I(N__47590));
    LocalMux I__8756 (
            .O(N__47590),
            .I(N__47587));
    Odrv4 I__8755 (
            .O(N__47587),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n271 ));
    InMux I__8754 (
            .O(N__47584),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17630 ));
    CascadeMux I__8753 (
            .O(N__47581),
            .I(N__47578));
    InMux I__8752 (
            .O(N__47578),
            .I(N__47575));
    LocalMux I__8751 (
            .O(N__47575),
            .I(N__47572));
    Odrv4 I__8750 (
            .O(N__47572),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n320 ));
    InMux I__8749 (
            .O(N__47569),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17631 ));
    InMux I__8748 (
            .O(N__47566),
            .I(N__47563));
    LocalMux I__8747 (
            .O(N__47563),
            .I(N__47560));
    Odrv4 I__8746 (
            .O(N__47560),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n369 ));
    InMux I__8745 (
            .O(N__47557),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17632 ));
    InMux I__8744 (
            .O(N__47554),
            .I(N__47551));
    LocalMux I__8743 (
            .O(N__47551),
            .I(N__47548));
    Odrv4 I__8742 (
            .O(N__47548),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n418 ));
    InMux I__8741 (
            .O(N__47545),
            .I(bfn_19_8_0_));
    CascadeMux I__8740 (
            .O(N__47542),
            .I(N__47539));
    InMux I__8739 (
            .O(N__47539),
            .I(N__47536));
    LocalMux I__8738 (
            .O(N__47536),
            .I(N__47533));
    Odrv12 I__8737 (
            .O(N__47533),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n467 ));
    InMux I__8736 (
            .O(N__47530),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17634 ));
    InMux I__8735 (
            .O(N__47527),
            .I(N__47524));
    LocalMux I__8734 (
            .O(N__47524),
            .I(N__47521));
    Odrv4 I__8733 (
            .O(N__47521),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n516 ));
    InMux I__8732 (
            .O(N__47518),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17635 ));
    CascadeMux I__8731 (
            .O(N__47515),
            .I(N__47512));
    InMux I__8730 (
            .O(N__47512),
            .I(N__47509));
    LocalMux I__8729 (
            .O(N__47509),
            .I(N__47506));
    Odrv12 I__8728 (
            .O(N__47506),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n565 ));
    InMux I__8727 (
            .O(N__47503),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17636 ));
    InMux I__8726 (
            .O(N__47500),
            .I(N__47497));
    LocalMux I__8725 (
            .O(N__47497),
            .I(N__47494));
    Odrv4 I__8724 (
            .O(N__47494),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n614 ));
    InMux I__8723 (
            .O(N__47491),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17637 ));
    InMux I__8722 (
            .O(N__47488),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17651 ));
    InMux I__8721 (
            .O(N__47485),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17652 ));
    InMux I__8720 (
            .O(N__47482),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17653 ));
    CascadeMux I__8719 (
            .O(N__47479),
            .I(N__47476));
    InMux I__8718 (
            .O(N__47476),
            .I(N__47473));
    LocalMux I__8717 (
            .O(N__47473),
            .I(N__47469));
    InMux I__8716 (
            .O(N__47472),
            .I(N__47466));
    Span4Mux_v I__8715 (
            .O(N__47469),
            .I(N__47463));
    LocalMux I__8714 (
            .O(N__47466),
            .I(N__47460));
    Odrv4 I__8713 (
            .O(N__47463),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n769 ));
    Odrv12 I__8712 (
            .O(N__47460),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n769 ));
    InMux I__8711 (
            .O(N__47455),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17654 ));
    InMux I__8710 (
            .O(N__47452),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n771 ));
    CascadeMux I__8709 (
            .O(N__47449),
            .I(N__47446));
    InMux I__8708 (
            .O(N__47446),
            .I(N__47443));
    LocalMux I__8707 (
            .O(N__47443),
            .I(N__47440));
    Odrv4 I__8706 (
            .O(N__47440),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510 ));
    InMux I__8705 (
            .O(N__47437),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17626 ));
    InMux I__8704 (
            .O(N__47434),
            .I(N__47431));
    LocalMux I__8703 (
            .O(N__47431),
            .I(N__47428));
    Odrv4 I__8702 (
            .O(N__47428),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n124 ));
    InMux I__8701 (
            .O(N__47425),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17627 ));
    CascadeMux I__8700 (
            .O(N__47422),
            .I(N__47419));
    InMux I__8699 (
            .O(N__47419),
            .I(N__47416));
    LocalMux I__8698 (
            .O(N__47416),
            .I(N__47413));
    Odrv12 I__8697 (
            .O(N__47413),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n173 ));
    InMux I__8696 (
            .O(N__47410),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17628 ));
    InMux I__8695 (
            .O(N__47407),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17642 ));
    InMux I__8694 (
            .O(N__47404),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17643 ));
    InMux I__8693 (
            .O(N__47401),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17644 ));
    InMux I__8692 (
            .O(N__47398),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17645 ));
    InMux I__8691 (
            .O(N__47395),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17646 ));
    InMux I__8690 (
            .O(N__47392),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17647 ));
    InMux I__8689 (
            .O(N__47389),
            .I(bfn_19_6_0_));
    InMux I__8688 (
            .O(N__47386),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17649 ));
    InMux I__8687 (
            .O(N__47383),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17650 ));
    InMux I__8686 (
            .O(N__47380),
            .I(N__47377));
    LocalMux I__8685 (
            .O(N__47377),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n534 ));
    InMux I__8684 (
            .O(N__47374),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18363 ));
    InMux I__8683 (
            .O(N__47371),
            .I(N__47368));
    LocalMux I__8682 (
            .O(N__47368),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n583 ));
    InMux I__8681 (
            .O(N__47365),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18364 ));
    InMux I__8680 (
            .O(N__47362),
            .I(N__47359));
    LocalMux I__8679 (
            .O(N__47359),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n632 ));
    InMux I__8678 (
            .O(N__47356),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18365 ));
    CascadeMux I__8677 (
            .O(N__47353),
            .I(N__47350));
    InMux I__8676 (
            .O(N__47350),
            .I(N__47347));
    LocalMux I__8675 (
            .O(N__47347),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n681 ));
    InMux I__8674 (
            .O(N__47344),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18366 ));
    InMux I__8673 (
            .O(N__47341),
            .I(N__47338));
    LocalMux I__8672 (
            .O(N__47338),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n730 ));
    InMux I__8671 (
            .O(N__47335),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18367 ));
    InMux I__8670 (
            .O(N__47332),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791 ));
    InMux I__8669 (
            .O(N__47329),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17641 ));
    CascadeMux I__8668 (
            .O(N__47326),
            .I(N__47323));
    InMux I__8667 (
            .O(N__47323),
            .I(N__47320));
    LocalMux I__8666 (
            .O(N__47320),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n93 ));
    InMux I__8665 (
            .O(N__47317),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18354 ));
    CascadeMux I__8664 (
            .O(N__47314),
            .I(N__47311));
    InMux I__8663 (
            .O(N__47311),
            .I(N__47308));
    LocalMux I__8662 (
            .O(N__47308),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n142 ));
    InMux I__8661 (
            .O(N__47305),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18355 ));
    CascadeMux I__8660 (
            .O(N__47302),
            .I(N__47299));
    InMux I__8659 (
            .O(N__47299),
            .I(N__47296));
    LocalMux I__8658 (
            .O(N__47296),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n191 ));
    InMux I__8657 (
            .O(N__47293),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18356 ));
    InMux I__8656 (
            .O(N__47290),
            .I(N__47287));
    LocalMux I__8655 (
            .O(N__47287),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n240 ));
    InMux I__8654 (
            .O(N__47284),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18357 ));
    InMux I__8653 (
            .O(N__47281),
            .I(N__47278));
    LocalMux I__8652 (
            .O(N__47278),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n289 ));
    InMux I__8651 (
            .O(N__47275),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18358 ));
    InMux I__8650 (
            .O(N__47272),
            .I(N__47269));
    LocalMux I__8649 (
            .O(N__47269),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n338 ));
    InMux I__8648 (
            .O(N__47266),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18359 ));
    InMux I__8647 (
            .O(N__47263),
            .I(N__47260));
    LocalMux I__8646 (
            .O(N__47260),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n387 ));
    InMux I__8645 (
            .O(N__47257),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18360 ));
    InMux I__8644 (
            .O(N__47254),
            .I(N__47251));
    LocalMux I__8643 (
            .O(N__47251),
            .I(N__47248));
    Odrv4 I__8642 (
            .O(N__47248),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n436 ));
    InMux I__8641 (
            .O(N__47245),
            .I(bfn_18_27_0_));
    InMux I__8640 (
            .O(N__47242),
            .I(N__47239));
    LocalMux I__8639 (
            .O(N__47239),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n485 ));
    InMux I__8638 (
            .O(N__47236),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18362 ));
    CascadeMux I__8637 (
            .O(N__47233),
            .I(N__47230));
    InMux I__8636 (
            .O(N__47230),
            .I(N__47227));
    LocalMux I__8635 (
            .O(N__47227),
            .I(N__47224));
    Span12Mux_h I__8634 (
            .O(N__47224),
            .I(N__47221));
    Odrv12 I__8633 (
            .O(N__47221),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24 ));
    InMux I__8632 (
            .O(N__47218),
            .I(bfn_18_25_0_));
    InMux I__8631 (
            .O(N__47215),
            .I(N__47212));
    LocalMux I__8630 (
            .O(N__47212),
            .I(N__47209));
    Span12Mux_s9_v I__8629 (
            .O(N__47209),
            .I(N__47206));
    Odrv12 I__8628 (
            .O(N__47206),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25 ));
    InMux I__8627 (
            .O(N__47203),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15907 ));
    CascadeMux I__8626 (
            .O(N__47200),
            .I(N__47197));
    InMux I__8625 (
            .O(N__47197),
            .I(N__47194));
    LocalMux I__8624 (
            .O(N__47194),
            .I(N__47191));
    Span4Mux_v I__8623 (
            .O(N__47191),
            .I(N__47188));
    Sp12to4 I__8622 (
            .O(N__47188),
            .I(N__47185));
    Odrv12 I__8621 (
            .O(N__47185),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26 ));
    InMux I__8620 (
            .O(N__47182),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15908 ));
    InMux I__8619 (
            .O(N__47179),
            .I(N__47176));
    LocalMux I__8618 (
            .O(N__47176),
            .I(N__47173));
    Span4Mux_v I__8617 (
            .O(N__47173),
            .I(N__47170));
    Span4Mux_h I__8616 (
            .O(N__47170),
            .I(N__47167));
    Odrv4 I__8615 (
            .O(N__47167),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27 ));
    InMux I__8614 (
            .O(N__47164),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15909 ));
    CascadeMux I__8613 (
            .O(N__47161),
            .I(N__47158));
    InMux I__8612 (
            .O(N__47158),
            .I(N__47155));
    LocalMux I__8611 (
            .O(N__47155),
            .I(N__47152));
    Span4Mux_v I__8610 (
            .O(N__47152),
            .I(N__47149));
    Span4Mux_h I__8609 (
            .O(N__47149),
            .I(N__47146));
    Odrv4 I__8608 (
            .O(N__47146),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28 ));
    InMux I__8607 (
            .O(N__47143),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15910 ));
    InMux I__8606 (
            .O(N__47140),
            .I(N__47137));
    LocalMux I__8605 (
            .O(N__47137),
            .I(N__47134));
    Span4Mux_v I__8604 (
            .O(N__47134),
            .I(N__47131));
    Span4Mux_h I__8603 (
            .O(N__47131),
            .I(N__47128));
    Odrv4 I__8602 (
            .O(N__47128),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29 ));
    InMux I__8601 (
            .O(N__47125),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15911 ));
    InMux I__8600 (
            .O(N__47122),
            .I(N__47119));
    LocalMux I__8599 (
            .O(N__47119),
            .I(N__47116));
    Span4Mux_v I__8598 (
            .O(N__47116),
            .I(N__47113));
    Span4Mux_h I__8597 (
            .O(N__47113),
            .I(N__47110));
    Odrv4 I__8596 (
            .O(N__47110),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30 ));
    InMux I__8595 (
            .O(N__47107),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15912 ));
    CascadeMux I__8594 (
            .O(N__47104),
            .I(N__47101));
    InMux I__8593 (
            .O(N__47101),
            .I(N__47098));
    LocalMux I__8592 (
            .O(N__47098),
            .I(N__47095));
    Span12Mux_h I__8591 (
            .O(N__47095),
            .I(N__47092));
    Odrv12 I__8590 (
            .O(N__47092),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15 ));
    InMux I__8589 (
            .O(N__47089),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15897 ));
    InMux I__8588 (
            .O(N__47086),
            .I(N__47083));
    LocalMux I__8587 (
            .O(N__47083),
            .I(N__47080));
    Span12Mux_h I__8586 (
            .O(N__47080),
            .I(N__47077));
    Odrv12 I__8585 (
            .O(N__47077),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16 ));
    InMux I__8584 (
            .O(N__47074),
            .I(bfn_18_24_0_));
    CascadeMux I__8583 (
            .O(N__47071),
            .I(N__47068));
    InMux I__8582 (
            .O(N__47068),
            .I(N__47065));
    LocalMux I__8581 (
            .O(N__47065),
            .I(N__47062));
    Span4Mux_v I__8580 (
            .O(N__47062),
            .I(N__47059));
    Span4Mux_h I__8579 (
            .O(N__47059),
            .I(N__47056));
    Odrv4 I__8578 (
            .O(N__47056),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17 ));
    InMux I__8577 (
            .O(N__47053),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15899 ));
    CascadeMux I__8576 (
            .O(N__47050),
            .I(N__47047));
    InMux I__8575 (
            .O(N__47047),
            .I(N__47044));
    LocalMux I__8574 (
            .O(N__47044),
            .I(N__47041));
    Span4Mux_v I__8573 (
            .O(N__47041),
            .I(N__47038));
    Span4Mux_h I__8572 (
            .O(N__47038),
            .I(N__47035));
    Odrv4 I__8571 (
            .O(N__47035),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18 ));
    InMux I__8570 (
            .O(N__47032),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15900 ));
    InMux I__8569 (
            .O(N__47029),
            .I(N__47026));
    LocalMux I__8568 (
            .O(N__47026),
            .I(N__47023));
    Span4Mux_h I__8567 (
            .O(N__47023),
            .I(N__47020));
    Span4Mux_h I__8566 (
            .O(N__47020),
            .I(N__47017));
    Odrv4 I__8565 (
            .O(N__47017),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19 ));
    InMux I__8564 (
            .O(N__47014),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15901 ));
    CascadeMux I__8563 (
            .O(N__47011),
            .I(N__47008));
    InMux I__8562 (
            .O(N__47008),
            .I(N__47005));
    LocalMux I__8561 (
            .O(N__47005),
            .I(N__47002));
    Span4Mux_v I__8560 (
            .O(N__47002),
            .I(N__46999));
    Span4Mux_h I__8559 (
            .O(N__46999),
            .I(N__46996));
    Odrv4 I__8558 (
            .O(N__46996),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20 ));
    InMux I__8557 (
            .O(N__46993),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15902 ));
    CascadeMux I__8556 (
            .O(N__46990),
            .I(N__46987));
    InMux I__8555 (
            .O(N__46987),
            .I(N__46984));
    LocalMux I__8554 (
            .O(N__46984),
            .I(N__46981));
    Span4Mux_v I__8553 (
            .O(N__46981),
            .I(N__46978));
    Span4Mux_h I__8552 (
            .O(N__46978),
            .I(N__46975));
    Odrv4 I__8551 (
            .O(N__46975),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21 ));
    InMux I__8550 (
            .O(N__46972),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15903 ));
    CascadeMux I__8549 (
            .O(N__46969),
            .I(N__46966));
    InMux I__8548 (
            .O(N__46966),
            .I(N__46963));
    LocalMux I__8547 (
            .O(N__46963),
            .I(N__46960));
    Span4Mux_v I__8546 (
            .O(N__46960),
            .I(N__46957));
    Span4Mux_h I__8545 (
            .O(N__46957),
            .I(N__46954));
    Odrv4 I__8544 (
            .O(N__46954),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22 ));
    InMux I__8543 (
            .O(N__46951),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15904 ));
    CascadeMux I__8542 (
            .O(N__46948),
            .I(N__46945));
    InMux I__8541 (
            .O(N__46945),
            .I(N__46942));
    LocalMux I__8540 (
            .O(N__46942),
            .I(N__46939));
    Span4Mux_v I__8539 (
            .O(N__46939),
            .I(N__46936));
    Span4Mux_h I__8538 (
            .O(N__46936),
            .I(N__46933));
    Odrv4 I__8537 (
            .O(N__46933),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23 ));
    InMux I__8536 (
            .O(N__46930),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15905 ));
    CascadeMux I__8535 (
            .O(N__46927),
            .I(N__46924));
    InMux I__8534 (
            .O(N__46924),
            .I(N__46921));
    LocalMux I__8533 (
            .O(N__46921),
            .I(N__46918));
    Span4Mux_h I__8532 (
            .O(N__46918),
            .I(N__46915));
    Odrv4 I__8531 (
            .O(N__46915),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7 ));
    InMux I__8530 (
            .O(N__46912),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15889 ));
    CascadeMux I__8529 (
            .O(N__46909),
            .I(N__46906));
    InMux I__8528 (
            .O(N__46906),
            .I(N__46903));
    LocalMux I__8527 (
            .O(N__46903),
            .I(N__46900));
    Odrv4 I__8526 (
            .O(N__46900),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8 ));
    InMux I__8525 (
            .O(N__46897),
            .I(bfn_18_23_0_));
    CascadeMux I__8524 (
            .O(N__46894),
            .I(N__46891));
    InMux I__8523 (
            .O(N__46891),
            .I(N__46888));
    LocalMux I__8522 (
            .O(N__46888),
            .I(N__46885));
    Span4Mux_v I__8521 (
            .O(N__46885),
            .I(N__46882));
    Odrv4 I__8520 (
            .O(N__46882),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9 ));
    InMux I__8519 (
            .O(N__46879),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15891 ));
    CascadeMux I__8518 (
            .O(N__46876),
            .I(N__46873));
    InMux I__8517 (
            .O(N__46873),
            .I(N__46870));
    LocalMux I__8516 (
            .O(N__46870),
            .I(N__46867));
    Span4Mux_v I__8515 (
            .O(N__46867),
            .I(N__46864));
    Odrv4 I__8514 (
            .O(N__46864),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10 ));
    InMux I__8513 (
            .O(N__46861),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15892 ));
    CascadeMux I__8512 (
            .O(N__46858),
            .I(N__46855));
    InMux I__8511 (
            .O(N__46855),
            .I(N__46852));
    LocalMux I__8510 (
            .O(N__46852),
            .I(N__46849));
    Span4Mux_h I__8509 (
            .O(N__46849),
            .I(N__46846));
    Odrv4 I__8508 (
            .O(N__46846),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11 ));
    InMux I__8507 (
            .O(N__46843),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15893 ));
    CascadeMux I__8506 (
            .O(N__46840),
            .I(N__46837));
    InMux I__8505 (
            .O(N__46837),
            .I(N__46834));
    LocalMux I__8504 (
            .O(N__46834),
            .I(N__46831));
    Span4Mux_h I__8503 (
            .O(N__46831),
            .I(N__46828));
    Odrv4 I__8502 (
            .O(N__46828),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12 ));
    InMux I__8501 (
            .O(N__46825),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15894 ));
    CascadeMux I__8500 (
            .O(N__46822),
            .I(N__46819));
    InMux I__8499 (
            .O(N__46819),
            .I(N__46816));
    LocalMux I__8498 (
            .O(N__46816),
            .I(N__46813));
    Span4Mux_h I__8497 (
            .O(N__46813),
            .I(N__46810));
    Odrv4 I__8496 (
            .O(N__46810),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13 ));
    InMux I__8495 (
            .O(N__46807),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15895 ));
    InMux I__8494 (
            .O(N__46804),
            .I(N__46801));
    LocalMux I__8493 (
            .O(N__46801),
            .I(N__46798));
    Span4Mux_h I__8492 (
            .O(N__46798),
            .I(N__46795));
    Odrv4 I__8491 (
            .O(N__46795),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14 ));
    InMux I__8490 (
            .O(N__46792),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15896 ));
    InMux I__8489 (
            .O(N__46789),
            .I(N__46786));
    LocalMux I__8488 (
            .O(N__46786),
            .I(N__46782));
    InMux I__8487 (
            .O(N__46785),
            .I(N__46779));
    Odrv4 I__8486 (
            .O(N__46782),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28 ));
    LocalMux I__8485 (
            .O(N__46779),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28 ));
    InMux I__8484 (
            .O(N__46774),
            .I(N__46770));
    InMux I__8483 (
            .O(N__46773),
            .I(N__46767));
    LocalMux I__8482 (
            .O(N__46770),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20174 ));
    LocalMux I__8481 (
            .O(N__46767),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20174 ));
    CascadeMux I__8480 (
            .O(N__46762),
            .I(N__46759));
    InMux I__8479 (
            .O(N__46759),
            .I(N__46756));
    LocalMux I__8478 (
            .O(N__46756),
            .I(N__46753));
    Span4Mux_v I__8477 (
            .O(N__46753),
            .I(N__46750));
    Odrv4 I__8476 (
            .O(N__46750),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1 ));
    InMux I__8475 (
            .O(N__46747),
            .I(N__46743));
    InMux I__8474 (
            .O(N__46746),
            .I(N__46740));
    LocalMux I__8473 (
            .O(N__46743),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2 ));
    LocalMux I__8472 (
            .O(N__46740),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2 ));
    InMux I__8471 (
            .O(N__46735),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15883 ));
    CascadeMux I__8470 (
            .O(N__46732),
            .I(N__46729));
    InMux I__8469 (
            .O(N__46729),
            .I(N__46726));
    LocalMux I__8468 (
            .O(N__46726),
            .I(N__46723));
    Span4Mux_v I__8467 (
            .O(N__46723),
            .I(N__46720));
    Odrv4 I__8466 (
            .O(N__46720),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2 ));
    CascadeMux I__8465 (
            .O(N__46717),
            .I(N__46713));
    InMux I__8464 (
            .O(N__46716),
            .I(N__46710));
    InMux I__8463 (
            .O(N__46713),
            .I(N__46707));
    LocalMux I__8462 (
            .O(N__46710),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3 ));
    LocalMux I__8461 (
            .O(N__46707),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3 ));
    InMux I__8460 (
            .O(N__46702),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15884 ));
    InMux I__8459 (
            .O(N__46699),
            .I(N__46696));
    LocalMux I__8458 (
            .O(N__46696),
            .I(N__46693));
    Span4Mux_h I__8457 (
            .O(N__46693),
            .I(N__46690));
    Odrv4 I__8456 (
            .O(N__46690),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3 ));
    CascadeMux I__8455 (
            .O(N__46687),
            .I(N__46684));
    InMux I__8454 (
            .O(N__46684),
            .I(N__46680));
    InMux I__8453 (
            .O(N__46683),
            .I(N__46677));
    LocalMux I__8452 (
            .O(N__46680),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4 ));
    LocalMux I__8451 (
            .O(N__46677),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4 ));
    InMux I__8450 (
            .O(N__46672),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15885 ));
    CascadeMux I__8449 (
            .O(N__46669),
            .I(N__46666));
    InMux I__8448 (
            .O(N__46666),
            .I(N__46663));
    LocalMux I__8447 (
            .O(N__46663),
            .I(N__46660));
    Span4Mux_h I__8446 (
            .O(N__46660),
            .I(N__46657));
    Span4Mux_v I__8445 (
            .O(N__46657),
            .I(N__46654));
    Odrv4 I__8444 (
            .O(N__46654),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4 ));
    InMux I__8443 (
            .O(N__46651),
            .I(N__46647));
    InMux I__8442 (
            .O(N__46650),
            .I(N__46644));
    LocalMux I__8441 (
            .O(N__46647),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5 ));
    LocalMux I__8440 (
            .O(N__46644),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5 ));
    InMux I__8439 (
            .O(N__46639),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15886 ));
    CascadeMux I__8438 (
            .O(N__46636),
            .I(N__46633));
    InMux I__8437 (
            .O(N__46633),
            .I(N__46630));
    LocalMux I__8436 (
            .O(N__46630),
            .I(N__46627));
    Span4Mux_h I__8435 (
            .O(N__46627),
            .I(N__46624));
    Odrv4 I__8434 (
            .O(N__46624),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5 ));
    InMux I__8433 (
            .O(N__46621),
            .I(N__46617));
    InMux I__8432 (
            .O(N__46620),
            .I(N__46614));
    LocalMux I__8431 (
            .O(N__46617),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6 ));
    LocalMux I__8430 (
            .O(N__46614),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6 ));
    InMux I__8429 (
            .O(N__46609),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15887 ));
    CascadeMux I__8428 (
            .O(N__46606),
            .I(N__46603));
    InMux I__8427 (
            .O(N__46603),
            .I(N__46600));
    LocalMux I__8426 (
            .O(N__46600),
            .I(N__46597));
    Span4Mux_h I__8425 (
            .O(N__46597),
            .I(N__46594));
    Odrv4 I__8424 (
            .O(N__46594),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6 ));
    InMux I__8423 (
            .O(N__46591),
            .I(N__46587));
    InMux I__8422 (
            .O(N__46590),
            .I(N__46584));
    LocalMux I__8421 (
            .O(N__46587),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7 ));
    LocalMux I__8420 (
            .O(N__46584),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7 ));
    InMux I__8419 (
            .O(N__46579),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15888 ));
    CascadeMux I__8418 (
            .O(N__46576),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_ ));
    InMux I__8417 (
            .O(N__46573),
            .I(N__46569));
    InMux I__8416 (
            .O(N__46572),
            .I(N__46566));
    LocalMux I__8415 (
            .O(N__46569),
            .I(N__46563));
    LocalMux I__8414 (
            .O(N__46566),
            .I(N__46560));
    Odrv4 I__8413 (
            .O(N__46563),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24 ));
    Odrv4 I__8412 (
            .O(N__46560),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24 ));
    InMux I__8411 (
            .O(N__46555),
            .I(N__46551));
    InMux I__8410 (
            .O(N__46554),
            .I(N__46548));
    LocalMux I__8409 (
            .O(N__46551),
            .I(N__46545));
    LocalMux I__8408 (
            .O(N__46548),
            .I(N__46542));
    Odrv12 I__8407 (
            .O(N__46545),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26 ));
    Odrv12 I__8406 (
            .O(N__46542),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26 ));
    InMux I__8405 (
            .O(N__46537),
            .I(N__46534));
    LocalMux I__8404 (
            .O(N__46534),
            .I(N__46531));
    Odrv4 I__8403 (
            .O(N__46531),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102 ));
    CascadeMux I__8402 (
            .O(N__46528),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_ ));
    InMux I__8401 (
            .O(N__46525),
            .I(N__46522));
    LocalMux I__8400 (
            .O(N__46522),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890 ));
    InMux I__8399 (
            .O(N__46519),
            .I(N__46515));
    InMux I__8398 (
            .O(N__46518),
            .I(N__46512));
    LocalMux I__8397 (
            .O(N__46515),
            .I(N__46509));
    LocalMux I__8396 (
            .O(N__46512),
            .I(N__46506));
    Span4Mux_v I__8395 (
            .O(N__46509),
            .I(N__46503));
    Odrv4 I__8394 (
            .O(N__46506),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21 ));
    Odrv4 I__8393 (
            .O(N__46503),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21 ));
    CascadeMux I__8392 (
            .O(N__46498),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_ ));
    InMux I__8391 (
            .O(N__46495),
            .I(N__46492));
    LocalMux I__8390 (
            .O(N__46492),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362 ));
    InMux I__8389 (
            .O(N__46489),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17759 ));
    InMux I__8388 (
            .O(N__46486),
            .I(N__46483));
    LocalMux I__8387 (
            .O(N__46483),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n501 ));
    InMux I__8386 (
            .O(N__46480),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17760 ));
    InMux I__8385 (
            .O(N__46477),
            .I(N__46474));
    LocalMux I__8384 (
            .O(N__46474),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n550 ));
    InMux I__8383 (
            .O(N__46471),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17761 ));
    InMux I__8382 (
            .O(N__46468),
            .I(N__46465));
    LocalMux I__8381 (
            .O(N__46465),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n599 ));
    InMux I__8380 (
            .O(N__46462),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17762 ));
    CascadeMux I__8379 (
            .O(N__46459),
            .I(N__46456));
    InMux I__8378 (
            .O(N__46456),
            .I(N__46453));
    LocalMux I__8377 (
            .O(N__46453),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347 ));
    InMux I__8376 (
            .O(N__46450),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17763 ));
    CascadeMux I__8375 (
            .O(N__46447),
            .I(N__46444));
    InMux I__8374 (
            .O(N__46444),
            .I(N__46441));
    LocalMux I__8373 (
            .O(N__46441),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n697 ));
    InMux I__8372 (
            .O(N__46438),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17764 ));
    InMux I__8371 (
            .O(N__46435),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n747 ));
    InMux I__8370 (
            .O(N__46432),
            .I(N__46429));
    LocalMux I__8369 (
            .O(N__46429),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108 ));
    CascadeMux I__8368 (
            .O(N__46426),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_ ));
    InMux I__8367 (
            .O(N__46423),
            .I(N__46420));
    LocalMux I__8366 (
            .O(N__46420),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n60 ));
    InMux I__8365 (
            .O(N__46417),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17751 ));
    InMux I__8364 (
            .O(N__46414),
            .I(N__46411));
    LocalMux I__8363 (
            .O(N__46411),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383 ));
    InMux I__8362 (
            .O(N__46408),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17752 ));
    CascadeMux I__8361 (
            .O(N__46405),
            .I(N__46402));
    InMux I__8360 (
            .O(N__46402),
            .I(N__46399));
    LocalMux I__8359 (
            .O(N__46399),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375 ));
    InMux I__8358 (
            .O(N__46396),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17753 ));
    InMux I__8357 (
            .O(N__46393),
            .I(N__46390));
    LocalMux I__8356 (
            .O(N__46390),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n207 ));
    InMux I__8355 (
            .O(N__46387),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17754 ));
    InMux I__8354 (
            .O(N__46384),
            .I(N__46381));
    LocalMux I__8353 (
            .O(N__46381),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n256 ));
    InMux I__8352 (
            .O(N__46378),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17755 ));
    InMux I__8351 (
            .O(N__46375),
            .I(N__46372));
    LocalMux I__8350 (
            .O(N__46372),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n305 ));
    InMux I__8349 (
            .O(N__46369),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17756 ));
    CascadeMux I__8348 (
            .O(N__46366),
            .I(N__46363));
    InMux I__8347 (
            .O(N__46363),
            .I(N__46360));
    LocalMux I__8346 (
            .O(N__46360),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367 ));
    InMux I__8345 (
            .O(N__46357),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17757 ));
    InMux I__8344 (
            .O(N__46354),
            .I(N__46351));
    LocalMux I__8343 (
            .O(N__46351),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365 ));
    InMux I__8342 (
            .O(N__46348),
            .I(bfn_18_19_0_));
    InMux I__8341 (
            .O(N__46345),
            .I(N__46342));
    LocalMux I__8340 (
            .O(N__46342),
            .I(N__46339));
    Odrv12 I__8339 (
            .O(N__46339),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500 ));
    InMux I__8338 (
            .O(N__46336),
            .I(bfn_18_17_0_));
    InMux I__8337 (
            .O(N__46333),
            .I(N__46330));
    LocalMux I__8336 (
            .O(N__46330),
            .I(N__46327));
    Odrv4 I__8335 (
            .O(N__46327),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499 ));
    InMux I__8334 (
            .O(N__46324),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17834 ));
    InMux I__8333 (
            .O(N__46321),
            .I(N__46318));
    LocalMux I__8332 (
            .O(N__46318),
            .I(N__46315));
    Odrv4 I__8331 (
            .O(N__46315),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498 ));
    InMux I__8330 (
            .O(N__46312),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17835 ));
    InMux I__8329 (
            .O(N__46309),
            .I(N__46306));
    LocalMux I__8328 (
            .O(N__46306),
            .I(N__46303));
    Odrv12 I__8327 (
            .O(N__46303),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497 ));
    InMux I__8326 (
            .O(N__46300),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17836 ));
    InMux I__8325 (
            .O(N__46297),
            .I(N__46294));
    LocalMux I__8324 (
            .O(N__46294),
            .I(N__46291));
    Odrv4 I__8323 (
            .O(N__46291),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496 ));
    InMux I__8322 (
            .O(N__46288),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17837 ));
    InMux I__8321 (
            .O(N__46285),
            .I(N__46282));
    LocalMux I__8320 (
            .O(N__46282),
            .I(N__46279));
    Odrv4 I__8319 (
            .O(N__46279),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494 ));
    InMux I__8318 (
            .O(N__46276),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17838 ));
    CascadeMux I__8317 (
            .O(N__46273),
            .I(N__46270));
    InMux I__8316 (
            .O(N__46270),
            .I(N__46267));
    LocalMux I__8315 (
            .O(N__46267),
            .I(N__46264));
    Odrv4 I__8314 (
            .O(N__46264),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493 ));
    InMux I__8313 (
            .O(N__46261),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17839 ));
    InMux I__8312 (
            .O(N__46258),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n767 ));
    InMux I__8311 (
            .O(N__46255),
            .I(N__46252));
    LocalMux I__8310 (
            .O(N__46252),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n75 ));
    InMux I__8309 (
            .O(N__46249),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17826 ));
    InMux I__8308 (
            .O(N__46246),
            .I(N__46243));
    LocalMux I__8307 (
            .O(N__46243),
            .I(N__46240));
    Odrv4 I__8306 (
            .O(N__46240),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507 ));
    InMux I__8305 (
            .O(N__46237),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17827 ));
    InMux I__8304 (
            .O(N__46234),
            .I(N__46231));
    LocalMux I__8303 (
            .O(N__46231),
            .I(N__46228));
    Odrv12 I__8302 (
            .O(N__46228),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506 ));
    InMux I__8301 (
            .O(N__46225),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17828 ));
    InMux I__8300 (
            .O(N__46222),
            .I(N__46219));
    LocalMux I__8299 (
            .O(N__46219),
            .I(N__46216));
    Odrv4 I__8298 (
            .O(N__46216),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505 ));
    InMux I__8297 (
            .O(N__46213),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17829 ));
    InMux I__8296 (
            .O(N__46210),
            .I(N__46207));
    LocalMux I__8295 (
            .O(N__46207),
            .I(N__46204));
    Odrv4 I__8294 (
            .O(N__46204),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503 ));
    InMux I__8293 (
            .O(N__46201),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17830 ));
    InMux I__8292 (
            .O(N__46198),
            .I(N__46195));
    LocalMux I__8291 (
            .O(N__46195),
            .I(N__46192));
    Odrv12 I__8290 (
            .O(N__46192),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502 ));
    InMux I__8289 (
            .O(N__46189),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17831 ));
    CascadeMux I__8288 (
            .O(N__46186),
            .I(N__46183));
    InMux I__8287 (
            .O(N__46183),
            .I(N__46180));
    LocalMux I__8286 (
            .O(N__46180),
            .I(N__46177));
    Odrv4 I__8285 (
            .O(N__46177),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501 ));
    InMux I__8284 (
            .O(N__46174),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17832 ));
    InMux I__8283 (
            .O(N__46171),
            .I(N__46168));
    LocalMux I__8282 (
            .O(N__46168),
            .I(N__46165));
    Odrv4 I__8281 (
            .O(N__46165),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473 ));
    InMux I__8280 (
            .O(N__46162),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17847 ));
    InMux I__8279 (
            .O(N__46159),
            .I(N__46156));
    LocalMux I__8278 (
            .O(N__46156),
            .I(N__46153));
    Odrv4 I__8277 (
            .O(N__46153),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465 ));
    InMux I__8276 (
            .O(N__46150),
            .I(bfn_18_15_0_));
    InMux I__8275 (
            .O(N__46147),
            .I(N__46144));
    LocalMux I__8274 (
            .O(N__46144),
            .I(N__46141));
    Odrv4 I__8273 (
            .O(N__46141),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463 ));
    InMux I__8272 (
            .O(N__46138),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17849 ));
    InMux I__8271 (
            .O(N__46135),
            .I(N__46132));
    LocalMux I__8270 (
            .O(N__46132),
            .I(N__46129));
    Odrv4 I__8269 (
            .O(N__46129),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461 ));
    InMux I__8268 (
            .O(N__46126),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17850 ));
    InMux I__8267 (
            .O(N__46123),
            .I(N__46120));
    LocalMux I__8266 (
            .O(N__46120),
            .I(N__46117));
    Odrv12 I__8265 (
            .O(N__46117),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460 ));
    InMux I__8264 (
            .O(N__46114),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17851 ));
    InMux I__8263 (
            .O(N__46111),
            .I(N__46108));
    LocalMux I__8262 (
            .O(N__46108),
            .I(N__46105));
    Odrv12 I__8261 (
            .O(N__46105),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459 ));
    InMux I__8260 (
            .O(N__46102),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17852 ));
    CascadeMux I__8259 (
            .O(N__46099),
            .I(N__46096));
    InMux I__8258 (
            .O(N__46096),
            .I(N__46093));
    LocalMux I__8257 (
            .O(N__46093),
            .I(N__46090));
    Span4Mux_v I__8256 (
            .O(N__46090),
            .I(N__46087));
    Odrv4 I__8255 (
            .O(N__46087),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n666 ));
    InMux I__8254 (
            .O(N__46084),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17853 ));
    CascadeMux I__8253 (
            .O(N__46081),
            .I(N__46078));
    InMux I__8252 (
            .O(N__46078),
            .I(N__46075));
    LocalMux I__8251 (
            .O(N__46075),
            .I(N__46072));
    Odrv4 I__8250 (
            .O(N__46072),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n715 ));
    InMux I__8249 (
            .O(N__46069),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17854 ));
    InMux I__8248 (
            .O(N__46066),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353 ));
    InMux I__8247 (
            .O(N__46063),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17880 ));
    InMux I__8246 (
            .O(N__46060),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n775 ));
    InMux I__8245 (
            .O(N__46057),
            .I(N__46054));
    LocalMux I__8244 (
            .O(N__46054),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480 ));
    InMux I__8243 (
            .O(N__46051),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17841 ));
    InMux I__8242 (
            .O(N__46048),
            .I(N__46045));
    LocalMux I__8241 (
            .O(N__46045),
            .I(N__46042));
    Odrv4 I__8240 (
            .O(N__46042),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479 ));
    InMux I__8239 (
            .O(N__46039),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17842 ));
    InMux I__8238 (
            .O(N__46036),
            .I(N__46033));
    LocalMux I__8237 (
            .O(N__46033),
            .I(N__46030));
    Odrv4 I__8236 (
            .O(N__46030),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478 ));
    InMux I__8235 (
            .O(N__46027),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17843 ));
    InMux I__8234 (
            .O(N__46024),
            .I(N__46021));
    LocalMux I__8233 (
            .O(N__46021),
            .I(N__46018));
    Odrv12 I__8232 (
            .O(N__46018),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477 ));
    InMux I__8231 (
            .O(N__46015),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17844 ));
    InMux I__8230 (
            .O(N__46012),
            .I(N__46009));
    LocalMux I__8229 (
            .O(N__46009),
            .I(N__46006));
    Odrv4 I__8228 (
            .O(N__46006),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476 ));
    InMux I__8227 (
            .O(N__46003),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17845 ));
    CascadeMux I__8226 (
            .O(N__46000),
            .I(N__45997));
    InMux I__8225 (
            .O(N__45997),
            .I(N__45994));
    LocalMux I__8224 (
            .O(N__45994),
            .I(N__45991));
    Odrv4 I__8223 (
            .O(N__45991),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475 ));
    InMux I__8222 (
            .O(N__45988),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17846 ));
    CascadeMux I__8221 (
            .O(N__45985),
            .I(N__45982));
    InMux I__8220 (
            .O(N__45982),
            .I(N__45979));
    LocalMux I__8219 (
            .O(N__45979),
            .I(N__45976));
    Odrv4 I__8218 (
            .O(N__45976),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443 ));
    InMux I__8217 (
            .O(N__45973),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17872 ));
    InMux I__8216 (
            .O(N__45970),
            .I(N__45967));
    LocalMux I__8215 (
            .O(N__45967),
            .I(N__45964));
    Odrv4 I__8214 (
            .O(N__45964),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438 ));
    InMux I__8213 (
            .O(N__45961),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17873 ));
    InMux I__8212 (
            .O(N__45958),
            .I(N__45955));
    LocalMux I__8211 (
            .O(N__45955),
            .I(N__45952));
    Odrv4 I__8210 (
            .O(N__45952),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435 ));
    InMux I__8209 (
            .O(N__45949),
            .I(bfn_18_13_0_));
    InMux I__8208 (
            .O(N__45946),
            .I(N__45943));
    LocalMux I__8207 (
            .O(N__45943),
            .I(N__45940));
    Odrv4 I__8206 (
            .O(N__45940),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431 ));
    InMux I__8205 (
            .O(N__45937),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17875 ));
    InMux I__8204 (
            .O(N__45934),
            .I(N__45931));
    LocalMux I__8203 (
            .O(N__45931),
            .I(N__45928));
    Odrv4 I__8202 (
            .O(N__45928),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430 ));
    InMux I__8201 (
            .O(N__45925),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17876 ));
    InMux I__8200 (
            .O(N__45922),
            .I(N__45919));
    LocalMux I__8199 (
            .O(N__45919),
            .I(N__45916));
    Odrv12 I__8198 (
            .O(N__45916),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n571 ));
    InMux I__8197 (
            .O(N__45913),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17877 ));
    InMux I__8196 (
            .O(N__45910),
            .I(N__45907));
    LocalMux I__8195 (
            .O(N__45907),
            .I(N__45904));
    Odrv4 I__8194 (
            .O(N__45904),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n620 ));
    InMux I__8193 (
            .O(N__45901),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17878 ));
    CascadeMux I__8192 (
            .O(N__45898),
            .I(N__45895));
    InMux I__8191 (
            .O(N__45895),
            .I(N__45892));
    LocalMux I__8190 (
            .O(N__45892),
            .I(N__45889));
    Span4Mux_v I__8189 (
            .O(N__45889),
            .I(N__45886));
    Odrv4 I__8188 (
            .O(N__45886),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n669 ));
    InMux I__8187 (
            .O(N__45883),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17879 ));
    InMux I__8186 (
            .O(N__45880),
            .I(N__45877));
    LocalMux I__8185 (
            .O(N__45877),
            .I(N__45874));
    Odrv12 I__8184 (
            .O(N__45874),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n718 ));
    InMux I__8183 (
            .O(N__45871),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17894 ));
    InMux I__8182 (
            .O(N__45868),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17895 ));
    InMux I__8181 (
            .O(N__45865),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n779 ));
    InMux I__8180 (
            .O(N__45862),
            .I(N__45859));
    LocalMux I__8179 (
            .O(N__45859),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457 ));
    InMux I__8178 (
            .O(N__45856),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17867 ));
    InMux I__8177 (
            .O(N__45853),
            .I(N__45850));
    LocalMux I__8176 (
            .O(N__45850),
            .I(N__45847));
    Odrv4 I__8175 (
            .O(N__45847),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453 ));
    InMux I__8174 (
            .O(N__45844),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17868 ));
    InMux I__8173 (
            .O(N__45841),
            .I(N__45838));
    LocalMux I__8172 (
            .O(N__45838),
            .I(N__45835));
    Odrv12 I__8171 (
            .O(N__45835),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452 ));
    InMux I__8170 (
            .O(N__45832),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17869 ));
    InMux I__8169 (
            .O(N__45829),
            .I(N__45826));
    LocalMux I__8168 (
            .O(N__45826),
            .I(N__45823));
    Odrv4 I__8167 (
            .O(N__45823),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450 ));
    InMux I__8166 (
            .O(N__45820),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17870 ));
    InMux I__8165 (
            .O(N__45817),
            .I(N__45814));
    LocalMux I__8164 (
            .O(N__45814),
            .I(N__45811));
    Odrv4 I__8163 (
            .O(N__45811),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448 ));
    InMux I__8162 (
            .O(N__45808),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17871 ));
    InMux I__8161 (
            .O(N__45805),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17885 ));
    InMux I__8160 (
            .O(N__45802),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17886 ));
    InMux I__8159 (
            .O(N__45799),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17887 ));
    InMux I__8158 (
            .O(N__45796),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17888 ));
    InMux I__8157 (
            .O(N__45793),
            .I(bfn_18_11_0_));
    InMux I__8156 (
            .O(N__45790),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17890 ));
    InMux I__8155 (
            .O(N__45787),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17891 ));
    InMux I__8154 (
            .O(N__45784),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17892 ));
    InMux I__8153 (
            .O(N__45781),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17893 ));
    InMux I__8152 (
            .O(N__45778),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17952 ));
    CascadeMux I__8151 (
            .O(N__45775),
            .I(N__45771));
    InMux I__8150 (
            .O(N__45774),
            .I(N__45768));
    InMux I__8149 (
            .O(N__45771),
            .I(N__45765));
    LocalMux I__8148 (
            .O(N__45768),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n785 ));
    LocalMux I__8147 (
            .O(N__45765),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n785 ));
    InMux I__8146 (
            .O(N__45760),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17953 ));
    CascadeMux I__8145 (
            .O(N__45757),
            .I(N__45752));
    InMux I__8144 (
            .O(N__45756),
            .I(N__45749));
    InMux I__8143 (
            .O(N__45755),
            .I(N__45746));
    InMux I__8142 (
            .O(N__45752),
            .I(N__45743));
    LocalMux I__8141 (
            .O(N__45749),
            .I(N__45738));
    LocalMux I__8140 (
            .O(N__45746),
            .I(N__45738));
    LocalMux I__8139 (
            .O(N__45743),
            .I(N__45735));
    Odrv4 I__8138 (
            .O(N__45738),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n789 ));
    Odrv4 I__8137 (
            .O(N__45735),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n789 ));
    InMux I__8136 (
            .O(N__45730),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17954 ));
    InMux I__8135 (
            .O(N__45727),
            .I(N__45724));
    LocalMux I__8134 (
            .O(N__45724),
            .I(n793));
    InMux I__8133 (
            .O(N__45721),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17955 ));
    InMux I__8132 (
            .O(N__45718),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n795 ));
    CascadeMux I__8131 (
            .O(N__45715),
            .I(N__45712));
    InMux I__8130 (
            .O(N__45712),
            .I(N__45709));
    LocalMux I__8129 (
            .O(N__45709),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389 ));
    InMux I__8128 (
            .O(N__45706),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17882 ));
    InMux I__8127 (
            .O(N__45703),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17883 ));
    InMux I__8126 (
            .O(N__45700),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17884 ));
    InMux I__8125 (
            .O(N__45697),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17944 ));
    InMux I__8124 (
            .O(N__45694),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17945 ));
    InMux I__8123 (
            .O(N__45691),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17946 ));
    InMux I__8122 (
            .O(N__45688),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17947 ));
    InMux I__8121 (
            .O(N__45685),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17948 ));
    InMux I__8120 (
            .O(N__45682),
            .I(bfn_18_9_0_));
    InMux I__8119 (
            .O(N__45679),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17950 ));
    InMux I__8118 (
            .O(N__45676),
            .I(N__45673));
    LocalMux I__8117 (
            .O(N__45673),
            .I(N__45669));
    InMux I__8116 (
            .O(N__45672),
            .I(N__45666));
    Odrv4 I__8115 (
            .O(N__45669),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n777 ));
    LocalMux I__8114 (
            .O(N__45666),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n777 ));
    InMux I__8113 (
            .O(N__45661),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17951 ));
    InMux I__8112 (
            .O(N__45658),
            .I(N__45655));
    LocalMux I__8111 (
            .O(N__45655),
            .I(N__45651));
    InMux I__8110 (
            .O(N__45654),
            .I(N__45648));
    Odrv4 I__8109 (
            .O(N__45651),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n781 ));
    LocalMux I__8108 (
            .O(N__45648),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n781 ));
    InMux I__8107 (
            .O(N__45643),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17274 ));
    CascadeMux I__8106 (
            .O(N__45640),
            .I(N__45636));
    CascadeMux I__8105 (
            .O(N__45639),
            .I(N__45633));
    InMux I__8104 (
            .O(N__45636),
            .I(N__45629));
    InMux I__8103 (
            .O(N__45633),
            .I(N__45624));
    InMux I__8102 (
            .O(N__45632),
            .I(N__45624));
    LocalMux I__8101 (
            .O(N__45629),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n427 ));
    LocalMux I__8100 (
            .O(N__45624),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n427 ));
    InMux I__8099 (
            .O(N__45619),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17275 ));
    InMux I__8098 (
            .O(N__45616),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352 ));
    InMux I__8097 (
            .O(N__45613),
            .I(N__45610));
    LocalMux I__8096 (
            .O(N__45610),
            .I(N__45606));
    InMux I__8095 (
            .O(N__45609),
            .I(N__45603));
    Span4Mux_v I__8094 (
            .O(N__45606),
            .I(N__45598));
    LocalMux I__8093 (
            .O(N__45603),
            .I(N__45598));
    Odrv4 I__8092 (
            .O(N__45598),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23 ));
    InMux I__8091 (
            .O(N__45595),
            .I(N__45589));
    InMux I__8090 (
            .O(N__45594),
            .I(N__45589));
    LocalMux I__8089 (
            .O(N__45589),
            .I(N__45586));
    Odrv12 I__8088 (
            .O(N__45586),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19 ));
    InMux I__8087 (
            .O(N__45583),
            .I(N__45579));
    InMux I__8086 (
            .O(N__45582),
            .I(N__45576));
    LocalMux I__8085 (
            .O(N__45579),
            .I(N__45571));
    LocalMux I__8084 (
            .O(N__45576),
            .I(N__45571));
    Odrv4 I__8083 (
            .O(N__45571),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22 ));
    InMux I__8082 (
            .O(N__45568),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17942 ));
    InMux I__8081 (
            .O(N__45565),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17943 ));
    CascadeMux I__8080 (
            .O(N__45562),
            .I(N__45559));
    InMux I__8079 (
            .O(N__45559),
            .I(N__45556));
    LocalMux I__8078 (
            .O(N__45556),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n84 ));
    InMux I__8077 (
            .O(N__45553),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17266 ));
    InMux I__8076 (
            .O(N__45550),
            .I(N__45547));
    LocalMux I__8075 (
            .O(N__45547),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n133 ));
    InMux I__8074 (
            .O(N__45544),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17267 ));
    CascadeMux I__8073 (
            .O(N__45541),
            .I(N__45538));
    InMux I__8072 (
            .O(N__45538),
            .I(N__45535));
    LocalMux I__8071 (
            .O(N__45535),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n182 ));
    InMux I__8070 (
            .O(N__45532),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17268 ));
    InMux I__8069 (
            .O(N__45529),
            .I(N__45526));
    LocalMux I__8068 (
            .O(N__45526),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n231 ));
    InMux I__8067 (
            .O(N__45523),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17269 ));
    CascadeMux I__8066 (
            .O(N__45520),
            .I(N__45517));
    InMux I__8065 (
            .O(N__45517),
            .I(N__45514));
    LocalMux I__8064 (
            .O(N__45514),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n280 ));
    InMux I__8063 (
            .O(N__45511),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17270 ));
    InMux I__8062 (
            .O(N__45508),
            .I(N__45505));
    LocalMux I__8061 (
            .O(N__45505),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n329 ));
    InMux I__8060 (
            .O(N__45502),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17271 ));
    CascadeMux I__8059 (
            .O(N__45499),
            .I(N__45496));
    InMux I__8058 (
            .O(N__45496),
            .I(N__45493));
    LocalMux I__8057 (
            .O(N__45493),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n378 ));
    InMux I__8056 (
            .O(N__45490),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17272 ));
    InMux I__8055 (
            .O(N__45487),
            .I(bfn_18_6_0_));
    InMux I__8054 (
            .O(N__45484),
            .I(N__45481));
    LocalMux I__8053 (
            .O(N__45481),
            .I(N__45478));
    Span4Mux_h I__8052 (
            .O(N__45478),
            .I(N__45474));
    InMux I__8051 (
            .O(N__45477),
            .I(N__45471));
    Span4Mux_h I__8050 (
            .O(N__45474),
            .I(N__45468));
    LocalMux I__8049 (
            .O(N__45471),
            .I(N__45465));
    Odrv4 I__8048 (
            .O(N__45468),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n769 ));
    Odrv4 I__8047 (
            .O(N__45465),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n769 ));
    InMux I__8046 (
            .O(N__45460),
            .I(bfn_17_26_0_));
    InMux I__8045 (
            .O(N__45457),
            .I(N__45453));
    InMux I__8044 (
            .O(N__45456),
            .I(N__45450));
    LocalMux I__8043 (
            .O(N__45453),
            .I(N__45447));
    LocalMux I__8042 (
            .O(N__45450),
            .I(N__45444));
    Span4Mux_v I__8041 (
            .O(N__45447),
            .I(N__45441));
    Span4Mux_v I__8040 (
            .O(N__45444),
            .I(N__45438));
    Odrv4 I__8039 (
            .O(N__45441),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n773 ));
    Odrv4 I__8038 (
            .O(N__45438),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n773 ));
    InMux I__8037 (
            .O(N__45433),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18377 ));
    InMux I__8036 (
            .O(N__45430),
            .I(N__45427));
    LocalMux I__8035 (
            .O(N__45427),
            .I(N__45423));
    InMux I__8034 (
            .O(N__45426),
            .I(N__45420));
    Span4Mux_h I__8033 (
            .O(N__45423),
            .I(N__45417));
    LocalMux I__8032 (
            .O(N__45420),
            .I(N__45414));
    Span4Mux_v I__8031 (
            .O(N__45417),
            .I(N__45409));
    Span4Mux_v I__8030 (
            .O(N__45414),
            .I(N__45409));
    Odrv4 I__8029 (
            .O(N__45409),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n777 ));
    InMux I__8028 (
            .O(N__45406),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18378 ));
    InMux I__8027 (
            .O(N__45403),
            .I(N__45400));
    LocalMux I__8026 (
            .O(N__45400),
            .I(N__45396));
    InMux I__8025 (
            .O(N__45399),
            .I(N__45393));
    Span4Mux_v I__8024 (
            .O(N__45396),
            .I(N__45390));
    LocalMux I__8023 (
            .O(N__45393),
            .I(N__45387));
    Odrv4 I__8022 (
            .O(N__45390),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n781 ));
    Odrv12 I__8021 (
            .O(N__45387),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n781 ));
    InMux I__8020 (
            .O(N__45382),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18379 ));
    CascadeMux I__8019 (
            .O(N__45379),
            .I(N__45376));
    InMux I__8018 (
            .O(N__45376),
            .I(N__45372));
    InMux I__8017 (
            .O(N__45375),
            .I(N__45369));
    LocalMux I__8016 (
            .O(N__45372),
            .I(N__45366));
    LocalMux I__8015 (
            .O(N__45369),
            .I(N__45363));
    Odrv12 I__8014 (
            .O(N__45366),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n785 ));
    Odrv4 I__8013 (
            .O(N__45363),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n785 ));
    InMux I__8012 (
            .O(N__45358),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18380 ));
    CascadeMux I__8011 (
            .O(N__45355),
            .I(N__45352));
    InMux I__8010 (
            .O(N__45352),
            .I(N__45349));
    LocalMux I__8009 (
            .O(N__45349),
            .I(N__45346));
    Odrv12 I__8008 (
            .O(N__45346),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n789 ));
    InMux I__8007 (
            .O(N__45343),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18381 ));
    InMux I__8006 (
            .O(N__45340),
            .I(N__45337));
    LocalMux I__8005 (
            .O(N__45337),
            .I(N__45334));
    Odrv12 I__8004 (
            .O(N__45334),
            .I(n793_adj_2424));
    InMux I__8003 (
            .O(N__45331),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18382 ));
    InMux I__8002 (
            .O(N__45328),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n795 ));
    CascadeMux I__8001 (
            .O(N__45325),
            .I(N__45322));
    InMux I__8000 (
            .O(N__45322),
            .I(N__45318));
    InMux I__7999 (
            .O(N__45321),
            .I(N__45315));
    LocalMux I__7998 (
            .O(N__45318),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n737 ));
    LocalMux I__7997 (
            .O(N__45315),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n737 ));
    InMux I__7996 (
            .O(N__45310),
            .I(N__45307));
    LocalMux I__7995 (
            .O(N__45307),
            .I(N__45304));
    Span4Mux_v I__7994 (
            .O(N__45304),
            .I(N__45300));
    InMux I__7993 (
            .O(N__45303),
            .I(N__45297));
    Odrv4 I__7992 (
            .O(N__45300),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n741 ));
    LocalMux I__7991 (
            .O(N__45297),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n741 ));
    InMux I__7990 (
            .O(N__45292),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18369 ));
    CascadeMux I__7989 (
            .O(N__45289),
            .I(N__45286));
    InMux I__7988 (
            .O(N__45286),
            .I(N__45283));
    LocalMux I__7987 (
            .O(N__45283),
            .I(N__45279));
    InMux I__7986 (
            .O(N__45282),
            .I(N__45276));
    Odrv4 I__7985 (
            .O(N__45279),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n745 ));
    LocalMux I__7984 (
            .O(N__45276),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n745 ));
    InMux I__7983 (
            .O(N__45271),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18370 ));
    InMux I__7982 (
            .O(N__45268),
            .I(N__45265));
    LocalMux I__7981 (
            .O(N__45265),
            .I(N__45262));
    Span4Mux_v I__7980 (
            .O(N__45262),
            .I(N__45259));
    Sp12to4 I__7979 (
            .O(N__45259),
            .I(N__45255));
    InMux I__7978 (
            .O(N__45258),
            .I(N__45252));
    Span12Mux_h I__7977 (
            .O(N__45255),
            .I(N__45247));
    LocalMux I__7976 (
            .O(N__45252),
            .I(N__45247));
    Odrv12 I__7975 (
            .O(N__45247),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n749 ));
    InMux I__7974 (
            .O(N__45244),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18371 ));
    InMux I__7973 (
            .O(N__45241),
            .I(N__45238));
    LocalMux I__7972 (
            .O(N__45238),
            .I(N__45234));
    InMux I__7971 (
            .O(N__45237),
            .I(N__45231));
    Span4Mux_v I__7970 (
            .O(N__45234),
            .I(N__45228));
    LocalMux I__7969 (
            .O(N__45231),
            .I(N__45225));
    Odrv4 I__7968 (
            .O(N__45228),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n753 ));
    Odrv4 I__7967 (
            .O(N__45225),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n753 ));
    InMux I__7966 (
            .O(N__45220),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18372 ));
    InMux I__7965 (
            .O(N__45217),
            .I(N__45214));
    LocalMux I__7964 (
            .O(N__45214),
            .I(N__45210));
    InMux I__7963 (
            .O(N__45213),
            .I(N__45207));
    Span4Mux_h I__7962 (
            .O(N__45210),
            .I(N__45204));
    LocalMux I__7961 (
            .O(N__45207),
            .I(N__45201));
    Odrv4 I__7960 (
            .O(N__45204),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n757 ));
    Odrv12 I__7959 (
            .O(N__45201),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n757 ));
    InMux I__7958 (
            .O(N__45196),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18373 ));
    InMux I__7957 (
            .O(N__45193),
            .I(N__45190));
    LocalMux I__7956 (
            .O(N__45190),
            .I(N__45186));
    InMux I__7955 (
            .O(N__45189),
            .I(N__45183));
    Span4Mux_v I__7954 (
            .O(N__45186),
            .I(N__45180));
    LocalMux I__7953 (
            .O(N__45183),
            .I(N__45177));
    Odrv4 I__7952 (
            .O(N__45180),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n761 ));
    Odrv4 I__7951 (
            .O(N__45177),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n761 ));
    InMux I__7950 (
            .O(N__45172),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18374 ));
    InMux I__7949 (
            .O(N__45169),
            .I(N__45166));
    LocalMux I__7948 (
            .O(N__45166),
            .I(N__45163));
    Span4Mux_h I__7947 (
            .O(N__45163),
            .I(N__45159));
    InMux I__7946 (
            .O(N__45162),
            .I(N__45156));
    Odrv4 I__7945 (
            .O(N__45159),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n765 ));
    LocalMux I__7944 (
            .O(N__45156),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n765 ));
    InMux I__7943 (
            .O(N__45151),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18375 ));
    InMux I__7942 (
            .O(N__45148),
            .I(N__45142));
    InMux I__7941 (
            .O(N__45147),
            .I(N__45142));
    LocalMux I__7940 (
            .O(N__45142),
            .I(N__45139));
    Span4Mux_v I__7939 (
            .O(N__45139),
            .I(N__45136));
    Odrv4 I__7938 (
            .O(N__45136),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20 ));
    InMux I__7937 (
            .O(N__45133),
            .I(N__45130));
    LocalMux I__7936 (
            .O(N__45130),
            .I(N__45116));
    InMux I__7935 (
            .O(N__45129),
            .I(N__45113));
    InMux I__7934 (
            .O(N__45128),
            .I(N__45108));
    InMux I__7933 (
            .O(N__45127),
            .I(N__45108));
    InMux I__7932 (
            .O(N__45126),
            .I(N__45101));
    InMux I__7931 (
            .O(N__45125),
            .I(N__45101));
    InMux I__7930 (
            .O(N__45124),
            .I(N__45101));
    InMux I__7929 (
            .O(N__45123),
            .I(N__45094));
    InMux I__7928 (
            .O(N__45122),
            .I(N__45094));
    InMux I__7927 (
            .O(N__45121),
            .I(N__45094));
    InMux I__7926 (
            .O(N__45120),
            .I(N__45089));
    InMux I__7925 (
            .O(N__45119),
            .I(N__45089));
    Odrv4 I__7924 (
            .O(N__45116),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7923 (
            .O(N__45113),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7922 (
            .O(N__45108),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7921 (
            .O(N__45101),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7920 (
            .O(N__45094),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7919 (
            .O(N__45089),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ));
    InMux I__7918 (
            .O(N__45076),
            .I(N__45073));
    LocalMux I__7917 (
            .O(N__45073),
            .I(N__45069));
    InMux I__7916 (
            .O(N__45072),
            .I(N__45066));
    Span4Mux_v I__7915 (
            .O(N__45069),
            .I(N__45063));
    LocalMux I__7914 (
            .O(N__45066),
            .I(N__45060));
    Odrv4 I__7913 (
            .O(N__45063),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18 ));
    Odrv4 I__7912 (
            .O(N__45060),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18 ));
    InMux I__7911 (
            .O(N__45055),
            .I(N__45052));
    LocalMux I__7910 (
            .O(N__45052),
            .I(N__45044));
    InMux I__7909 (
            .O(N__45051),
            .I(N__45041));
    InMux I__7908 (
            .O(N__45050),
            .I(N__45036));
    InMux I__7907 (
            .O(N__45049),
            .I(N__45036));
    InMux I__7906 (
            .O(N__45048),
            .I(N__45031));
    InMux I__7905 (
            .O(N__45047),
            .I(N__45031));
    Odrv4 I__7904 (
            .O(N__45044),
            .I(Error_sub_temp_30_adj_2385));
    LocalMux I__7903 (
            .O(N__45041),
            .I(Error_sub_temp_30_adj_2385));
    LocalMux I__7902 (
            .O(N__45036),
            .I(Error_sub_temp_30_adj_2385));
    LocalMux I__7901 (
            .O(N__45031),
            .I(Error_sub_temp_30_adj_2385));
    InMux I__7900 (
            .O(N__45022),
            .I(N__45019));
    LocalMux I__7899 (
            .O(N__45019),
            .I(N__45015));
    InMux I__7898 (
            .O(N__45018),
            .I(N__45012));
    Span4Mux_v I__7897 (
            .O(N__45015),
            .I(N__45007));
    LocalMux I__7896 (
            .O(N__45012),
            .I(N__45007));
    Odrv4 I__7895 (
            .O(N__45007),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16 ));
    InMux I__7894 (
            .O(N__45004),
            .I(N__45001));
    LocalMux I__7893 (
            .O(N__45001),
            .I(N__44998));
    Span4Mux_v I__7892 (
            .O(N__44998),
            .I(N__44994));
    InMux I__7891 (
            .O(N__44997),
            .I(N__44991));
    Odrv4 I__7890 (
            .O(N__44994),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23 ));
    LocalMux I__7889 (
            .O(N__44991),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23 ));
    CascadeMux I__7888 (
            .O(N__44986),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_ ));
    InMux I__7887 (
            .O(N__44983),
            .I(N__44980));
    LocalMux I__7886 (
            .O(N__44980),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743 ));
    CascadeMux I__7885 (
            .O(N__44977),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_ ));
    CascadeMux I__7884 (
            .O(N__44974),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_ ));
    InMux I__7883 (
            .O(N__44971),
            .I(N__44968));
    LocalMux I__7882 (
            .O(N__44968),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22 ));
    CascadeMux I__7881 (
            .O(N__44965),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_ ));
    InMux I__7880 (
            .O(N__44962),
            .I(N__44959));
    LocalMux I__7879 (
            .O(N__44959),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812 ));
    CascadeMux I__7878 (
            .O(N__44956),
            .I(N__44943));
    InMux I__7877 (
            .O(N__44955),
            .I(N__44937));
    InMux I__7876 (
            .O(N__44954),
            .I(N__44937));
    InMux I__7875 (
            .O(N__44953),
            .I(N__44934));
    InMux I__7874 (
            .O(N__44952),
            .I(N__44925));
    InMux I__7873 (
            .O(N__44951),
            .I(N__44925));
    InMux I__7872 (
            .O(N__44950),
            .I(N__44925));
    InMux I__7871 (
            .O(N__44949),
            .I(N__44925));
    InMux I__7870 (
            .O(N__44948),
            .I(N__44918));
    InMux I__7869 (
            .O(N__44947),
            .I(N__44918));
    InMux I__7868 (
            .O(N__44946),
            .I(N__44918));
    InMux I__7867 (
            .O(N__44943),
            .I(N__44913));
    InMux I__7866 (
            .O(N__44942),
            .I(N__44913));
    LocalMux I__7865 (
            .O(N__44937),
            .I(N__44908));
    LocalMux I__7864 (
            .O(N__44934),
            .I(N__44901));
    LocalMux I__7863 (
            .O(N__44925),
            .I(N__44901));
    LocalMux I__7862 (
            .O(N__44918),
            .I(N__44901));
    LocalMux I__7861 (
            .O(N__44913),
            .I(N__44898));
    InMux I__7860 (
            .O(N__44912),
            .I(N__44895));
    InMux I__7859 (
            .O(N__44911),
            .I(N__44890));
    Span4Mux_v I__7858 (
            .O(N__44908),
            .I(N__44885));
    Span4Mux_v I__7857 (
            .O(N__44901),
            .I(N__44885));
    Span4Mux_v I__7856 (
            .O(N__44898),
            .I(N__44880));
    LocalMux I__7855 (
            .O(N__44895),
            .I(N__44880));
    InMux I__7854 (
            .O(N__44894),
            .I(N__44877));
    CascadeMux I__7853 (
            .O(N__44893),
            .I(N__44874));
    LocalMux I__7852 (
            .O(N__44890),
            .I(N__44871));
    Span4Mux_h I__7851 (
            .O(N__44885),
            .I(N__44864));
    Span4Mux_h I__7850 (
            .O(N__44880),
            .I(N__44864));
    LocalMux I__7849 (
            .O(N__44877),
            .I(N__44864));
    InMux I__7848 (
            .O(N__44874),
            .I(N__44861));
    Span4Mux_v I__7847 (
            .O(N__44871),
            .I(N__44857));
    Span4Mux_v I__7846 (
            .O(N__44864),
            .I(N__44852));
    LocalMux I__7845 (
            .O(N__44861),
            .I(N__44852));
    CascadeMux I__7844 (
            .O(N__44860),
            .I(N__44849));
    Span4Mux_h I__7843 (
            .O(N__44857),
            .I(N__44846));
    Span4Mux_v I__7842 (
            .O(N__44852),
            .I(N__44843));
    InMux I__7841 (
            .O(N__44849),
            .I(N__44840));
    Odrv4 I__7840 (
            .O(N__44846),
            .I(Amp25_out1_14));
    Odrv4 I__7839 (
            .O(N__44843),
            .I(Amp25_out1_14));
    LocalMux I__7838 (
            .O(N__44840),
            .I(Amp25_out1_14));
    InMux I__7837 (
            .O(N__44833),
            .I(N__44829));
    CascadeMux I__7836 (
            .O(N__44832),
            .I(N__44824));
    LocalMux I__7835 (
            .O(N__44829),
            .I(N__44818));
    InMux I__7834 (
            .O(N__44828),
            .I(N__44815));
    InMux I__7833 (
            .O(N__44827),
            .I(N__44808));
    InMux I__7832 (
            .O(N__44824),
            .I(N__44808));
    InMux I__7831 (
            .O(N__44823),
            .I(N__44808));
    InMux I__7830 (
            .O(N__44822),
            .I(N__44802));
    InMux I__7829 (
            .O(N__44821),
            .I(N__44802));
    Span4Mux_v I__7828 (
            .O(N__44818),
            .I(N__44795));
    LocalMux I__7827 (
            .O(N__44815),
            .I(N__44795));
    LocalMux I__7826 (
            .O(N__44808),
            .I(N__44795));
    InMux I__7825 (
            .O(N__44807),
            .I(N__44792));
    LocalMux I__7824 (
            .O(N__44802),
            .I(n142_adj_2422));
    Odrv4 I__7823 (
            .O(N__44795),
            .I(n142_adj_2422));
    LocalMux I__7822 (
            .O(N__44792),
            .I(n142_adj_2422));
    InMux I__7821 (
            .O(N__44785),
            .I(N__44782));
    LocalMux I__7820 (
            .O(N__44782),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763 ));
    InMux I__7819 (
            .O(N__44779),
            .I(N__44776));
    LocalMux I__7818 (
            .O(N__44776),
            .I(N__44773));
    Odrv12 I__7817 (
            .O(N__44773),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727 ));
    CascadeMux I__7816 (
            .O(N__44770),
            .I(n141_adj_2421_cascade_));
    InMux I__7815 (
            .O(N__44767),
            .I(N__44759));
    InMux I__7814 (
            .O(N__44766),
            .I(N__44759));
    InMux I__7813 (
            .O(N__44765),
            .I(N__44754));
    InMux I__7812 (
            .O(N__44764),
            .I(N__44754));
    LocalMux I__7811 (
            .O(N__44759),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761 ));
    LocalMux I__7810 (
            .O(N__44754),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761 ));
    InMux I__7809 (
            .O(N__44749),
            .I(N__44745));
    InMux I__7808 (
            .O(N__44748),
            .I(N__44742));
    LocalMux I__7807 (
            .O(N__44745),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19 ));
    LocalMux I__7806 (
            .O(N__44742),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19 ));
    InMux I__7805 (
            .O(N__44737),
            .I(N__44734));
    LocalMux I__7804 (
            .O(N__44734),
            .I(N__44731));
    Odrv12 I__7803 (
            .O(N__44731),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n602 ));
    InMux I__7802 (
            .O(N__44728),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17777 ));
    CascadeMux I__7801 (
            .O(N__44725),
            .I(N__44722));
    InMux I__7800 (
            .O(N__44722),
            .I(N__44719));
    LocalMux I__7799 (
            .O(N__44719),
            .I(N__44716));
    Odrv4 I__7798 (
            .O(N__44716),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474 ));
    InMux I__7797 (
            .O(N__44713),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17778 ));
    CascadeMux I__7796 (
            .O(N__44710),
            .I(N__44707));
    InMux I__7795 (
            .O(N__44707),
            .I(N__44704));
    LocalMux I__7794 (
            .O(N__44704),
            .I(N__44701));
    Odrv4 I__7793 (
            .O(N__44701),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455 ));
    InMux I__7792 (
            .O(N__44698),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17779 ));
    InMux I__7791 (
            .O(N__44695),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n751 ));
    CascadeMux I__7790 (
            .O(N__44692),
            .I(n142_adj_2422_cascade_));
    CascadeMux I__7789 (
            .O(N__44689),
            .I(N__44684));
    InMux I__7788 (
            .O(N__44688),
            .I(N__44677));
    InMux I__7787 (
            .O(N__44687),
            .I(N__44677));
    InMux I__7786 (
            .O(N__44684),
            .I(N__44677));
    LocalMux I__7785 (
            .O(N__44677),
            .I(N__44674));
    Odrv4 I__7784 (
            .O(N__44674),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755 ));
    CascadeMux I__7783 (
            .O(N__44671),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_ ));
    InMux I__7782 (
            .O(N__44668),
            .I(N__44662));
    InMux I__7781 (
            .O(N__44667),
            .I(N__44662));
    LocalMux I__7780 (
            .O(N__44662),
            .I(N__44659));
    Odrv4 I__7779 (
            .O(N__44659),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756 ));
    InMux I__7778 (
            .O(N__44656),
            .I(N__44653));
    LocalMux I__7777 (
            .O(N__44653),
            .I(N__44650));
    Odrv4 I__7776 (
            .O(N__44650),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n161 ));
    InMux I__7775 (
            .O(N__44647),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17768 ));
    InMux I__7774 (
            .O(N__44644),
            .I(N__44641));
    LocalMux I__7773 (
            .O(N__44641),
            .I(N__44638));
    Odrv12 I__7772 (
            .O(N__44638),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n210 ));
    InMux I__7771 (
            .O(N__44635),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17769 ));
    InMux I__7770 (
            .O(N__44632),
            .I(N__44629));
    LocalMux I__7769 (
            .O(N__44629),
            .I(N__44626));
    Odrv4 I__7768 (
            .O(N__44626),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n259 ));
    InMux I__7767 (
            .O(N__44623),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17770 ));
    InMux I__7766 (
            .O(N__44620),
            .I(N__44617));
    LocalMux I__7765 (
            .O(N__44617),
            .I(N__44614));
    Odrv4 I__7764 (
            .O(N__44614),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368 ));
    InMux I__7763 (
            .O(N__44611),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17771 ));
    CascadeMux I__7762 (
            .O(N__44608),
            .I(N__44605));
    InMux I__7761 (
            .O(N__44605),
            .I(N__44602));
    LocalMux I__7760 (
            .O(N__44602),
            .I(N__44599));
    Odrv4 I__7759 (
            .O(N__44599),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366 ));
    InMux I__7758 (
            .O(N__44596),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17772 ));
    InMux I__7757 (
            .O(N__44593),
            .I(N__44590));
    LocalMux I__7756 (
            .O(N__44590),
            .I(N__44587));
    Odrv12 I__7755 (
            .O(N__44587),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363 ));
    InMux I__7754 (
            .O(N__44584),
            .I(bfn_17_19_0_));
    InMux I__7753 (
            .O(N__44581),
            .I(N__44578));
    LocalMux I__7752 (
            .O(N__44578),
            .I(N__44575));
    Odrv12 I__7751 (
            .O(N__44575),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350 ));
    InMux I__7750 (
            .O(N__44572),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17774 ));
    CascadeMux I__7749 (
            .O(N__44569),
            .I(N__44566));
    InMux I__7748 (
            .O(N__44566),
            .I(N__44563));
    LocalMux I__7747 (
            .O(N__44563),
            .I(N__44560));
    Odrv12 I__7746 (
            .O(N__44560),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n504 ));
    InMux I__7745 (
            .O(N__44557),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17775 ));
    InMux I__7744 (
            .O(N__44554),
            .I(N__44551));
    LocalMux I__7743 (
            .O(N__44551),
            .I(N__44548));
    Odrv4 I__7742 (
            .O(N__44548),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n553 ));
    InMux I__7741 (
            .O(N__44545),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17776 ));
    InMux I__7740 (
            .O(N__44542),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17790 ));
    InMux I__7739 (
            .O(N__44539),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17791 ));
    InMux I__7738 (
            .O(N__44536),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17792 ));
    InMux I__7737 (
            .O(N__44533),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17793 ));
    InMux I__7736 (
            .O(N__44530),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17794 ));
    InMux I__7735 (
            .O(N__44527),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n755 ));
    InMux I__7734 (
            .O(N__44524),
            .I(N__44521));
    LocalMux I__7733 (
            .O(N__44521),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384 ));
    InMux I__7732 (
            .O(N__44518),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17766 ));
    InMux I__7731 (
            .O(N__44515),
            .I(N__44512));
    LocalMux I__7730 (
            .O(N__44512),
            .I(N__44509));
    Odrv12 I__7729 (
            .O(N__44509),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n112 ));
    InMux I__7728 (
            .O(N__44506),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17767 ));
    InMux I__7727 (
            .O(N__44503),
            .I(N__44500));
    LocalMux I__7726 (
            .O(N__44500),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433 ));
    InMux I__7725 (
            .O(N__44497),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17781 ));
    InMux I__7724 (
            .O(N__44494),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17782 ));
    InMux I__7723 (
            .O(N__44491),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17783 ));
    InMux I__7722 (
            .O(N__44488),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17784 ));
    InMux I__7721 (
            .O(N__44485),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17785 ));
    InMux I__7720 (
            .O(N__44482),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17786 ));
    InMux I__7719 (
            .O(N__44479),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17787 ));
    InMux I__7718 (
            .O(N__44476),
            .I(bfn_17_16_0_));
    InMux I__7717 (
            .O(N__44473),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17789 ));
    CascadeMux I__7716 (
            .O(N__44470),
            .I(\foc.u_Park_Transform.n7_cascade_ ));
    InMux I__7715 (
            .O(N__44467),
            .I(N__44464));
    LocalMux I__7714 (
            .O(N__44464),
            .I(N__44460));
    InMux I__7713 (
            .O(N__44463),
            .I(N__44457));
    Span4Mux_v I__7712 (
            .O(N__44460),
            .I(N__44454));
    LocalMux I__7711 (
            .O(N__44457),
            .I(N__44451));
    Span4Mux_h I__7710 (
            .O(N__44454),
            .I(N__44448));
    Span4Mux_v I__7709 (
            .O(N__44451),
            .I(N__44445));
    Odrv4 I__7708 (
            .O(N__44448),
            .I(\foc.u_Park_Transform.n791 ));
    Odrv4 I__7707 (
            .O(N__44445),
            .I(\foc.u_Park_Transform.n791 ));
    CascadeMux I__7706 (
            .O(N__44440),
            .I(\foc.u_Park_Transform.n4_cascade_ ));
    InMux I__7705 (
            .O(N__44437),
            .I(N__44431));
    InMux I__7704 (
            .O(N__44436),
            .I(N__44428));
    InMux I__7703 (
            .O(N__44435),
            .I(N__44423));
    InMux I__7702 (
            .O(N__44434),
            .I(N__44423));
    LocalMux I__7701 (
            .O(N__44431),
            .I(N__44419));
    LocalMux I__7700 (
            .O(N__44428),
            .I(N__44414));
    LocalMux I__7699 (
            .O(N__44423),
            .I(N__44414));
    InMux I__7698 (
            .O(N__44422),
            .I(N__44411));
    Span4Mux_v I__7697 (
            .O(N__44419),
            .I(N__44406));
    Span12Mux_v I__7696 (
            .O(N__44414),
            .I(N__44401));
    LocalMux I__7695 (
            .O(N__44411),
            .I(N__44401));
    InMux I__7694 (
            .O(N__44410),
            .I(N__44396));
    InMux I__7693 (
            .O(N__44409),
            .I(N__44396));
    Sp12to4 I__7692 (
            .O(N__44406),
            .I(N__44387));
    Span12Mux_h I__7691 (
            .O(N__44401),
            .I(N__44387));
    LocalMux I__7690 (
            .O(N__44396),
            .I(N__44384));
    InMux I__7689 (
            .O(N__44395),
            .I(N__44375));
    InMux I__7688 (
            .O(N__44394),
            .I(N__44375));
    InMux I__7687 (
            .O(N__44393),
            .I(N__44375));
    InMux I__7686 (
            .O(N__44392),
            .I(N__44375));
    Odrv12 I__7685 (
            .O(N__44387),
            .I(Look_Up_Table_out1_1_13));
    Odrv4 I__7684 (
            .O(N__44384),
            .I(Look_Up_Table_out1_1_13));
    LocalMux I__7683 (
            .O(N__44375),
            .I(Look_Up_Table_out1_1_13));
    InMux I__7682 (
            .O(N__44368),
            .I(N__44365));
    LocalMux I__7681 (
            .O(N__44365),
            .I(N__44361));
    InMux I__7680 (
            .O(N__44364),
            .I(N__44358));
    Odrv4 I__7679 (
            .O(N__44361),
            .I(\foc.u_Park_Transform.n14 ));
    LocalMux I__7678 (
            .O(N__44358),
            .I(\foc.u_Park_Transform.n14 ));
    CascadeMux I__7677 (
            .O(N__44353),
            .I(n628_cascade_));
    CascadeMux I__7676 (
            .O(N__44350),
            .I(N__44346));
    InMux I__7675 (
            .O(N__44349),
            .I(N__44341));
    InMux I__7674 (
            .O(N__44346),
            .I(N__44341));
    LocalMux I__7673 (
            .O(N__44341),
            .I(N__44336));
    InMux I__7672 (
            .O(N__44340),
            .I(N__44333));
    InMux I__7671 (
            .O(N__44339),
            .I(N__44330));
    Odrv4 I__7670 (
            .O(N__44336),
            .I(\foc.u_Park_Transform.n12 ));
    LocalMux I__7669 (
            .O(N__44333),
            .I(\foc.u_Park_Transform.n12 ));
    LocalMux I__7668 (
            .O(N__44330),
            .I(\foc.u_Park_Transform.n12 ));
    InMux I__7667 (
            .O(N__44323),
            .I(N__44320));
    LocalMux I__7666 (
            .O(N__44320),
            .I(N__44310));
    InMux I__7665 (
            .O(N__44319),
            .I(N__44305));
    InMux I__7664 (
            .O(N__44318),
            .I(N__44305));
    InMux I__7663 (
            .O(N__44317),
            .I(N__44298));
    InMux I__7662 (
            .O(N__44316),
            .I(N__44298));
    InMux I__7661 (
            .O(N__44315),
            .I(N__44298));
    InMux I__7660 (
            .O(N__44314),
            .I(N__44293));
    InMux I__7659 (
            .O(N__44313),
            .I(N__44293));
    Span4Mux_h I__7658 (
            .O(N__44310),
            .I(N__44288));
    LocalMux I__7657 (
            .O(N__44305),
            .I(N__44285));
    LocalMux I__7656 (
            .O(N__44298),
            .I(N__44282));
    LocalMux I__7655 (
            .O(N__44293),
            .I(N__44279));
    InMux I__7654 (
            .O(N__44292),
            .I(N__44274));
    InMux I__7653 (
            .O(N__44291),
            .I(N__44274));
    Span4Mux_v I__7652 (
            .O(N__44288),
            .I(N__44271));
    Span4Mux_h I__7651 (
            .O(N__44285),
            .I(N__44268));
    Span4Mux_h I__7650 (
            .O(N__44282),
            .I(N__44261));
    Span4Mux_h I__7649 (
            .O(N__44279),
            .I(N__44261));
    LocalMux I__7648 (
            .O(N__44274),
            .I(N__44261));
    Odrv4 I__7647 (
            .O(N__44271),
            .I(n142));
    Odrv4 I__7646 (
            .O(N__44268),
            .I(n142));
    Odrv4 I__7645 (
            .O(N__44261),
            .I(n142));
    InMux I__7644 (
            .O(N__44254),
            .I(N__44250));
    InMux I__7643 (
            .O(N__44253),
            .I(N__44247));
    LocalMux I__7642 (
            .O(N__44250),
            .I(N__44242));
    LocalMux I__7641 (
            .O(N__44247),
            .I(N__44242));
    Span4Mux_v I__7640 (
            .O(N__44242),
            .I(N__44236));
    InMux I__7639 (
            .O(N__44241),
            .I(N__44233));
    InMux I__7638 (
            .O(N__44240),
            .I(N__44230));
    InMux I__7637 (
            .O(N__44239),
            .I(N__44227));
    Sp12to4 I__7636 (
            .O(N__44236),
            .I(N__44217));
    LocalMux I__7635 (
            .O(N__44233),
            .I(N__44217));
    LocalMux I__7634 (
            .O(N__44230),
            .I(N__44217));
    LocalMux I__7633 (
            .O(N__44227),
            .I(N__44214));
    InMux I__7632 (
            .O(N__44226),
            .I(N__44209));
    InMux I__7631 (
            .O(N__44225),
            .I(N__44209));
    InMux I__7630 (
            .O(N__44224),
            .I(N__44206));
    Odrv12 I__7629 (
            .O(N__44217),
            .I(n628));
    Odrv12 I__7628 (
            .O(N__44214),
            .I(n628));
    LocalMux I__7627 (
            .O(N__44209),
            .I(n628));
    LocalMux I__7626 (
            .O(N__44206),
            .I(n628));
    CascadeMux I__7625 (
            .O(N__44197),
            .I(\foc.u_Park_Transform.n18_cascade_ ));
    InMux I__7624 (
            .O(N__44194),
            .I(N__44191));
    LocalMux I__7623 (
            .O(N__44191),
            .I(\foc.u_Park_Transform.n19845 ));
    InMux I__7622 (
            .O(N__44188),
            .I(N__44183));
    InMux I__7621 (
            .O(N__44187),
            .I(N__44178));
    InMux I__7620 (
            .O(N__44186),
            .I(N__44178));
    LocalMux I__7619 (
            .O(N__44183),
            .I(N__44175));
    LocalMux I__7618 (
            .O(N__44178),
            .I(N__44172));
    Odrv12 I__7617 (
            .O(N__44175),
            .I(\foc.u_Park_Transform.n26 ));
    Odrv12 I__7616 (
            .O(N__44172),
            .I(\foc.u_Park_Transform.n26 ));
    InMux I__7615 (
            .O(N__44167),
            .I(N__44161));
    InMux I__7614 (
            .O(N__44166),
            .I(N__44161));
    LocalMux I__7613 (
            .O(N__44161),
            .I(N__44158));
    Span4Mux_v I__7612 (
            .O(N__44158),
            .I(N__44155));
    Odrv4 I__7611 (
            .O(N__44155),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28 ));
    InMux I__7610 (
            .O(N__44152),
            .I(N__44146));
    InMux I__7609 (
            .O(N__44151),
            .I(N__44146));
    LocalMux I__7608 (
            .O(N__44146),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n4 ));
    InMux I__7607 (
            .O(N__44143),
            .I(N__44133));
    InMux I__7606 (
            .O(N__44142),
            .I(N__44133));
    InMux I__7605 (
            .O(N__44141),
            .I(N__44130));
    InMux I__7604 (
            .O(N__44140),
            .I(N__44123));
    InMux I__7603 (
            .O(N__44139),
            .I(N__44123));
    InMux I__7602 (
            .O(N__44138),
            .I(N__44123));
    LocalMux I__7601 (
            .O(N__44133),
            .I(N__44116));
    LocalMux I__7600 (
            .O(N__44130),
            .I(N__44116));
    LocalMux I__7599 (
            .O(N__44123),
            .I(N__44116));
    Span4Mux_v I__7598 (
            .O(N__44116),
            .I(N__44111));
    InMux I__7597 (
            .O(N__44115),
            .I(N__44108));
    InMux I__7596 (
            .O(N__44114),
            .I(N__44105));
    Odrv4 I__7595 (
            .O(N__44111),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7594 (
            .O(N__44108),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29 ));
    LocalMux I__7593 (
            .O(N__44105),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29 ));
    CascadeMux I__7592 (
            .O(N__44098),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_ ));
    CascadeMux I__7591 (
            .O(N__44095),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_ ));
    CascadeMux I__7590 (
            .O(N__44092),
            .I(N__44088));
    CascadeMux I__7589 (
            .O(N__44091),
            .I(N__44083));
    InMux I__7588 (
            .O(N__44088),
            .I(N__44078));
    InMux I__7587 (
            .O(N__44087),
            .I(N__44078));
    InMux I__7586 (
            .O(N__44086),
            .I(N__44073));
    InMux I__7585 (
            .O(N__44083),
            .I(N__44073));
    LocalMux I__7584 (
            .O(N__44078),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n12 ));
    LocalMux I__7583 (
            .O(N__44073),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n12 ));
    InMux I__7582 (
            .O(N__44068),
            .I(N__44065));
    LocalMux I__7581 (
            .O(N__44065),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19273 ));
    InMux I__7580 (
            .O(N__44062),
            .I(N__44047));
    InMux I__7579 (
            .O(N__44061),
            .I(N__44047));
    InMux I__7578 (
            .O(N__44060),
            .I(N__44047));
    InMux I__7577 (
            .O(N__44059),
            .I(N__44047));
    InMux I__7576 (
            .O(N__44058),
            .I(N__44042));
    InMux I__7575 (
            .O(N__44057),
            .I(N__44042));
    InMux I__7574 (
            .O(N__44056),
            .I(N__44039));
    LocalMux I__7573 (
            .O(N__44047),
            .I(n142_adj_2419));
    LocalMux I__7572 (
            .O(N__44042),
            .I(n142_adj_2419));
    LocalMux I__7571 (
            .O(N__44039),
            .I(n142_adj_2419));
    CascadeMux I__7570 (
            .O(N__44032),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_ ));
    InMux I__7569 (
            .O(N__44029),
            .I(N__44026));
    LocalMux I__7568 (
            .O(N__44026),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19269 ));
    CascadeMux I__7567 (
            .O(N__44023),
            .I(N__44020));
    InMux I__7566 (
            .O(N__44020),
            .I(N__44017));
    LocalMux I__7565 (
            .O(N__44017),
            .I(N__44014));
    Odrv4 I__7564 (
            .O(N__44014),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n283 ));
    InMux I__7563 (
            .O(N__44011),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18170 ));
    CascadeMux I__7562 (
            .O(N__44008),
            .I(N__44004));
    CascadeMux I__7561 (
            .O(N__44007),
            .I(N__44000));
    InMux I__7560 (
            .O(N__44004),
            .I(N__43995));
    InMux I__7559 (
            .O(N__44003),
            .I(N__43995));
    InMux I__7558 (
            .O(N__44000),
            .I(N__43992));
    LocalMux I__7557 (
            .O(N__43995),
            .I(N__43987));
    LocalMux I__7556 (
            .O(N__43992),
            .I(N__43987));
    Odrv4 I__7555 (
            .O(N__43987),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n332 ));
    InMux I__7554 (
            .O(N__43984),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18171 ));
    InMux I__7553 (
            .O(N__43981),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18172 ));
    InMux I__7552 (
            .O(N__43978),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n787 ));
    InMux I__7551 (
            .O(N__43975),
            .I(N__43972));
    LocalMux I__7550 (
            .O(N__43972),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n188 ));
    CascadeMux I__7549 (
            .O(N__43969),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_ ));
    InMux I__7548 (
            .O(N__43966),
            .I(N__43963));
    LocalMux I__7547 (
            .O(N__43963),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n139 ));
    CascadeMux I__7546 (
            .O(N__43960),
            .I(N__43956));
    CascadeMux I__7545 (
            .O(N__43959),
            .I(N__43953));
    InMux I__7544 (
            .O(N__43956),
            .I(N__43949));
    InMux I__7543 (
            .O(N__43953),
            .I(N__43944));
    InMux I__7542 (
            .O(N__43952),
            .I(N__43944));
    LocalMux I__7541 (
            .O(N__43949),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n237 ));
    LocalMux I__7540 (
            .O(N__43944),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n237 ));
    InMux I__7539 (
            .O(N__43939),
            .I(N__43933));
    InMux I__7538 (
            .O(N__43938),
            .I(N__43933));
    LocalMux I__7537 (
            .O(N__43933),
            .I(N__43930));
    Span4Mux_v I__7536 (
            .O(N__43930),
            .I(N__43927));
    Odrv4 I__7535 (
            .O(N__43927),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27 ));
    InMux I__7534 (
            .O(N__43924),
            .I(N__43918));
    InMux I__7533 (
            .O(N__43923),
            .I(N__43918));
    LocalMux I__7532 (
            .O(N__43918),
            .I(N__43915));
    Odrv12 I__7531 (
            .O(N__43915),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21 ));
    CascadeMux I__7530 (
            .O(N__43912),
            .I(N__43909));
    InMux I__7529 (
            .O(N__43909),
            .I(N__43906));
    LocalMux I__7528 (
            .O(N__43906),
            .I(N__43903));
    Sp12to4 I__7527 (
            .O(N__43903),
            .I(N__43900));
    Odrv12 I__7526 (
            .O(N__43900),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400 ));
    InMux I__7525 (
            .O(N__43897),
            .I(N__43894));
    LocalMux I__7524 (
            .O(N__43894),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n90 ));
    InMux I__7523 (
            .O(N__43891),
            .I(N__43888));
    LocalMux I__7522 (
            .O(N__43888),
            .I(N__43885));
    Odrv4 I__7521 (
            .O(N__43885),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399 ));
    InMux I__7520 (
            .O(N__43882),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18167 ));
    CascadeMux I__7519 (
            .O(N__43879),
            .I(N__43876));
    InMux I__7518 (
            .O(N__43876),
            .I(N__43873));
    LocalMux I__7517 (
            .O(N__43873),
            .I(N__43870));
    Odrv4 I__7516 (
            .O(N__43870),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398 ));
    InMux I__7515 (
            .O(N__43867),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18168 ));
    InMux I__7514 (
            .O(N__43864),
            .I(N__43861));
    LocalMux I__7513 (
            .O(N__43861),
            .I(N__43858));
    Odrv4 I__7512 (
            .O(N__43858),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397 ));
    InMux I__7511 (
            .O(N__43855),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18169 ));
    InMux I__7510 (
            .O(N__43852),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18138 ));
    InMux I__7509 (
            .O(N__43849),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18139 ));
    InMux I__7508 (
            .O(N__43846),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18140 ));
    InMux I__7507 (
            .O(N__43843),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18141 ));
    InMux I__7506 (
            .O(N__43840),
            .I(bfn_17_6_0_));
    InMux I__7505 (
            .O(N__43837),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349 ));
    InMux I__7504 (
            .O(N__43834),
            .I(N__43828));
    InMux I__7503 (
            .O(N__43833),
            .I(N__43828));
    LocalMux I__7502 (
            .O(N__43828),
            .I(N__43825));
    Span4Mux_v I__7501 (
            .O(N__43825),
            .I(N__43822));
    Odrv4 I__7500 (
            .O(N__43822),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26 ));
    InMux I__7499 (
            .O(N__43819),
            .I(N__43816));
    LocalMux I__7498 (
            .O(N__43816),
            .I(N__43813));
    Odrv12 I__7497 (
            .O(N__43813),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703 ));
    CascadeMux I__7496 (
            .O(N__43810),
            .I(N__43807));
    InMux I__7495 (
            .O(N__43807),
            .I(N__43804));
    LocalMux I__7494 (
            .O(N__43804),
            .I(N__43801));
    Odrv12 I__7493 (
            .O(N__43801),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n642 ));
    InMux I__7492 (
            .O(N__43798),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18013 ));
    InMux I__7491 (
            .O(N__43795),
            .I(N__43792));
    LocalMux I__7490 (
            .O(N__43792),
            .I(N__43789));
    Odrv4 I__7489 (
            .O(N__43789),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702 ));
    InMux I__7488 (
            .O(N__43786),
            .I(N__43783));
    LocalMux I__7487 (
            .O(N__43783),
            .I(N__43780));
    Span4Mux_v I__7486 (
            .O(N__43780),
            .I(N__43777));
    Odrv4 I__7485 (
            .O(N__43777),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717 ));
    InMux I__7484 (
            .O(N__43774),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18014 ));
    CascadeMux I__7483 (
            .O(N__43771),
            .I(N__43768));
    InMux I__7482 (
            .O(N__43768),
            .I(N__43765));
    LocalMux I__7481 (
            .O(N__43765),
            .I(N__43762));
    Odrv4 I__7480 (
            .O(N__43762),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701 ));
    InMux I__7479 (
            .O(N__43759),
            .I(N__43756));
    LocalMux I__7478 (
            .O(N__43756),
            .I(N__43753));
    Span12Mux_h I__7477 (
            .O(N__43753),
            .I(N__43750));
    Odrv12 I__7476 (
            .O(N__43750),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715 ));
    InMux I__7475 (
            .O(N__43747),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18015 ));
    InMux I__7474 (
            .O(N__43744),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716 ));
    CascadeMux I__7473 (
            .O(N__43741),
            .I(N__43738));
    InMux I__7472 (
            .O(N__43738),
            .I(N__43735));
    LocalMux I__7471 (
            .O(N__43735),
            .I(N__43732));
    Span12Mux_v I__7470 (
            .O(N__43732),
            .I(N__43729));
    Odrv12 I__7469 (
            .O(N__43729),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO ));
    InMux I__7468 (
            .O(N__43726),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18135 ));
    InMux I__7467 (
            .O(N__43723),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18136 ));
    InMux I__7466 (
            .O(N__43720),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18137 ));
    InMux I__7465 (
            .O(N__43717),
            .I(N__43714));
    LocalMux I__7464 (
            .O(N__43714),
            .I(N__43711));
    Odrv4 I__7463 (
            .O(N__43711),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711 ));
    InMux I__7462 (
            .O(N__43708),
            .I(N__43705));
    LocalMux I__7461 (
            .O(N__43705),
            .I(N__43702));
    Odrv12 I__7460 (
            .O(N__43702),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n250 ));
    InMux I__7459 (
            .O(N__43699),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18005 ));
    InMux I__7458 (
            .O(N__43696),
            .I(N__43693));
    LocalMux I__7457 (
            .O(N__43693),
            .I(N__43690));
    Odrv4 I__7456 (
            .O(N__43690),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710 ));
    CascadeMux I__7455 (
            .O(N__43687),
            .I(N__43684));
    InMux I__7454 (
            .O(N__43684),
            .I(N__43681));
    LocalMux I__7453 (
            .O(N__43681),
            .I(N__43678));
    Odrv12 I__7452 (
            .O(N__43678),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n299 ));
    InMux I__7451 (
            .O(N__43675),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18006 ));
    InMux I__7450 (
            .O(N__43672),
            .I(N__43669));
    LocalMux I__7449 (
            .O(N__43669),
            .I(N__43666));
    Odrv4 I__7448 (
            .O(N__43666),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709 ));
    InMux I__7447 (
            .O(N__43663),
            .I(N__43660));
    LocalMux I__7446 (
            .O(N__43660),
            .I(N__43657));
    Odrv12 I__7445 (
            .O(N__43657),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n348 ));
    InMux I__7444 (
            .O(N__43654),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18007 ));
    InMux I__7443 (
            .O(N__43651),
            .I(N__43648));
    LocalMux I__7442 (
            .O(N__43648),
            .I(N__43645));
    Odrv4 I__7441 (
            .O(N__43645),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708 ));
    InMux I__7440 (
            .O(N__43642),
            .I(N__43639));
    LocalMux I__7439 (
            .O(N__43639),
            .I(N__43636));
    Odrv12 I__7438 (
            .O(N__43636),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n397 ));
    InMux I__7437 (
            .O(N__43633),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18008 ));
    InMux I__7436 (
            .O(N__43630),
            .I(N__43627));
    LocalMux I__7435 (
            .O(N__43627),
            .I(N__43624));
    Odrv4 I__7434 (
            .O(N__43624),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707 ));
    InMux I__7433 (
            .O(N__43621),
            .I(N__43618));
    LocalMux I__7432 (
            .O(N__43618),
            .I(N__43615));
    Odrv12 I__7431 (
            .O(N__43615),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n446 ));
    InMux I__7430 (
            .O(N__43612),
            .I(bfn_16_28_0_));
    InMux I__7429 (
            .O(N__43609),
            .I(N__43606));
    LocalMux I__7428 (
            .O(N__43606),
            .I(N__43603));
    Odrv4 I__7427 (
            .O(N__43603),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706 ));
    InMux I__7426 (
            .O(N__43600),
            .I(N__43597));
    LocalMux I__7425 (
            .O(N__43597),
            .I(N__43594));
    Odrv12 I__7424 (
            .O(N__43594),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n495 ));
    InMux I__7423 (
            .O(N__43591),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18010 ));
    InMux I__7422 (
            .O(N__43588),
            .I(N__43585));
    LocalMux I__7421 (
            .O(N__43585),
            .I(N__43582));
    Odrv4 I__7420 (
            .O(N__43582),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705 ));
    InMux I__7419 (
            .O(N__43579),
            .I(N__43576));
    LocalMux I__7418 (
            .O(N__43576),
            .I(N__43573));
    Odrv12 I__7417 (
            .O(N__43573),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n544 ));
    InMux I__7416 (
            .O(N__43570),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18011 ));
    InMux I__7415 (
            .O(N__43567),
            .I(N__43564));
    LocalMux I__7414 (
            .O(N__43564),
            .I(N__43561));
    Odrv12 I__7413 (
            .O(N__43561),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704 ));
    InMux I__7412 (
            .O(N__43558),
            .I(N__43555));
    LocalMux I__7411 (
            .O(N__43555),
            .I(N__43552));
    Odrv12 I__7410 (
            .O(N__43552),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n593 ));
    InMux I__7409 (
            .O(N__43549),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18012 ));
    InMux I__7408 (
            .O(N__43546),
            .I(N__43543));
    LocalMux I__7407 (
            .O(N__43543),
            .I(N__43540));
    Odrv12 I__7406 (
            .O(N__43540),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687 ));
    InMux I__7405 (
            .O(N__43537),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18028 ));
    CascadeMux I__7404 (
            .O(N__43534),
            .I(N__43531));
    InMux I__7403 (
            .O(N__43531),
            .I(N__43528));
    LocalMux I__7402 (
            .O(N__43528),
            .I(N__43525));
    Odrv12 I__7401 (
            .O(N__43525),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686 ));
    InMux I__7400 (
            .O(N__43522),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18029 ));
    InMux I__7399 (
            .O(N__43519),
            .I(N__43516));
    LocalMux I__7398 (
            .O(N__43516),
            .I(N__43513));
    Odrv12 I__7397 (
            .O(N__43513),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685 ));
    InMux I__7396 (
            .O(N__43510),
            .I(N__43507));
    LocalMux I__7395 (
            .O(N__43507),
            .I(N__43504));
    Span4Mux_h I__7394 (
            .O(N__43504),
            .I(N__43501));
    Span4Mux_v I__7393 (
            .O(N__43501),
            .I(N__43498));
    Odrv4 I__7392 (
            .O(N__43498),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699 ));
    InMux I__7391 (
            .O(N__43495),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18030 ));
    InMux I__7390 (
            .O(N__43492),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700 ));
    CascadeMux I__7389 (
            .O(N__43489),
            .I(N__43486));
    InMux I__7388 (
            .O(N__43486),
            .I(N__43483));
    LocalMux I__7387 (
            .O(N__43483),
            .I(N__43480));
    Span4Mux_h I__7386 (
            .O(N__43480),
            .I(N__43477));
    Span4Mux_v I__7385 (
            .O(N__43477),
            .I(N__43474));
    Odrv4 I__7384 (
            .O(N__43474),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO ));
    CascadeMux I__7383 (
            .O(N__43471),
            .I(N__43468));
    InMux I__7382 (
            .O(N__43468),
            .I(N__43465));
    LocalMux I__7381 (
            .O(N__43465),
            .I(N__43462));
    Span4Mux_v I__7380 (
            .O(N__43462),
            .I(N__43459));
    Odrv4 I__7379 (
            .O(N__43459),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n54 ));
    CascadeMux I__7378 (
            .O(N__43456),
            .I(N__43453));
    InMux I__7377 (
            .O(N__43453),
            .I(N__43450));
    LocalMux I__7376 (
            .O(N__43450),
            .I(N__43447));
    Odrv4 I__7375 (
            .O(N__43447),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714 ));
    InMux I__7374 (
            .O(N__43444),
            .I(N__43441));
    LocalMux I__7373 (
            .O(N__43441),
            .I(N__43438));
    Odrv12 I__7372 (
            .O(N__43438),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n103 ));
    InMux I__7371 (
            .O(N__43435),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18002 ));
    InMux I__7370 (
            .O(N__43432),
            .I(N__43429));
    LocalMux I__7369 (
            .O(N__43429),
            .I(N__43426));
    Odrv4 I__7368 (
            .O(N__43426),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713 ));
    CascadeMux I__7367 (
            .O(N__43423),
            .I(N__43420));
    InMux I__7366 (
            .O(N__43420),
            .I(N__43417));
    LocalMux I__7365 (
            .O(N__43417),
            .I(N__43414));
    Odrv12 I__7364 (
            .O(N__43414),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n152 ));
    InMux I__7363 (
            .O(N__43411),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18003 ));
    InMux I__7362 (
            .O(N__43408),
            .I(N__43405));
    LocalMux I__7361 (
            .O(N__43405),
            .I(N__43402));
    Odrv12 I__7360 (
            .O(N__43402),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712 ));
    InMux I__7359 (
            .O(N__43399),
            .I(N__43396));
    LocalMux I__7358 (
            .O(N__43396),
            .I(N__43393));
    Odrv12 I__7357 (
            .O(N__43393),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n201 ));
    InMux I__7356 (
            .O(N__43390),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18004 ));
    CascadeMux I__7355 (
            .O(N__43387),
            .I(N__43384));
    InMux I__7354 (
            .O(N__43384),
            .I(N__43381));
    LocalMux I__7353 (
            .O(N__43381),
            .I(N__43378));
    Odrv12 I__7352 (
            .O(N__43378),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696 ));
    InMux I__7351 (
            .O(N__43375),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18019 ));
    InMux I__7350 (
            .O(N__43372),
            .I(N__43369));
    LocalMux I__7349 (
            .O(N__43369),
            .I(N__43366));
    Odrv4 I__7348 (
            .O(N__43366),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695 ));
    InMux I__7347 (
            .O(N__43363),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18020 ));
    CascadeMux I__7346 (
            .O(N__43360),
            .I(N__43357));
    InMux I__7345 (
            .O(N__43357),
            .I(N__43354));
    LocalMux I__7344 (
            .O(N__43354),
            .I(N__43351));
    Odrv4 I__7343 (
            .O(N__43351),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694 ));
    InMux I__7342 (
            .O(N__43348),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18021 ));
    InMux I__7341 (
            .O(N__43345),
            .I(N__43342));
    LocalMux I__7340 (
            .O(N__43342),
            .I(N__43339));
    Odrv12 I__7339 (
            .O(N__43339),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693 ));
    InMux I__7338 (
            .O(N__43336),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18022 ));
    CascadeMux I__7337 (
            .O(N__43333),
            .I(N__43330));
    InMux I__7336 (
            .O(N__43330),
            .I(N__43327));
    LocalMux I__7335 (
            .O(N__43327),
            .I(N__43324));
    Odrv4 I__7334 (
            .O(N__43324),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692 ));
    InMux I__7333 (
            .O(N__43321),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18023 ));
    InMux I__7332 (
            .O(N__43318),
            .I(N__43315));
    LocalMux I__7331 (
            .O(N__43315),
            .I(N__43312));
    Span4Mux_h I__7330 (
            .O(N__43312),
            .I(N__43309));
    Odrv4 I__7329 (
            .O(N__43309),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691 ));
    InMux I__7328 (
            .O(N__43306),
            .I(bfn_16_26_0_));
    CascadeMux I__7327 (
            .O(N__43303),
            .I(N__43300));
    InMux I__7326 (
            .O(N__43300),
            .I(N__43297));
    LocalMux I__7325 (
            .O(N__43297),
            .I(N__43294));
    Odrv4 I__7324 (
            .O(N__43294),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690 ));
    InMux I__7323 (
            .O(N__43291),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18025 ));
    InMux I__7322 (
            .O(N__43288),
            .I(N__43285));
    LocalMux I__7321 (
            .O(N__43285),
            .I(N__43282));
    Odrv4 I__7320 (
            .O(N__43282),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689 ));
    InMux I__7319 (
            .O(N__43279),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18026 ));
    CascadeMux I__7318 (
            .O(N__43276),
            .I(N__43273));
    InMux I__7317 (
            .O(N__43273),
            .I(N__43270));
    LocalMux I__7316 (
            .O(N__43270),
            .I(N__43267));
    Odrv12 I__7315 (
            .O(N__43267),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688 ));
    InMux I__7314 (
            .O(N__43264),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18027 ));
    InMux I__7313 (
            .O(N__43261),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17996 ));
    InMux I__7312 (
            .O(N__43258),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17997 ));
    InMux I__7311 (
            .O(N__43255),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17998 ));
    InMux I__7310 (
            .O(N__43252),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17999 ));
    CascadeMux I__7309 (
            .O(N__43249),
            .I(N__43246));
    InMux I__7308 (
            .O(N__43246),
            .I(N__43242));
    InMux I__7307 (
            .O(N__43245),
            .I(N__43239));
    LocalMux I__7306 (
            .O(N__43242),
            .I(N__43234));
    LocalMux I__7305 (
            .O(N__43239),
            .I(N__43234));
    Span4Mux_v I__7304 (
            .O(N__43234),
            .I(N__43231));
    Odrv4 I__7303 (
            .O(N__43231),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718 ));
    InMux I__7302 (
            .O(N__43228),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18000 ));
    InMux I__7301 (
            .O(N__43225),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n739 ));
    CascadeMux I__7300 (
            .O(N__43222),
            .I(N__43219));
    InMux I__7299 (
            .O(N__43219),
            .I(N__43216));
    LocalMux I__7298 (
            .O(N__43216),
            .I(N__43213));
    Span4Mux_h I__7297 (
            .O(N__43213),
            .I(N__43210));
    Odrv4 I__7296 (
            .O(N__43210),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO ));
    CascadeMux I__7295 (
            .O(N__43207),
            .I(N__43204));
    InMux I__7294 (
            .O(N__43204),
            .I(N__43201));
    LocalMux I__7293 (
            .O(N__43201),
            .I(N__43198));
    Odrv12 I__7292 (
            .O(N__43198),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698 ));
    InMux I__7291 (
            .O(N__43195),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18017 ));
    InMux I__7290 (
            .O(N__43192),
            .I(N__43189));
    LocalMux I__7289 (
            .O(N__43189),
            .I(N__43186));
    Odrv4 I__7288 (
            .O(N__43186),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697 ));
    InMux I__7287 (
            .O(N__43183),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18018 ));
    InMux I__7286 (
            .O(N__43180),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17987 ));
    InMux I__7285 (
            .O(N__43177),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17988 ));
    InMux I__7284 (
            .O(N__43174),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17989 ));
    InMux I__7283 (
            .O(N__43171),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17990 ));
    InMux I__7282 (
            .O(N__43168),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17991 ));
    InMux I__7281 (
            .O(N__43165),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17992 ));
    InMux I__7280 (
            .O(N__43162),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17993 ));
    InMux I__7279 (
            .O(N__43159),
            .I(bfn_16_24_0_));
    InMux I__7278 (
            .O(N__43156),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17995 ));
    InMux I__7277 (
            .O(N__43153),
            .I(N__43147));
    InMux I__7276 (
            .O(N__43152),
            .I(N__43147));
    LocalMux I__7275 (
            .O(N__43147),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27 ));
    InMux I__7274 (
            .O(N__43144),
            .I(N__43138));
    InMux I__7273 (
            .O(N__43143),
            .I(N__43138));
    LocalMux I__7272 (
            .O(N__43138),
            .I(N__43135));
    Odrv4 I__7271 (
            .O(N__43135),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25 ));
    InMux I__7270 (
            .O(N__43132),
            .I(N__43126));
    InMux I__7269 (
            .O(N__43131),
            .I(N__43126));
    LocalMux I__7268 (
            .O(N__43126),
            .I(N__43123));
    Odrv12 I__7267 (
            .O(N__43123),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22 ));
    InMux I__7266 (
            .O(N__43120),
            .I(N__43117));
    LocalMux I__7265 (
            .O(N__43117),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n7 ));
    InMux I__7264 (
            .O(N__43114),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15742 ));
    InMux I__7263 (
            .O(N__43111),
            .I(N__43108));
    LocalMux I__7262 (
            .O(N__43108),
            .I(N__43105));
    Span4Mux_v I__7261 (
            .O(N__43105),
            .I(N__43102));
    Odrv4 I__7260 (
            .O(N__43102),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n6 ));
    InMux I__7259 (
            .O(N__43099),
            .I(bfn_16_21_0_));
    InMux I__7258 (
            .O(N__43096),
            .I(N__43093));
    LocalMux I__7257 (
            .O(N__43093),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n5 ));
    InMux I__7256 (
            .O(N__43090),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15744 ));
    InMux I__7255 (
            .O(N__43087),
            .I(N__43084));
    LocalMux I__7254 (
            .O(N__43084),
            .I(N__43081));
    Span4Mux_v I__7253 (
            .O(N__43081),
            .I(N__43078));
    Odrv4 I__7252 (
            .O(N__43078),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4 ));
    InMux I__7251 (
            .O(N__43075),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15745 ));
    InMux I__7250 (
            .O(N__43072),
            .I(N__43069));
    LocalMux I__7249 (
            .O(N__43069),
            .I(N__43066));
    Span4Mux_v I__7248 (
            .O(N__43066),
            .I(N__43063));
    Odrv4 I__7247 (
            .O(N__43063),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n3 ));
    InMux I__7246 (
            .O(N__43060),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15746 ));
    InMux I__7245 (
            .O(N__43057),
            .I(N__43054));
    LocalMux I__7244 (
            .O(N__43054),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n2 ));
    InMux I__7243 (
            .O(N__43051),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15747 ));
    InMux I__7242 (
            .O(N__43048),
            .I(N__43045));
    LocalMux I__7241 (
            .O(N__43045),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725 ));
    CascadeMux I__7240 (
            .O(N__43042),
            .I(N__43038));
    CascadeMux I__7239 (
            .O(N__43041),
            .I(N__43035));
    InMux I__7238 (
            .O(N__43038),
            .I(N__43031));
    InMux I__7237 (
            .O(N__43035),
            .I(N__43026));
    InMux I__7236 (
            .O(N__43034),
            .I(N__43026));
    LocalMux I__7235 (
            .O(N__43031),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720 ));
    LocalMux I__7234 (
            .O(N__43026),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720 ));
    InMux I__7233 (
            .O(N__43021),
            .I(N__43018));
    LocalMux I__7232 (
            .O(N__43018),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15 ));
    InMux I__7231 (
            .O(N__43015),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15734 ));
    InMux I__7230 (
            .O(N__43012),
            .I(N__43009));
    LocalMux I__7229 (
            .O(N__43009),
            .I(N__43006));
    Odrv4 I__7228 (
            .O(N__43006),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n14 ));
    InMux I__7227 (
            .O(N__43003),
            .I(bfn_16_20_0_));
    InMux I__7226 (
            .O(N__43000),
            .I(N__42997));
    LocalMux I__7225 (
            .O(N__42997),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n13 ));
    InMux I__7224 (
            .O(N__42994),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15736 ));
    InMux I__7223 (
            .O(N__42991),
            .I(N__42988));
    LocalMux I__7222 (
            .O(N__42988),
            .I(N__42985));
    Odrv4 I__7221 (
            .O(N__42985),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n12 ));
    InMux I__7220 (
            .O(N__42982),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15737 ));
    InMux I__7219 (
            .O(N__42979),
            .I(N__42976));
    LocalMux I__7218 (
            .O(N__42976),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n11 ));
    InMux I__7217 (
            .O(N__42973),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15738 ));
    InMux I__7216 (
            .O(N__42970),
            .I(N__42967));
    LocalMux I__7215 (
            .O(N__42967),
            .I(N__42964));
    Odrv12 I__7214 (
            .O(N__42964),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10 ));
    InMux I__7213 (
            .O(N__42961),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15739 ));
    InMux I__7212 (
            .O(N__42958),
            .I(N__42955));
    LocalMux I__7211 (
            .O(N__42955),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n9 ));
    InMux I__7210 (
            .O(N__42952),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15740 ));
    InMux I__7209 (
            .O(N__42949),
            .I(N__42946));
    LocalMux I__7208 (
            .O(N__42946),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n8 ));
    InMux I__7207 (
            .O(N__42943),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15741 ));
    InMux I__7206 (
            .O(N__42940),
            .I(N__42937));
    LocalMux I__7205 (
            .O(N__42937),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n24 ));
    InMux I__7204 (
            .O(N__42934),
            .I(N__42931));
    LocalMux I__7203 (
            .O(N__42931),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n23 ));
    InMux I__7202 (
            .O(N__42928),
            .I(N__42925));
    LocalMux I__7201 (
            .O(N__42925),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n22 ));
    InMux I__7200 (
            .O(N__42922),
            .I(N__42919));
    LocalMux I__7199 (
            .O(N__42919),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752 ));
    InMux I__7198 (
            .O(N__42916),
            .I(N__42913));
    LocalMux I__7197 (
            .O(N__42913),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20 ));
    InMux I__7196 (
            .O(N__42910),
            .I(N__42907));
    LocalMux I__7195 (
            .O(N__42907),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19 ));
    InMux I__7194 (
            .O(N__42904),
            .I(N__42901));
    LocalMux I__7193 (
            .O(N__42901),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751 ));
    InMux I__7192 (
            .O(N__42898),
            .I(N__42895));
    LocalMux I__7191 (
            .O(N__42895),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17 ));
    InMux I__7190 (
            .O(N__42892),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15732 ));
    InMux I__7189 (
            .O(N__42889),
            .I(N__42886));
    LocalMux I__7188 (
            .O(N__42886),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n16 ));
    InMux I__7187 (
            .O(N__42883),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15733 ));
    InMux I__7186 (
            .O(N__42880),
            .I(N__42877));
    LocalMux I__7185 (
            .O(N__42877),
            .I(N__42874));
    Odrv4 I__7184 (
            .O(N__42874),
            .I(\foc.qCurrent_5 ));
    InMux I__7183 (
            .O(N__42871),
            .I(N__42868));
    LocalMux I__7182 (
            .O(N__42868),
            .I(N__42865));
    Odrv4 I__7181 (
            .O(N__42865),
            .I(\foc.qCurrent_9 ));
    InMux I__7180 (
            .O(N__42862),
            .I(N__42859));
    LocalMux I__7179 (
            .O(N__42859),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n30 ));
    InMux I__7178 (
            .O(N__42856),
            .I(N__42853));
    LocalMux I__7177 (
            .O(N__42853),
            .I(N__42850));
    Span4Mux_v I__7176 (
            .O(N__42850),
            .I(N__42846));
    CascadeMux I__7175 (
            .O(N__42849),
            .I(N__42843));
    Sp12to4 I__7174 (
            .O(N__42846),
            .I(N__42840));
    InMux I__7173 (
            .O(N__42843),
            .I(N__42837));
    Span12Mux_h I__7172 (
            .O(N__42840),
            .I(N__42834));
    LocalMux I__7171 (
            .O(N__42837),
            .I(N__42831));
    Odrv12 I__7170 (
            .O(N__42834),
            .I(\foc.u_DQ_Current_Control.n31 ));
    Odrv4 I__7169 (
            .O(N__42831),
            .I(\foc.u_DQ_Current_Control.n31 ));
    InMux I__7168 (
            .O(N__42826),
            .I(N__42823));
    LocalMux I__7167 (
            .O(N__42823),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n29 ));
    InMux I__7166 (
            .O(N__42820),
            .I(N__42817));
    LocalMux I__7165 (
            .O(N__42817),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n28 ));
    InMux I__7164 (
            .O(N__42814),
            .I(N__42811));
    LocalMux I__7163 (
            .O(N__42811),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753 ));
    InMux I__7162 (
            .O(N__42808),
            .I(N__42805));
    LocalMux I__7161 (
            .O(N__42805),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n26 ));
    InMux I__7160 (
            .O(N__42802),
            .I(N__42799));
    LocalMux I__7159 (
            .O(N__42799),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n25 ));
    InMux I__7158 (
            .O(N__42796),
            .I(N__42793));
    LocalMux I__7157 (
            .O(N__42793),
            .I(N__42790));
    Span4Mux_v I__7156 (
            .O(N__42790),
            .I(N__42786));
    InMux I__7155 (
            .O(N__42789),
            .I(N__42783));
    Span4Mux_v I__7154 (
            .O(N__42786),
            .I(N__42778));
    LocalMux I__7153 (
            .O(N__42783),
            .I(N__42778));
    Span4Mux_h I__7152 (
            .O(N__42778),
            .I(N__42775));
    Odrv4 I__7151 (
            .O(N__42775),
            .I(\foc.u_Park_Transform.n745 ));
    CascadeMux I__7150 (
            .O(N__42772),
            .I(N__42769));
    InMux I__7149 (
            .O(N__42769),
            .I(N__42766));
    LocalMux I__7148 (
            .O(N__42766),
            .I(\foc.u_Park_Transform.n697 ));
    InMux I__7147 (
            .O(N__42763),
            .I(N__42760));
    LocalMux I__7146 (
            .O(N__42760),
            .I(N__42757));
    Span4Mux_h I__7145 (
            .O(N__42757),
            .I(N__42754));
    Odrv4 I__7144 (
            .O(N__42754),
            .I(\foc.u_Park_Transform.n746_adj_2011 ));
    InMux I__7143 (
            .O(N__42751),
            .I(\foc.u_Park_Transform.n17051 ));
    InMux I__7142 (
            .O(N__42748),
            .I(\foc.u_Park_Transform.n747_adj_2012 ));
    CascadeMux I__7141 (
            .O(N__42745),
            .I(N__42742));
    InMux I__7140 (
            .O(N__42742),
            .I(N__42739));
    LocalMux I__7139 (
            .O(N__42739),
            .I(N__42736));
    Span4Mux_v I__7138 (
            .O(N__42736),
            .I(N__42733));
    Span4Mux_v I__7137 (
            .O(N__42733),
            .I(N__42730));
    Odrv4 I__7136 (
            .O(N__42730),
            .I(\foc.u_Park_Transform.n747_adj_2012_THRU_CO ));
    CascadeMux I__7135 (
            .O(N__42727),
            .I(\foc.u_Park_Transform.n6_cascade_ ));
    InMux I__7134 (
            .O(N__42724),
            .I(N__42721));
    LocalMux I__7133 (
            .O(N__42721),
            .I(N__42718));
    Span4Mux_v I__7132 (
            .O(N__42718),
            .I(N__42715));
    Sp12to4 I__7131 (
            .O(N__42715),
            .I(N__42711));
    InMux I__7130 (
            .O(N__42714),
            .I(N__42708));
    Odrv12 I__7129 (
            .O(N__42711),
            .I(\foc.Look_Up_Table_out1_1_2 ));
    LocalMux I__7128 (
            .O(N__42708),
            .I(\foc.Look_Up_Table_out1_1_2 ));
    CascadeMux I__7127 (
            .O(N__42703),
            .I(N__42693));
    CascadeMux I__7126 (
            .O(N__42702),
            .I(N__42689));
    CascadeMux I__7125 (
            .O(N__42701),
            .I(N__42685));
    CascadeMux I__7124 (
            .O(N__42700),
            .I(N__42680));
    CascadeMux I__7123 (
            .O(N__42699),
            .I(N__42677));
    CascadeMux I__7122 (
            .O(N__42698),
            .I(N__42674));
    CascadeMux I__7121 (
            .O(N__42697),
            .I(N__42671));
    CascadeMux I__7120 (
            .O(N__42696),
            .I(N__42667));
    InMux I__7119 (
            .O(N__42693),
            .I(N__42653));
    InMux I__7118 (
            .O(N__42692),
            .I(N__42653));
    InMux I__7117 (
            .O(N__42689),
            .I(N__42653));
    InMux I__7116 (
            .O(N__42688),
            .I(N__42653));
    InMux I__7115 (
            .O(N__42685),
            .I(N__42653));
    InMux I__7114 (
            .O(N__42684),
            .I(N__42653));
    InMux I__7113 (
            .O(N__42683),
            .I(N__42648));
    InMux I__7112 (
            .O(N__42680),
            .I(N__42648));
    InMux I__7111 (
            .O(N__42677),
            .I(N__42645));
    InMux I__7110 (
            .O(N__42674),
            .I(N__42634));
    InMux I__7109 (
            .O(N__42671),
            .I(N__42634));
    InMux I__7108 (
            .O(N__42670),
            .I(N__42634));
    InMux I__7107 (
            .O(N__42667),
            .I(N__42634));
    InMux I__7106 (
            .O(N__42666),
            .I(N__42634));
    LocalMux I__7105 (
            .O(N__42653),
            .I(N__42623));
    LocalMux I__7104 (
            .O(N__42648),
            .I(N__42623));
    LocalMux I__7103 (
            .O(N__42645),
            .I(N__42618));
    LocalMux I__7102 (
            .O(N__42634),
            .I(N__42618));
    InMux I__7101 (
            .O(N__42633),
            .I(N__42615));
    CascadeMux I__7100 (
            .O(N__42632),
            .I(N__42612));
    CascadeMux I__7099 (
            .O(N__42631),
            .I(N__42608));
    CascadeMux I__7098 (
            .O(N__42630),
            .I(N__42604));
    CascadeMux I__7097 (
            .O(N__42629),
            .I(N__42600));
    CascadeMux I__7096 (
            .O(N__42628),
            .I(N__42597));
    Span4Mux_h I__7095 (
            .O(N__42623),
            .I(N__42590));
    Span4Mux_h I__7094 (
            .O(N__42618),
            .I(N__42585));
    LocalMux I__7093 (
            .O(N__42615),
            .I(N__42585));
    InMux I__7092 (
            .O(N__42612),
            .I(N__42570));
    InMux I__7091 (
            .O(N__42611),
            .I(N__42570));
    InMux I__7090 (
            .O(N__42608),
            .I(N__42570));
    InMux I__7089 (
            .O(N__42607),
            .I(N__42570));
    InMux I__7088 (
            .O(N__42604),
            .I(N__42570));
    InMux I__7087 (
            .O(N__42603),
            .I(N__42570));
    InMux I__7086 (
            .O(N__42600),
            .I(N__42570));
    InMux I__7085 (
            .O(N__42597),
            .I(N__42567));
    CascadeMux I__7084 (
            .O(N__42596),
            .I(N__42564));
    CascadeMux I__7083 (
            .O(N__42595),
            .I(N__42560));
    CascadeMux I__7082 (
            .O(N__42594),
            .I(N__42556));
    CascadeMux I__7081 (
            .O(N__42593),
            .I(N__42552));
    Span4Mux_v I__7080 (
            .O(N__42590),
            .I(N__42549));
    Span4Mux_v I__7079 (
            .O(N__42585),
            .I(N__42542));
    LocalMux I__7078 (
            .O(N__42570),
            .I(N__42542));
    LocalMux I__7077 (
            .O(N__42567),
            .I(N__42542));
    InMux I__7076 (
            .O(N__42564),
            .I(N__42529));
    InMux I__7075 (
            .O(N__42563),
            .I(N__42529));
    InMux I__7074 (
            .O(N__42560),
            .I(N__42529));
    InMux I__7073 (
            .O(N__42559),
            .I(N__42529));
    InMux I__7072 (
            .O(N__42556),
            .I(N__42529));
    InMux I__7071 (
            .O(N__42555),
            .I(N__42529));
    InMux I__7070 (
            .O(N__42552),
            .I(N__42526));
    Odrv4 I__7069 (
            .O(N__42549),
            .I(\foc.u_Park_Transform.n595 ));
    Odrv4 I__7068 (
            .O(N__42542),
            .I(\foc.u_Park_Transform.n595 ));
    LocalMux I__7067 (
            .O(N__42529),
            .I(\foc.u_Park_Transform.n595 ));
    LocalMux I__7066 (
            .O(N__42526),
            .I(\foc.u_Park_Transform.n595 ));
    InMux I__7065 (
            .O(N__42517),
            .I(N__42511));
    InMux I__7064 (
            .O(N__42516),
            .I(N__42511));
    LocalMux I__7063 (
            .O(N__42511),
            .I(N__42508));
    Span4Mux_h I__7062 (
            .O(N__42508),
            .I(N__42504));
    InMux I__7061 (
            .O(N__42507),
            .I(N__42501));
    Odrv4 I__7060 (
            .O(N__42504),
            .I(n4));
    LocalMux I__7059 (
            .O(N__42501),
            .I(n4));
    InMux I__7058 (
            .O(N__42496),
            .I(N__42493));
    LocalMux I__7057 (
            .O(N__42493),
            .I(N__42490));
    Odrv12 I__7056 (
            .O(N__42490),
            .I(\foc.qCurrent_10 ));
    InMux I__7055 (
            .O(N__42487),
            .I(N__42484));
    LocalMux I__7054 (
            .O(N__42484),
            .I(N__42481));
    Odrv12 I__7053 (
            .O(N__42481),
            .I(\foc.qCurrent_7 ));
    CascadeMux I__7052 (
            .O(N__42478),
            .I(N__42475));
    InMux I__7051 (
            .O(N__42475),
            .I(N__42472));
    LocalMux I__7050 (
            .O(N__42472),
            .I(\foc.u_Park_Transform.n305 ));
    CascadeMux I__7049 (
            .O(N__42469),
            .I(N__42466));
    InMux I__7048 (
            .O(N__42466),
            .I(N__42463));
    LocalMux I__7047 (
            .O(N__42463),
            .I(N__42460));
    Odrv4 I__7046 (
            .O(N__42460),
            .I(\foc.u_Park_Transform.n351 ));
    InMux I__7045 (
            .O(N__42457),
            .I(\foc.u_Park_Transform.n17043 ));
    InMux I__7044 (
            .O(N__42454),
            .I(N__42451));
    LocalMux I__7043 (
            .O(N__42451),
            .I(\foc.u_Park_Transform.n354 ));
    CascadeMux I__7042 (
            .O(N__42448),
            .I(N__42445));
    InMux I__7041 (
            .O(N__42445),
            .I(N__42442));
    LocalMux I__7040 (
            .O(N__42442),
            .I(N__42439));
    Span4Mux_v I__7039 (
            .O(N__42439),
            .I(N__42436));
    Odrv4 I__7038 (
            .O(N__42436),
            .I(\foc.u_Park_Transform.n400 ));
    InMux I__7037 (
            .O(N__42433),
            .I(\foc.u_Park_Transform.n17044 ));
    CascadeMux I__7036 (
            .O(N__42430),
            .I(N__42427));
    InMux I__7035 (
            .O(N__42427),
            .I(N__42424));
    LocalMux I__7034 (
            .O(N__42424),
            .I(\foc.u_Park_Transform.n403 ));
    InMux I__7033 (
            .O(N__42421),
            .I(N__42418));
    LocalMux I__7032 (
            .O(N__42418),
            .I(N__42415));
    Odrv4 I__7031 (
            .O(N__42415),
            .I(\foc.u_Park_Transform.n449 ));
    InMux I__7030 (
            .O(N__42412),
            .I(bfn_16_14_0_));
    InMux I__7029 (
            .O(N__42409),
            .I(N__42406));
    LocalMux I__7028 (
            .O(N__42406),
            .I(\foc.u_Park_Transform.n452 ));
    CascadeMux I__7027 (
            .O(N__42403),
            .I(N__42400));
    InMux I__7026 (
            .O(N__42400),
            .I(N__42397));
    LocalMux I__7025 (
            .O(N__42397),
            .I(N__42394));
    Span4Mux_h I__7024 (
            .O(N__42394),
            .I(N__42391));
    Odrv4 I__7023 (
            .O(N__42391),
            .I(\foc.u_Park_Transform.n498 ));
    InMux I__7022 (
            .O(N__42388),
            .I(\foc.u_Park_Transform.n17046 ));
    CascadeMux I__7021 (
            .O(N__42385),
            .I(N__42382));
    InMux I__7020 (
            .O(N__42382),
            .I(N__42379));
    LocalMux I__7019 (
            .O(N__42379),
            .I(\foc.u_Park_Transform.n501 ));
    InMux I__7018 (
            .O(N__42376),
            .I(N__42373));
    LocalMux I__7017 (
            .O(N__42373),
            .I(N__42370));
    Odrv4 I__7016 (
            .O(N__42370),
            .I(\foc.u_Park_Transform.n547 ));
    InMux I__7015 (
            .O(N__42367),
            .I(\foc.u_Park_Transform.n17047 ));
    InMux I__7014 (
            .O(N__42364),
            .I(N__42361));
    LocalMux I__7013 (
            .O(N__42361),
            .I(\foc.u_Park_Transform.n550 ));
    CascadeMux I__7012 (
            .O(N__42358),
            .I(N__42355));
    InMux I__7011 (
            .O(N__42355),
            .I(N__42352));
    LocalMux I__7010 (
            .O(N__42352),
            .I(N__42349));
    Odrv4 I__7009 (
            .O(N__42349),
            .I(\foc.u_Park_Transform.n596 ));
    InMux I__7008 (
            .O(N__42346),
            .I(\foc.u_Park_Transform.n17048 ));
    CascadeMux I__7007 (
            .O(N__42343),
            .I(N__42340));
    InMux I__7006 (
            .O(N__42340),
            .I(N__42337));
    LocalMux I__7005 (
            .O(N__42337),
            .I(\foc.u_Park_Transform.n599 ));
    CascadeMux I__7004 (
            .O(N__42334),
            .I(N__42331));
    InMux I__7003 (
            .O(N__42331),
            .I(N__42328));
    LocalMux I__7002 (
            .O(N__42328),
            .I(N__42325));
    Odrv4 I__7001 (
            .O(N__42325),
            .I(\foc.u_Park_Transform.n645 ));
    InMux I__7000 (
            .O(N__42322),
            .I(\foc.u_Park_Transform.n17049 ));
    InMux I__6999 (
            .O(N__42319),
            .I(N__42316));
    LocalMux I__6998 (
            .O(N__42316),
            .I(\foc.u_Park_Transform.n648 ));
    CascadeMux I__6997 (
            .O(N__42313),
            .I(N__42310));
    InMux I__6996 (
            .O(N__42310),
            .I(N__42307));
    LocalMux I__6995 (
            .O(N__42307),
            .I(N__42304));
    Span4Mux_h I__6994 (
            .O(N__42304),
            .I(N__42301));
    Odrv4 I__6993 (
            .O(N__42301),
            .I(\foc.u_Park_Transform.n694 ));
    InMux I__6992 (
            .O(N__42298),
            .I(\foc.u_Park_Transform.n17050 ));
    InMux I__6991 (
            .O(N__42295),
            .I(N__42292));
    LocalMux I__6990 (
            .O(N__42292),
            .I(N__42288));
    InMux I__6989 (
            .O(N__42291),
            .I(N__42285));
    Span4Mux_v I__6988 (
            .O(N__42288),
            .I(N__42282));
    LocalMux I__6987 (
            .O(N__42285),
            .I(N__42279));
    Span4Mux_h I__6986 (
            .O(N__42282),
            .I(N__42276));
    Span4Mux_v I__6985 (
            .O(N__42279),
            .I(N__42273));
    Odrv4 I__6984 (
            .O(N__42276),
            .I(\foc.u_Park_Transform.n749 ));
    Odrv4 I__6983 (
            .O(N__42273),
            .I(\foc.u_Park_Transform.n749 ));
    CascadeMux I__6982 (
            .O(N__42268),
            .I(N__42265));
    InMux I__6981 (
            .O(N__42265),
            .I(N__42262));
    LocalMux I__6980 (
            .O(N__42262),
            .I(N__42259));
    Odrv12 I__6979 (
            .O(N__42259),
            .I(\foc.u_Park_Transform.n700_adj_2141 ));
    InMux I__6978 (
            .O(N__42256),
            .I(N__42253));
    LocalMux I__6977 (
            .O(N__42253),
            .I(N__42250));
    Span4Mux_h I__6976 (
            .O(N__42250),
            .I(N__42247));
    Odrv4 I__6975 (
            .O(N__42247),
            .I(\foc.u_Park_Transform.n750 ));
    InMux I__6974 (
            .O(N__42244),
            .I(\foc.u_Park_Transform.n17219 ));
    InMux I__6973 (
            .O(N__42241),
            .I(\foc.u_Park_Transform.n751_adj_2142 ));
    CascadeMux I__6972 (
            .O(N__42238),
            .I(N__42235));
    InMux I__6971 (
            .O(N__42235),
            .I(N__42232));
    LocalMux I__6970 (
            .O(N__42232),
            .I(N__42229));
    Span4Mux_h I__6969 (
            .O(N__42229),
            .I(N__42226));
    Odrv4 I__6968 (
            .O(N__42226),
            .I(\foc.u_Park_Transform.n751_adj_2142_THRU_CO ));
    CascadeMux I__6967 (
            .O(N__42223),
            .I(N__42212));
    CascadeMux I__6966 (
            .O(N__42222),
            .I(N__42208));
    CascadeMux I__6965 (
            .O(N__42221),
            .I(N__42204));
    CascadeMux I__6964 (
            .O(N__42220),
            .I(N__42200));
    CascadeMux I__6963 (
            .O(N__42219),
            .I(N__42197));
    CascadeMux I__6962 (
            .O(N__42218),
            .I(N__42194));
    CascadeMux I__6961 (
            .O(N__42217),
            .I(N__42191));
    CascadeMux I__6960 (
            .O(N__42216),
            .I(N__42187));
    CascadeMux I__6959 (
            .O(N__42215),
            .I(N__42179));
    InMux I__6958 (
            .O(N__42212),
            .I(N__42164));
    InMux I__6957 (
            .O(N__42211),
            .I(N__42164));
    InMux I__6956 (
            .O(N__42208),
            .I(N__42164));
    InMux I__6955 (
            .O(N__42207),
            .I(N__42164));
    InMux I__6954 (
            .O(N__42204),
            .I(N__42164));
    InMux I__6953 (
            .O(N__42203),
            .I(N__42164));
    InMux I__6952 (
            .O(N__42200),
            .I(N__42164));
    InMux I__6951 (
            .O(N__42197),
            .I(N__42161));
    InMux I__6950 (
            .O(N__42194),
            .I(N__42150));
    InMux I__6949 (
            .O(N__42191),
            .I(N__42150));
    InMux I__6948 (
            .O(N__42190),
            .I(N__42150));
    InMux I__6947 (
            .O(N__42187),
            .I(N__42150));
    InMux I__6946 (
            .O(N__42186),
            .I(N__42150));
    CascadeMux I__6945 (
            .O(N__42185),
            .I(N__42147));
    CascadeMux I__6944 (
            .O(N__42184),
            .I(N__42143));
    CascadeMux I__6943 (
            .O(N__42183),
            .I(N__42139));
    InMux I__6942 (
            .O(N__42182),
            .I(N__42131));
    InMux I__6941 (
            .O(N__42179),
            .I(N__42127));
    LocalMux I__6940 (
            .O(N__42164),
            .I(N__42120));
    LocalMux I__6939 (
            .O(N__42161),
            .I(N__42120));
    LocalMux I__6938 (
            .O(N__42150),
            .I(N__42120));
    InMux I__6937 (
            .O(N__42147),
            .I(N__42107));
    InMux I__6936 (
            .O(N__42146),
            .I(N__42107));
    InMux I__6935 (
            .O(N__42143),
            .I(N__42107));
    InMux I__6934 (
            .O(N__42142),
            .I(N__42107));
    InMux I__6933 (
            .O(N__42139),
            .I(N__42107));
    InMux I__6932 (
            .O(N__42138),
            .I(N__42107));
    CascadeMux I__6931 (
            .O(N__42137),
            .I(N__42104));
    CascadeMux I__6930 (
            .O(N__42136),
            .I(N__42100));
    CascadeMux I__6929 (
            .O(N__42135),
            .I(N__42096));
    CascadeMux I__6928 (
            .O(N__42134),
            .I(N__42092));
    LocalMux I__6927 (
            .O(N__42131),
            .I(N__42088));
    InMux I__6926 (
            .O(N__42130),
            .I(N__42085));
    LocalMux I__6925 (
            .O(N__42127),
            .I(N__42082));
    Span4Mux_v I__6924 (
            .O(N__42120),
            .I(N__42077));
    LocalMux I__6923 (
            .O(N__42107),
            .I(N__42077));
    InMux I__6922 (
            .O(N__42104),
            .I(N__42060));
    InMux I__6921 (
            .O(N__42103),
            .I(N__42060));
    InMux I__6920 (
            .O(N__42100),
            .I(N__42060));
    InMux I__6919 (
            .O(N__42099),
            .I(N__42060));
    InMux I__6918 (
            .O(N__42096),
            .I(N__42060));
    InMux I__6917 (
            .O(N__42095),
            .I(N__42060));
    InMux I__6916 (
            .O(N__42092),
            .I(N__42060));
    InMux I__6915 (
            .O(N__42091),
            .I(N__42060));
    Span4Mux_v I__6914 (
            .O(N__42088),
            .I(N__42057));
    LocalMux I__6913 (
            .O(N__42085),
            .I(N__42054));
    Span4Mux_v I__6912 (
            .O(N__42082),
            .I(N__42047));
    Span4Mux_v I__6911 (
            .O(N__42077),
            .I(N__42047));
    LocalMux I__6910 (
            .O(N__42060),
            .I(N__42047));
    Odrv4 I__6909 (
            .O(N__42057),
            .I(\foc.u_Park_Transform.n598 ));
    Odrv12 I__6908 (
            .O(N__42054),
            .I(\foc.u_Park_Transform.n598 ));
    Odrv4 I__6907 (
            .O(N__42047),
            .I(\foc.u_Park_Transform.n598 ));
    InMux I__6906 (
            .O(N__42040),
            .I(N__42037));
    LocalMux I__6905 (
            .O(N__42037),
            .I(N__42034));
    Odrv4 I__6904 (
            .O(N__42034),
            .I(\foc.u_Park_Transform.n57 ));
    InMux I__6903 (
            .O(N__42031),
            .I(N__42028));
    LocalMux I__6902 (
            .O(N__42028),
            .I(\foc.u_Park_Transform.n60 ));
    CascadeMux I__6901 (
            .O(N__42025),
            .I(N__42022));
    InMux I__6900 (
            .O(N__42022),
            .I(N__42019));
    LocalMux I__6899 (
            .O(N__42019),
            .I(N__42016));
    Span4Mux_v I__6898 (
            .O(N__42016),
            .I(N__42013));
    Odrv4 I__6897 (
            .O(N__42013),
            .I(\foc.u_Park_Transform.n106 ));
    InMux I__6896 (
            .O(N__42010),
            .I(\foc.u_Park_Transform.n17038 ));
    CascadeMux I__6895 (
            .O(N__42007),
            .I(N__42004));
    InMux I__6894 (
            .O(N__42004),
            .I(N__42001));
    LocalMux I__6893 (
            .O(N__42001),
            .I(\foc.u_Park_Transform.n109 ));
    InMux I__6892 (
            .O(N__41998),
            .I(N__41995));
    LocalMux I__6891 (
            .O(N__41995),
            .I(N__41992));
    Odrv4 I__6890 (
            .O(N__41992),
            .I(\foc.u_Park_Transform.n155 ));
    InMux I__6889 (
            .O(N__41989),
            .I(\foc.u_Park_Transform.n17039 ));
    InMux I__6888 (
            .O(N__41986),
            .I(N__41983));
    LocalMux I__6887 (
            .O(N__41983),
            .I(\foc.u_Park_Transform.n158 ));
    CascadeMux I__6886 (
            .O(N__41980),
            .I(N__41977));
    InMux I__6885 (
            .O(N__41977),
            .I(N__41974));
    LocalMux I__6884 (
            .O(N__41974),
            .I(N__41971));
    Odrv4 I__6883 (
            .O(N__41971),
            .I(\foc.u_Park_Transform.n204 ));
    InMux I__6882 (
            .O(N__41968),
            .I(\foc.u_Park_Transform.n17040 ));
    CascadeMux I__6881 (
            .O(N__41965),
            .I(N__41962));
    InMux I__6880 (
            .O(N__41962),
            .I(N__41959));
    LocalMux I__6879 (
            .O(N__41959),
            .I(\foc.u_Park_Transform.n207 ));
    CascadeMux I__6878 (
            .O(N__41956),
            .I(N__41953));
    InMux I__6877 (
            .O(N__41953),
            .I(N__41950));
    LocalMux I__6876 (
            .O(N__41950),
            .I(N__41947));
    Odrv4 I__6875 (
            .O(N__41947),
            .I(\foc.u_Park_Transform.n253 ));
    InMux I__6874 (
            .O(N__41944),
            .I(\foc.u_Park_Transform.n17041 ));
    InMux I__6873 (
            .O(N__41941),
            .I(N__41938));
    LocalMux I__6872 (
            .O(N__41938),
            .I(\foc.u_Park_Transform.n256 ));
    CascadeMux I__6871 (
            .O(N__41935),
            .I(N__41932));
    InMux I__6870 (
            .O(N__41932),
            .I(N__41929));
    LocalMux I__6869 (
            .O(N__41929),
            .I(N__41926));
    Span4Mux_h I__6868 (
            .O(N__41926),
            .I(N__41923));
    Odrv4 I__6867 (
            .O(N__41923),
            .I(\foc.u_Park_Transform.n302 ));
    InMux I__6866 (
            .O(N__41920),
            .I(\foc.u_Park_Transform.n17042 ));
    InMux I__6865 (
            .O(N__41917),
            .I(N__41914));
    LocalMux I__6864 (
            .O(N__41914),
            .I(N__41911));
    Odrv4 I__6863 (
            .O(N__41911),
            .I(\foc.u_Park_Transform.n354_adj_2133 ));
    InMux I__6862 (
            .O(N__41908),
            .I(\foc.u_Park_Transform.n17211 ));
    InMux I__6861 (
            .O(N__41905),
            .I(N__41902));
    LocalMux I__6860 (
            .O(N__41902),
            .I(N__41899));
    Odrv12 I__6859 (
            .O(N__41899),
            .I(\foc.u_Park_Transform.n357_adj_2151 ));
    CascadeMux I__6858 (
            .O(N__41896),
            .I(N__41893));
    InMux I__6857 (
            .O(N__41893),
            .I(N__41890));
    LocalMux I__6856 (
            .O(N__41890),
            .I(N__41887));
    Span4Mux_v I__6855 (
            .O(N__41887),
            .I(N__41884));
    Odrv4 I__6854 (
            .O(N__41884),
            .I(\foc.u_Park_Transform.n403_adj_2132 ));
    InMux I__6853 (
            .O(N__41881),
            .I(\foc.u_Park_Transform.n17212 ));
    CascadeMux I__6852 (
            .O(N__41878),
            .I(N__41875));
    InMux I__6851 (
            .O(N__41875),
            .I(N__41872));
    LocalMux I__6850 (
            .O(N__41872),
            .I(N__41869));
    Span4Mux_h I__6849 (
            .O(N__41869),
            .I(N__41866));
    Odrv4 I__6848 (
            .O(N__41866),
            .I(\foc.u_Park_Transform.n406_adj_2150 ));
    InMux I__6847 (
            .O(N__41863),
            .I(N__41860));
    LocalMux I__6846 (
            .O(N__41860),
            .I(N__41857));
    Odrv4 I__6845 (
            .O(N__41857),
            .I(\foc.u_Park_Transform.n452_adj_2131 ));
    InMux I__6844 (
            .O(N__41854),
            .I(bfn_16_12_0_));
    InMux I__6843 (
            .O(N__41851),
            .I(N__41848));
    LocalMux I__6842 (
            .O(N__41848),
            .I(N__41845));
    Odrv12 I__6841 (
            .O(N__41845),
            .I(\foc.u_Park_Transform.n455_adj_2148 ));
    CascadeMux I__6840 (
            .O(N__41842),
            .I(N__41839));
    InMux I__6839 (
            .O(N__41839),
            .I(N__41836));
    LocalMux I__6838 (
            .O(N__41836),
            .I(N__41833));
    Odrv4 I__6837 (
            .O(N__41833),
            .I(\foc.u_Park_Transform.n501_adj_2130 ));
    InMux I__6836 (
            .O(N__41830),
            .I(\foc.u_Park_Transform.n17214 ));
    CascadeMux I__6835 (
            .O(N__41827),
            .I(N__41824));
    InMux I__6834 (
            .O(N__41824),
            .I(N__41821));
    LocalMux I__6833 (
            .O(N__41821),
            .I(N__41818));
    Odrv4 I__6832 (
            .O(N__41818),
            .I(\foc.u_Park_Transform.n504_adj_2147 ));
    InMux I__6831 (
            .O(N__41815),
            .I(N__41812));
    LocalMux I__6830 (
            .O(N__41812),
            .I(N__41809));
    Span4Mux_h I__6829 (
            .O(N__41809),
            .I(N__41806));
    Odrv4 I__6828 (
            .O(N__41806),
            .I(\foc.u_Park_Transform.n550_adj_2129 ));
    InMux I__6827 (
            .O(N__41803),
            .I(\foc.u_Park_Transform.n17215 ));
    InMux I__6826 (
            .O(N__41800),
            .I(N__41797));
    LocalMux I__6825 (
            .O(N__41797),
            .I(N__41794));
    Odrv12 I__6824 (
            .O(N__41794),
            .I(\foc.u_Park_Transform.n553_adj_2146 ));
    InMux I__6823 (
            .O(N__41791),
            .I(N__41788));
    LocalMux I__6822 (
            .O(N__41788),
            .I(N__41785));
    Odrv12 I__6821 (
            .O(N__41785),
            .I(\foc.u_Park_Transform.n599_adj_2128 ));
    InMux I__6820 (
            .O(N__41782),
            .I(\foc.u_Park_Transform.n17216 ));
    InMux I__6819 (
            .O(N__41779),
            .I(N__41776));
    LocalMux I__6818 (
            .O(N__41776),
            .I(N__41773));
    Odrv12 I__6817 (
            .O(N__41773),
            .I(\foc.u_Park_Transform.n602_adj_2144 ));
    InMux I__6816 (
            .O(N__41770),
            .I(N__41767));
    LocalMux I__6815 (
            .O(N__41767),
            .I(N__41764));
    Odrv12 I__6814 (
            .O(N__41764),
            .I(\foc.u_Park_Transform.n648_adj_2124 ));
    InMux I__6813 (
            .O(N__41761),
            .I(\foc.u_Park_Transform.n17217 ));
    InMux I__6812 (
            .O(N__41758),
            .I(N__41755));
    LocalMux I__6811 (
            .O(N__41755),
            .I(N__41752));
    Odrv4 I__6810 (
            .O(N__41752),
            .I(\foc.u_Park_Transform.n651_adj_2143 ));
    CascadeMux I__6809 (
            .O(N__41749),
            .I(N__41746));
    InMux I__6808 (
            .O(N__41746),
            .I(N__41743));
    LocalMux I__6807 (
            .O(N__41743),
            .I(N__41740));
    Odrv12 I__6806 (
            .O(N__41740),
            .I(\foc.u_Park_Transform.n697_adj_2121 ));
    InMux I__6805 (
            .O(N__41737),
            .I(\foc.u_Park_Transform.n17218 ));
    InMux I__6804 (
            .O(N__41734),
            .I(N__41731));
    LocalMux I__6803 (
            .O(N__41731),
            .I(N__41728));
    Span4Mux_v I__6802 (
            .O(N__41728),
            .I(N__41725));
    Odrv4 I__6801 (
            .O(N__41725),
            .I(\foc.dCurrent_27 ));
    InMux I__6800 (
            .O(N__41722),
            .I(N__41719));
    LocalMux I__6799 (
            .O(N__41719),
            .I(N__41716));
    Sp12to4 I__6798 (
            .O(N__41716),
            .I(N__41713));
    Odrv12 I__6797 (
            .O(N__41713),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n6 ));
    InMux I__6796 (
            .O(N__41710),
            .I(N__41704));
    CascadeMux I__6795 (
            .O(N__41709),
            .I(N__41701));
    CascadeMux I__6794 (
            .O(N__41708),
            .I(N__41697));
    CascadeMux I__6793 (
            .O(N__41707),
            .I(N__41693));
    LocalMux I__6792 (
            .O(N__41704),
            .I(N__41682));
    InMux I__6791 (
            .O(N__41701),
            .I(N__41669));
    InMux I__6790 (
            .O(N__41700),
            .I(N__41669));
    InMux I__6789 (
            .O(N__41697),
            .I(N__41669));
    InMux I__6788 (
            .O(N__41696),
            .I(N__41669));
    InMux I__6787 (
            .O(N__41693),
            .I(N__41669));
    InMux I__6786 (
            .O(N__41692),
            .I(N__41669));
    CascadeMux I__6785 (
            .O(N__41691),
            .I(N__41663));
    CascadeMux I__6784 (
            .O(N__41690),
            .I(N__41657));
    CascadeMux I__6783 (
            .O(N__41689),
            .I(N__41654));
    CascadeMux I__6782 (
            .O(N__41688),
            .I(N__41648));
    CascadeMux I__6781 (
            .O(N__41687),
            .I(N__41644));
    CascadeMux I__6780 (
            .O(N__41686),
            .I(N__41640));
    CascadeMux I__6779 (
            .O(N__41685),
            .I(N__41635));
    Span4Mux_v I__6778 (
            .O(N__41682),
            .I(N__41630));
    LocalMux I__6777 (
            .O(N__41669),
            .I(N__41630));
    InMux I__6776 (
            .O(N__41668),
            .I(N__41621));
    InMux I__6775 (
            .O(N__41667),
            .I(N__41621));
    InMux I__6774 (
            .O(N__41666),
            .I(N__41621));
    InMux I__6773 (
            .O(N__41663),
            .I(N__41621));
    InMux I__6772 (
            .O(N__41662),
            .I(N__41612));
    InMux I__6771 (
            .O(N__41661),
            .I(N__41612));
    InMux I__6770 (
            .O(N__41660),
            .I(N__41612));
    InMux I__6769 (
            .O(N__41657),
            .I(N__41612));
    InMux I__6768 (
            .O(N__41654),
            .I(N__41609));
    CascadeMux I__6767 (
            .O(N__41653),
            .I(N__41605));
    CascadeMux I__6766 (
            .O(N__41652),
            .I(N__41601));
    CascadeMux I__6765 (
            .O(N__41651),
            .I(N__41597));
    InMux I__6764 (
            .O(N__41648),
            .I(N__41584));
    InMux I__6763 (
            .O(N__41647),
            .I(N__41584));
    InMux I__6762 (
            .O(N__41644),
            .I(N__41584));
    InMux I__6761 (
            .O(N__41643),
            .I(N__41584));
    InMux I__6760 (
            .O(N__41640),
            .I(N__41584));
    InMux I__6759 (
            .O(N__41639),
            .I(N__41584));
    InMux I__6758 (
            .O(N__41638),
            .I(N__41579));
    InMux I__6757 (
            .O(N__41635),
            .I(N__41579));
    Span4Mux_h I__6756 (
            .O(N__41630),
            .I(N__41572));
    LocalMux I__6755 (
            .O(N__41621),
            .I(N__41572));
    LocalMux I__6754 (
            .O(N__41612),
            .I(N__41572));
    LocalMux I__6753 (
            .O(N__41609),
            .I(N__41569));
    InMux I__6752 (
            .O(N__41608),
            .I(N__41556));
    InMux I__6751 (
            .O(N__41605),
            .I(N__41556));
    InMux I__6750 (
            .O(N__41604),
            .I(N__41556));
    InMux I__6749 (
            .O(N__41601),
            .I(N__41556));
    InMux I__6748 (
            .O(N__41600),
            .I(N__41556));
    InMux I__6747 (
            .O(N__41597),
            .I(N__41556));
    LocalMux I__6746 (
            .O(N__41584),
            .I(N__41551));
    LocalMux I__6745 (
            .O(N__41579),
            .I(N__41551));
    Odrv4 I__6744 (
            .O(N__41572),
            .I(\foc.u_Park_Transform.n601 ));
    Odrv12 I__6743 (
            .O(N__41569),
            .I(\foc.u_Park_Transform.n601 ));
    LocalMux I__6742 (
            .O(N__41556),
            .I(\foc.u_Park_Transform.n601 ));
    Odrv4 I__6741 (
            .O(N__41551),
            .I(\foc.u_Park_Transform.n601 ));
    CascadeMux I__6740 (
            .O(N__41542),
            .I(N__41539));
    InMux I__6739 (
            .O(N__41539),
            .I(N__41536));
    LocalMux I__6738 (
            .O(N__41536),
            .I(N__41533));
    Odrv4 I__6737 (
            .O(N__41533),
            .I(\foc.u_Park_Transform.n60_adj_2140 ));
    InMux I__6736 (
            .O(N__41530),
            .I(N__41527));
    LocalMux I__6735 (
            .O(N__41527),
            .I(N__41524));
    Odrv4 I__6734 (
            .O(N__41524),
            .I(\foc.u_Park_Transform.n63_adj_2158 ));
    CascadeMux I__6733 (
            .O(N__41521),
            .I(N__41518));
    InMux I__6732 (
            .O(N__41518),
            .I(N__41515));
    LocalMux I__6731 (
            .O(N__41515),
            .I(N__41512));
    Odrv4 I__6730 (
            .O(N__41512),
            .I(\foc.u_Park_Transform.n109_adj_2139 ));
    InMux I__6729 (
            .O(N__41509),
            .I(\foc.u_Park_Transform.n17206 ));
    CascadeMux I__6728 (
            .O(N__41506),
            .I(N__41503));
    InMux I__6727 (
            .O(N__41503),
            .I(N__41500));
    LocalMux I__6726 (
            .O(N__41500),
            .I(N__41497));
    Odrv4 I__6725 (
            .O(N__41497),
            .I(\foc.u_Park_Transform.n112_adj_2157 ));
    InMux I__6724 (
            .O(N__41494),
            .I(N__41491));
    LocalMux I__6723 (
            .O(N__41491),
            .I(N__41488));
    Odrv12 I__6722 (
            .O(N__41488),
            .I(\foc.u_Park_Transform.n158_adj_2137 ));
    InMux I__6721 (
            .O(N__41485),
            .I(\foc.u_Park_Transform.n17207 ));
    InMux I__6720 (
            .O(N__41482),
            .I(N__41479));
    LocalMux I__6719 (
            .O(N__41479),
            .I(N__41476));
    Odrv4 I__6718 (
            .O(N__41476),
            .I(\foc.u_Park_Transform.n161_adj_2156 ));
    CascadeMux I__6717 (
            .O(N__41473),
            .I(N__41470));
    InMux I__6716 (
            .O(N__41470),
            .I(N__41467));
    LocalMux I__6715 (
            .O(N__41467),
            .I(N__41464));
    Odrv4 I__6714 (
            .O(N__41464),
            .I(\foc.u_Park_Transform.n207_adj_2136 ));
    InMux I__6713 (
            .O(N__41461),
            .I(\foc.u_Park_Transform.n17208 ));
    CascadeMux I__6712 (
            .O(N__41458),
            .I(N__41455));
    InMux I__6711 (
            .O(N__41455),
            .I(N__41452));
    LocalMux I__6710 (
            .O(N__41452),
            .I(N__41449));
    Odrv4 I__6709 (
            .O(N__41449),
            .I(\foc.u_Park_Transform.n210_adj_2155 ));
    InMux I__6708 (
            .O(N__41446),
            .I(N__41443));
    LocalMux I__6707 (
            .O(N__41443),
            .I(N__41440));
    Span4Mux_h I__6706 (
            .O(N__41440),
            .I(N__41437));
    Odrv4 I__6705 (
            .O(N__41437),
            .I(\foc.u_Park_Transform.n256_adj_2135 ));
    InMux I__6704 (
            .O(N__41434),
            .I(\foc.u_Park_Transform.n17209 ));
    InMux I__6703 (
            .O(N__41431),
            .I(N__41428));
    LocalMux I__6702 (
            .O(N__41428),
            .I(N__41425));
    Odrv12 I__6701 (
            .O(N__41425),
            .I(\foc.u_Park_Transform.n259_adj_2154 ));
    CascadeMux I__6700 (
            .O(N__41422),
            .I(N__41419));
    InMux I__6699 (
            .O(N__41419),
            .I(N__41416));
    LocalMux I__6698 (
            .O(N__41416),
            .I(N__41413));
    Span4Mux_v I__6697 (
            .O(N__41413),
            .I(N__41410));
    Odrv4 I__6696 (
            .O(N__41410),
            .I(\foc.u_Park_Transform.n305_adj_2134 ));
    InMux I__6695 (
            .O(N__41407),
            .I(\foc.u_Park_Transform.n17210 ));
    CascadeMux I__6694 (
            .O(N__41404),
            .I(N__41401));
    InMux I__6693 (
            .O(N__41401),
            .I(N__41398));
    LocalMux I__6692 (
            .O(N__41398),
            .I(N__41395));
    Odrv12 I__6691 (
            .O(N__41395),
            .I(\foc.u_Park_Transform.n308_adj_2153 ));
    InMux I__6690 (
            .O(N__41392),
            .I(N__41388));
    InMux I__6689 (
            .O(N__41391),
            .I(N__41385));
    LocalMux I__6688 (
            .O(N__41388),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18 ));
    LocalMux I__6687 (
            .O(N__41385),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18 ));
    InMux I__6686 (
            .O(N__41380),
            .I(N__41374));
    InMux I__6685 (
            .O(N__41379),
            .I(N__41374));
    LocalMux I__6684 (
            .O(N__41374),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25 ));
    InMux I__6683 (
            .O(N__41371),
            .I(N__41368));
    LocalMux I__6682 (
            .O(N__41368),
            .I(N__41364));
    InMux I__6681 (
            .O(N__41367),
            .I(N__41361));
    Odrv4 I__6680 (
            .O(N__41364),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17 ));
    LocalMux I__6679 (
            .O(N__41361),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17 ));
    InMux I__6678 (
            .O(N__41356),
            .I(N__41350));
    InMux I__6677 (
            .O(N__41355),
            .I(N__41350));
    LocalMux I__6676 (
            .O(N__41350),
            .I(N__41347));
    Odrv4 I__6675 (
            .O(N__41347),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24 ));
    InMux I__6674 (
            .O(N__41344),
            .I(N__41341));
    LocalMux I__6673 (
            .O(N__41341),
            .I(N__41338));
    Odrv4 I__6672 (
            .O(N__41338),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623 ));
    InMux I__6671 (
            .O(N__41335),
            .I(N__41332));
    LocalMux I__6670 (
            .O(N__41332),
            .I(N__41329));
    Odrv4 I__6669 (
            .O(N__41329),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638 ));
    InMux I__6668 (
            .O(N__41326),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18088 ));
    CascadeMux I__6667 (
            .O(N__41323),
            .I(N__41320));
    InMux I__6666 (
            .O(N__41320),
            .I(N__41317));
    LocalMux I__6665 (
            .O(N__41317),
            .I(N__41314));
    Odrv12 I__6664 (
            .O(N__41314),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622 ));
    CascadeMux I__6663 (
            .O(N__41311),
            .I(N__41308));
    InMux I__6662 (
            .O(N__41308),
            .I(N__41305));
    LocalMux I__6661 (
            .O(N__41305),
            .I(N__41302));
    Odrv4 I__6660 (
            .O(N__41302),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637 ));
    InMux I__6659 (
            .O(N__41299),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18089 ));
    CascadeMux I__6658 (
            .O(N__41296),
            .I(N__41293));
    InMux I__6657 (
            .O(N__41293),
            .I(N__41290));
    LocalMux I__6656 (
            .O(N__41290),
            .I(N__41287));
    Odrv12 I__6655 (
            .O(N__41287),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621 ));
    InMux I__6654 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__6653 (
            .O(N__41281),
            .I(N__41278));
    Span12Mux_v I__6652 (
            .O(N__41278),
            .I(N__41275));
    Odrv12 I__6651 (
            .O(N__41275),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635 ));
    InMux I__6650 (
            .O(N__41272),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18090 ));
    InMux I__6649 (
            .O(N__41269),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636 ));
    CascadeMux I__6648 (
            .O(N__41266),
            .I(N__41263));
    InMux I__6647 (
            .O(N__41263),
            .I(N__41260));
    LocalMux I__6646 (
            .O(N__41260),
            .I(N__41257));
    Span4Mux_h I__6645 (
            .O(N__41257),
            .I(N__41254));
    Odrv4 I__6644 (
            .O(N__41254),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO ));
    InMux I__6643 (
            .O(N__41251),
            .I(N__41245));
    InMux I__6642 (
            .O(N__41250),
            .I(N__41245));
    LocalMux I__6641 (
            .O(N__41245),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16 ));
    InMux I__6640 (
            .O(N__41242),
            .I(N__41238));
    InMux I__6639 (
            .O(N__41241),
            .I(N__41235));
    LocalMux I__6638 (
            .O(N__41238),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20 ));
    LocalMux I__6637 (
            .O(N__41235),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20 ));
    InMux I__6636 (
            .O(N__41230),
            .I(N__41227));
    LocalMux I__6635 (
            .O(N__41227),
            .I(N__41224));
    Odrv12 I__6634 (
            .O(N__41224),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631 ));
    CascadeMux I__6633 (
            .O(N__41221),
            .I(N__41218));
    InMux I__6632 (
            .O(N__41218),
            .I(N__41215));
    LocalMux I__6631 (
            .O(N__41215),
            .I(N__41212));
    Odrv4 I__6630 (
            .O(N__41212),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646 ));
    InMux I__6629 (
            .O(N__41209),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18080 ));
    CascadeMux I__6628 (
            .O(N__41206),
            .I(N__41203));
    InMux I__6627 (
            .O(N__41203),
            .I(N__41200));
    LocalMux I__6626 (
            .O(N__41200),
            .I(N__41197));
    Odrv4 I__6625 (
            .O(N__41197),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630 ));
    InMux I__6624 (
            .O(N__41194),
            .I(N__41191));
    LocalMux I__6623 (
            .O(N__41191),
            .I(N__41188));
    Odrv4 I__6622 (
            .O(N__41188),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645 ));
    InMux I__6621 (
            .O(N__41185),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18081 ));
    CascadeMux I__6620 (
            .O(N__41182),
            .I(N__41179));
    InMux I__6619 (
            .O(N__41179),
            .I(N__41176));
    LocalMux I__6618 (
            .O(N__41176),
            .I(N__41173));
    Odrv4 I__6617 (
            .O(N__41173),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629 ));
    CascadeMux I__6616 (
            .O(N__41170),
            .I(N__41167));
    InMux I__6615 (
            .O(N__41167),
            .I(N__41164));
    LocalMux I__6614 (
            .O(N__41164),
            .I(N__41161));
    Odrv4 I__6613 (
            .O(N__41161),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644 ));
    InMux I__6612 (
            .O(N__41158),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18082 ));
    InMux I__6611 (
            .O(N__41155),
            .I(N__41152));
    LocalMux I__6610 (
            .O(N__41152),
            .I(N__41149));
    Odrv12 I__6609 (
            .O(N__41149),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628 ));
    InMux I__6608 (
            .O(N__41146),
            .I(N__41143));
    LocalMux I__6607 (
            .O(N__41143),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643 ));
    InMux I__6606 (
            .O(N__41140),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18083 ));
    InMux I__6605 (
            .O(N__41137),
            .I(N__41134));
    LocalMux I__6604 (
            .O(N__41134),
            .I(N__41131));
    Span4Mux_v I__6603 (
            .O(N__41131),
            .I(N__41128));
    Odrv4 I__6602 (
            .O(N__41128),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627 ));
    CascadeMux I__6601 (
            .O(N__41125),
            .I(N__41122));
    InMux I__6600 (
            .O(N__41122),
            .I(N__41119));
    LocalMux I__6599 (
            .O(N__41119),
            .I(N__41116));
    Odrv4 I__6598 (
            .O(N__41116),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642 ));
    InMux I__6597 (
            .O(N__41113),
            .I(bfn_15_26_0_));
    CascadeMux I__6596 (
            .O(N__41110),
            .I(N__41107));
    InMux I__6595 (
            .O(N__41107),
            .I(N__41104));
    LocalMux I__6594 (
            .O(N__41104),
            .I(N__41101));
    Odrv4 I__6593 (
            .O(N__41101),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626 ));
    InMux I__6592 (
            .O(N__41098),
            .I(N__41095));
    LocalMux I__6591 (
            .O(N__41095),
            .I(N__41092));
    Odrv4 I__6590 (
            .O(N__41092),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641 ));
    InMux I__6589 (
            .O(N__41089),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18085 ));
    InMux I__6588 (
            .O(N__41086),
            .I(N__41083));
    LocalMux I__6587 (
            .O(N__41083),
            .I(N__41080));
    Odrv4 I__6586 (
            .O(N__41080),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625 ));
    CascadeMux I__6585 (
            .O(N__41077),
            .I(N__41074));
    InMux I__6584 (
            .O(N__41074),
            .I(N__41071));
    LocalMux I__6583 (
            .O(N__41071),
            .I(N__41068));
    Odrv4 I__6582 (
            .O(N__41068),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640 ));
    InMux I__6581 (
            .O(N__41065),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18086 ));
    CascadeMux I__6580 (
            .O(N__41062),
            .I(N__41059));
    InMux I__6579 (
            .O(N__41059),
            .I(N__41056));
    LocalMux I__6578 (
            .O(N__41056),
            .I(N__41053));
    Odrv12 I__6577 (
            .O(N__41053),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624 ));
    InMux I__6576 (
            .O(N__41050),
            .I(N__41047));
    LocalMux I__6575 (
            .O(N__41047),
            .I(N__41044));
    Odrv4 I__6574 (
            .O(N__41044),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639 ));
    InMux I__6573 (
            .O(N__41041),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18087 ));
    InMux I__6572 (
            .O(N__41038),
            .I(N__41035));
    LocalMux I__6571 (
            .O(N__41035),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654 ));
    InMux I__6570 (
            .O(N__41032),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18073 ));
    CascadeMux I__6569 (
            .O(N__41029),
            .I(N__41026));
    InMux I__6568 (
            .O(N__41026),
            .I(N__41023));
    LocalMux I__6567 (
            .O(N__41023),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653 ));
    InMux I__6566 (
            .O(N__41020),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18074 ));
    InMux I__6565 (
            .O(N__41017),
            .I(N__41014));
    LocalMux I__6564 (
            .O(N__41014),
            .I(N__41011));
    Span4Mux_v I__6563 (
            .O(N__41011),
            .I(N__41008));
    Odrv4 I__6562 (
            .O(N__41008),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651 ));
    InMux I__6561 (
            .O(N__41005),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18075 ));
    InMux I__6560 (
            .O(N__41002),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652 ));
    CascadeMux I__6559 (
            .O(N__40999),
            .I(N__40996));
    InMux I__6558 (
            .O(N__40996),
            .I(N__40993));
    LocalMux I__6557 (
            .O(N__40993),
            .I(N__40990));
    Span4Mux_h I__6556 (
            .O(N__40990),
            .I(N__40987));
    Odrv4 I__6555 (
            .O(N__40987),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO ));
    CascadeMux I__6554 (
            .O(N__40984),
            .I(N__40981));
    InMux I__6553 (
            .O(N__40981),
            .I(N__40978));
    LocalMux I__6552 (
            .O(N__40978),
            .I(N__40975));
    Odrv12 I__6551 (
            .O(N__40975),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650 ));
    CascadeMux I__6550 (
            .O(N__40972),
            .I(N__40969));
    InMux I__6549 (
            .O(N__40969),
            .I(N__40966));
    LocalMux I__6548 (
            .O(N__40966),
            .I(N__40963));
    Odrv12 I__6547 (
            .O(N__40963),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634 ));
    InMux I__6546 (
            .O(N__40960),
            .I(N__40957));
    LocalMux I__6545 (
            .O(N__40957),
            .I(N__40954));
    Odrv4 I__6544 (
            .O(N__40954),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649 ));
    InMux I__6543 (
            .O(N__40951),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18077 ));
    InMux I__6542 (
            .O(N__40948),
            .I(N__40945));
    LocalMux I__6541 (
            .O(N__40945),
            .I(N__40942));
    Odrv12 I__6540 (
            .O(N__40942),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633 ));
    CascadeMux I__6539 (
            .O(N__40939),
            .I(N__40936));
    InMux I__6538 (
            .O(N__40936),
            .I(N__40933));
    LocalMux I__6537 (
            .O(N__40933),
            .I(N__40930));
    Odrv12 I__6536 (
            .O(N__40930),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648 ));
    InMux I__6535 (
            .O(N__40927),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18078 ));
    CascadeMux I__6534 (
            .O(N__40924),
            .I(N__40921));
    InMux I__6533 (
            .O(N__40921),
            .I(N__40918));
    LocalMux I__6532 (
            .O(N__40918),
            .I(N__40915));
    Odrv12 I__6531 (
            .O(N__40915),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632 ));
    InMux I__6530 (
            .O(N__40912),
            .I(N__40909));
    LocalMux I__6529 (
            .O(N__40909),
            .I(N__40906));
    Odrv4 I__6528 (
            .O(N__40906),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647 ));
    InMux I__6527 (
            .O(N__40903),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18079 ));
    InMux I__6526 (
            .O(N__40900),
            .I(N__40897));
    LocalMux I__6525 (
            .O(N__40897),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662 ));
    InMux I__6524 (
            .O(N__40894),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18065 ));
    InMux I__6523 (
            .O(N__40891),
            .I(N__40888));
    LocalMux I__6522 (
            .O(N__40888),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661 ));
    InMux I__6521 (
            .O(N__40885),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18066 ));
    InMux I__6520 (
            .O(N__40882),
            .I(N__40879));
    LocalMux I__6519 (
            .O(N__40879),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660 ));
    InMux I__6518 (
            .O(N__40876),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18067 ));
    InMux I__6517 (
            .O(N__40873),
            .I(N__40870));
    LocalMux I__6516 (
            .O(N__40870),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659 ));
    InMux I__6515 (
            .O(N__40867),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18068 ));
    InMux I__6514 (
            .O(N__40864),
            .I(N__40861));
    LocalMux I__6513 (
            .O(N__40861),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658 ));
    InMux I__6512 (
            .O(N__40858),
            .I(bfn_15_24_0_));
    InMux I__6511 (
            .O(N__40855),
            .I(N__40852));
    LocalMux I__6510 (
            .O(N__40852),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657 ));
    InMux I__6509 (
            .O(N__40849),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18070 ));
    InMux I__6508 (
            .O(N__40846),
            .I(N__40843));
    LocalMux I__6507 (
            .O(N__40843),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656 ));
    InMux I__6506 (
            .O(N__40840),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18071 ));
    InMux I__6505 (
            .O(N__40837),
            .I(N__40834));
    LocalMux I__6504 (
            .O(N__40834),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655 ));
    InMux I__6503 (
            .O(N__40831),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18072 ));
    InMux I__6502 (
            .O(N__40828),
            .I(N__40825));
    LocalMux I__6501 (
            .O(N__40825),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729 ));
    CascadeMux I__6500 (
            .O(N__40822),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_ ));
    CascadeMux I__6499 (
            .O(N__40819),
            .I(N__40816));
    InMux I__6498 (
            .O(N__40816),
            .I(N__40813));
    LocalMux I__6497 (
            .O(N__40813),
            .I(N__40810));
    Span4Mux_v I__6496 (
            .O(N__40810),
            .I(N__40807));
    Odrv4 I__6495 (
            .O(N__40807),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732 ));
    InMux I__6494 (
            .O(N__40804),
            .I(N__40795));
    InMux I__6493 (
            .O(N__40803),
            .I(N__40795));
    InMux I__6492 (
            .O(N__40802),
            .I(N__40795));
    LocalMux I__6491 (
            .O(N__40795),
            .I(N__40792));
    Odrv4 I__6490 (
            .O(N__40792),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759 ));
    CascadeMux I__6489 (
            .O(N__40789),
            .I(N__40786));
    InMux I__6488 (
            .O(N__40786),
            .I(N__40783));
    LocalMux I__6487 (
            .O(N__40783),
            .I(N__40780));
    Span4Mux_v I__6486 (
            .O(N__40780),
            .I(N__40777));
    Odrv4 I__6485 (
            .O(N__40777),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733 ));
    InMux I__6484 (
            .O(N__40774),
            .I(N__40771));
    LocalMux I__6483 (
            .O(N__40771),
            .I(N__40768));
    Span4Mux_h I__6482 (
            .O(N__40768),
            .I(N__40765));
    Odrv4 I__6481 (
            .O(N__40765),
            .I(n794_adj_2425));
    InMux I__6480 (
            .O(N__40762),
            .I(N__40759));
    LocalMux I__6479 (
            .O(N__40759),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666 ));
    InMux I__6478 (
            .O(N__40756),
            .I(N__40753));
    LocalMux I__6477 (
            .O(N__40753),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665 ));
    InMux I__6476 (
            .O(N__40750),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18062 ));
    InMux I__6475 (
            .O(N__40747),
            .I(N__40744));
    LocalMux I__6474 (
            .O(N__40744),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664 ));
    InMux I__6473 (
            .O(N__40741),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18063 ));
    InMux I__6472 (
            .O(N__40738),
            .I(N__40735));
    LocalMux I__6471 (
            .O(N__40735),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663 ));
    InMux I__6470 (
            .O(N__40732),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18064 ));
    InMux I__6469 (
            .O(N__40729),
            .I(N__40726));
    LocalMux I__6468 (
            .O(N__40726),
            .I(\foc.qCurrent_25 ));
    InMux I__6467 (
            .O(N__40723),
            .I(N__40720));
    LocalMux I__6466 (
            .O(N__40720),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730 ));
    InMux I__6465 (
            .O(N__40717),
            .I(N__40714));
    LocalMux I__6464 (
            .O(N__40714),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728 ));
    InMux I__6463 (
            .O(N__40711),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17973 ));
    CascadeMux I__6462 (
            .O(N__40708),
            .I(N__40705));
    InMux I__6461 (
            .O(N__40705),
            .I(N__40702));
    LocalMux I__6460 (
            .O(N__40702),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726 ));
    InMux I__6459 (
            .O(N__40699),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17974 ));
    InMux I__6458 (
            .O(N__40696),
            .I(N__40693));
    LocalMux I__6457 (
            .O(N__40693),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724 ));
    InMux I__6456 (
            .O(N__40690),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17975 ));
    CascadeMux I__6455 (
            .O(N__40687),
            .I(N__40684));
    InMux I__6454 (
            .O(N__40684),
            .I(N__40681));
    LocalMux I__6453 (
            .O(N__40681),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723 ));
    InMux I__6452 (
            .O(N__40678),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17976 ));
    CascadeMux I__6451 (
            .O(N__40675),
            .I(N__40671));
    CascadeMux I__6450 (
            .O(N__40674),
            .I(N__40667));
    InMux I__6449 (
            .O(N__40671),
            .I(N__40664));
    InMux I__6448 (
            .O(N__40670),
            .I(N__40659));
    InMux I__6447 (
            .O(N__40667),
            .I(N__40659));
    LocalMux I__6446 (
            .O(N__40664),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722 ));
    LocalMux I__6445 (
            .O(N__40659),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722 ));
    InMux I__6444 (
            .O(N__40654),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17977 ));
    InMux I__6443 (
            .O(N__40651),
            .I(N__40648));
    LocalMux I__6442 (
            .O(N__40648),
            .I(N__40645));
    Span4Mux_h I__6441 (
            .O(N__40645),
            .I(N__40642));
    Odrv4 I__6440 (
            .O(N__40642),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719 ));
    InMux I__6439 (
            .O(N__40639),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17978 ));
    InMux I__6438 (
            .O(N__40636),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721 ));
    InMux I__6437 (
            .O(N__40633),
            .I(N__40630));
    LocalMux I__6436 (
            .O(N__40630),
            .I(N__40627));
    Span4Mux_h I__6435 (
            .O(N__40627),
            .I(N__40624));
    Odrv4 I__6434 (
            .O(N__40624),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO ));
    InMux I__6433 (
            .O(N__40621),
            .I(N__40618));
    LocalMux I__6432 (
            .O(N__40618),
            .I(\foc.qCurrent_26 ));
    InMux I__6431 (
            .O(N__40615),
            .I(N__40612));
    LocalMux I__6430 (
            .O(N__40612),
            .I(\foc.qCurrent_12 ));
    InMux I__6429 (
            .O(N__40609),
            .I(N__40606));
    LocalMux I__6428 (
            .O(N__40606),
            .I(\foc.qCurrent_28 ));
    InMux I__6427 (
            .O(N__40603),
            .I(N__40600));
    LocalMux I__6426 (
            .O(N__40600),
            .I(\foc.qCurrent_20 ));
    CascadeMux I__6425 (
            .O(N__40597),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_ ));
    InMux I__6424 (
            .O(N__40594),
            .I(N__40591));
    LocalMux I__6423 (
            .O(N__40591),
            .I(N__40588));
    Odrv4 I__6422 (
            .O(N__40588),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758 ));
    CascadeMux I__6421 (
            .O(N__40585),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_ ));
    InMux I__6420 (
            .O(N__40582),
            .I(N__40579));
    LocalMux I__6419 (
            .O(N__40579),
            .I(\foc.qCurrent_31 ));
    InMux I__6418 (
            .O(N__40576),
            .I(N__40573));
    LocalMux I__6417 (
            .O(N__40573),
            .I(\foc.qCurrent_16 ));
    InMux I__6416 (
            .O(N__40570),
            .I(N__40567));
    LocalMux I__6415 (
            .O(N__40567),
            .I(\foc.qCurrent_14 ));
    InMux I__6414 (
            .O(N__40564),
            .I(N__40561));
    LocalMux I__6413 (
            .O(N__40561),
            .I(\foc.qCurrent_4 ));
    InMux I__6412 (
            .O(N__40558),
            .I(N__40555));
    LocalMux I__6411 (
            .O(N__40555),
            .I(\foc.qCurrent_11 ));
    InMux I__6410 (
            .O(N__40552),
            .I(N__40549));
    LocalMux I__6409 (
            .O(N__40549),
            .I(\foc.qCurrent_15 ));
    InMux I__6408 (
            .O(N__40546),
            .I(N__40543));
    LocalMux I__6407 (
            .O(N__40543),
            .I(\foc.qCurrent_22 ));
    InMux I__6406 (
            .O(N__40540),
            .I(N__40537));
    LocalMux I__6405 (
            .O(N__40537),
            .I(\foc.qCurrent_17 ));
    InMux I__6404 (
            .O(N__40534),
            .I(N__40531));
    LocalMux I__6403 (
            .O(N__40531),
            .I(\foc.qCurrent_24 ));
    InMux I__6402 (
            .O(N__40528),
            .I(N__40525));
    LocalMux I__6401 (
            .O(N__40525),
            .I(\foc.qCurrent_27 ));
    InMux I__6400 (
            .O(N__40522),
            .I(N__40519));
    LocalMux I__6399 (
            .O(N__40519),
            .I(\foc.qCurrent_6 ));
    InMux I__6398 (
            .O(N__40516),
            .I(N__40513));
    LocalMux I__6397 (
            .O(N__40513),
            .I(N__40509));
    InMux I__6396 (
            .O(N__40512),
            .I(N__40506));
    Odrv12 I__6395 (
            .O(N__40509),
            .I(\foc.u_Park_Transform.n741 ));
    LocalMux I__6394 (
            .O(N__40506),
            .I(\foc.u_Park_Transform.n741 ));
    InMux I__6393 (
            .O(N__40501),
            .I(N__40498));
    LocalMux I__6392 (
            .O(N__40498),
            .I(N__40494));
    InMux I__6391 (
            .O(N__40497),
            .I(N__40491));
    Span4Mux_v I__6390 (
            .O(N__40494),
            .I(N__40486));
    LocalMux I__6389 (
            .O(N__40491),
            .I(N__40486));
    Span4Mux_h I__6388 (
            .O(N__40486),
            .I(N__40481));
    InMux I__6387 (
            .O(N__40485),
            .I(N__40476));
    InMux I__6386 (
            .O(N__40484),
            .I(N__40476));
    Span4Mux_v I__6385 (
            .O(N__40481),
            .I(N__40470));
    LocalMux I__6384 (
            .O(N__40476),
            .I(N__40470));
    InMux I__6383 (
            .O(N__40475),
            .I(N__40467));
    Odrv4 I__6382 (
            .O(N__40470),
            .I(Look_Up_Table_out1_1_14));
    LocalMux I__6381 (
            .O(N__40467),
            .I(Look_Up_Table_out1_1_14));
    InMux I__6380 (
            .O(N__40462),
            .I(N__40459));
    LocalMux I__6379 (
            .O(N__40459),
            .I(N__40454));
    InMux I__6378 (
            .O(N__40458),
            .I(N__40451));
    InMux I__6377 (
            .O(N__40457),
            .I(N__40448));
    Span4Mux_v I__6376 (
            .O(N__40454),
            .I(N__40443));
    LocalMux I__6375 (
            .O(N__40451),
            .I(N__40440));
    LocalMux I__6374 (
            .O(N__40448),
            .I(N__40437));
    InMux I__6373 (
            .O(N__40447),
            .I(N__40434));
    InMux I__6372 (
            .O(N__40446),
            .I(N__40431));
    Span4Mux_v I__6371 (
            .O(N__40443),
            .I(N__40426));
    Span4Mux_v I__6370 (
            .O(N__40440),
            .I(N__40426));
    Span4Mux_h I__6369 (
            .O(N__40437),
            .I(N__40421));
    LocalMux I__6368 (
            .O(N__40434),
            .I(N__40421));
    LocalMux I__6367 (
            .O(N__40431),
            .I(N__40418));
    Odrv4 I__6366 (
            .O(N__40426),
            .I(Look_Up_Table_out1_1_15));
    Odrv4 I__6365 (
            .O(N__40421),
            .I(Look_Up_Table_out1_1_15));
    Odrv12 I__6364 (
            .O(N__40418),
            .I(Look_Up_Table_out1_1_15));
    InMux I__6363 (
            .O(N__40411),
            .I(N__40408));
    LocalMux I__6362 (
            .O(N__40408),
            .I(\foc.qCurrent_8 ));
    InMux I__6361 (
            .O(N__40405),
            .I(N__40399));
    InMux I__6360 (
            .O(N__40404),
            .I(N__40399));
    LocalMux I__6359 (
            .O(N__40399),
            .I(N__40396));
    Span4Mux_v I__6358 (
            .O(N__40396),
            .I(N__40393));
    Odrv4 I__6357 (
            .O(N__40393),
            .I(\foc.Look_Up_Table_out1_1_1 ));
    InMux I__6356 (
            .O(N__40390),
            .I(N__40380));
    CascadeMux I__6355 (
            .O(N__40389),
            .I(N__40377));
    CascadeMux I__6354 (
            .O(N__40388),
            .I(N__40373));
    CascadeMux I__6353 (
            .O(N__40387),
            .I(N__40369));
    CascadeMux I__6352 (
            .O(N__40386),
            .I(N__40364));
    CascadeMux I__6351 (
            .O(N__40385),
            .I(N__40361));
    CascadeMux I__6350 (
            .O(N__40384),
            .I(N__40357));
    CascadeMux I__6349 (
            .O(N__40383),
            .I(N__40353));
    LocalMux I__6348 (
            .O(N__40380),
            .I(N__40345));
    InMux I__6347 (
            .O(N__40377),
            .I(N__40332));
    InMux I__6346 (
            .O(N__40376),
            .I(N__40332));
    InMux I__6345 (
            .O(N__40373),
            .I(N__40332));
    InMux I__6344 (
            .O(N__40372),
            .I(N__40332));
    InMux I__6343 (
            .O(N__40369),
            .I(N__40332));
    InMux I__6342 (
            .O(N__40368),
            .I(N__40332));
    InMux I__6341 (
            .O(N__40367),
            .I(N__40327));
    InMux I__6340 (
            .O(N__40364),
            .I(N__40327));
    InMux I__6339 (
            .O(N__40361),
            .I(N__40314));
    InMux I__6338 (
            .O(N__40360),
            .I(N__40314));
    InMux I__6337 (
            .O(N__40357),
            .I(N__40314));
    InMux I__6336 (
            .O(N__40356),
            .I(N__40314));
    InMux I__6335 (
            .O(N__40353),
            .I(N__40314));
    InMux I__6334 (
            .O(N__40352),
            .I(N__40314));
    CascadeMux I__6333 (
            .O(N__40351),
            .I(N__40308));
    CascadeMux I__6332 (
            .O(N__40350),
            .I(N__40304));
    InMux I__6331 (
            .O(N__40349),
            .I(N__40296));
    InMux I__6330 (
            .O(N__40348),
            .I(N__40296));
    Span4Mux_v I__6329 (
            .O(N__40345),
            .I(N__40287));
    LocalMux I__6328 (
            .O(N__40332),
            .I(N__40287));
    LocalMux I__6327 (
            .O(N__40327),
            .I(N__40287));
    LocalMux I__6326 (
            .O(N__40314),
            .I(N__40287));
    InMux I__6325 (
            .O(N__40313),
            .I(N__40284));
    InMux I__6324 (
            .O(N__40312),
            .I(N__40271));
    InMux I__6323 (
            .O(N__40311),
            .I(N__40271));
    InMux I__6322 (
            .O(N__40308),
            .I(N__40271));
    InMux I__6321 (
            .O(N__40307),
            .I(N__40271));
    InMux I__6320 (
            .O(N__40304),
            .I(N__40271));
    InMux I__6319 (
            .O(N__40303),
            .I(N__40271));
    CascadeMux I__6318 (
            .O(N__40302),
            .I(N__40266));
    CascadeMux I__6317 (
            .O(N__40301),
            .I(N__40262));
    LocalMux I__6316 (
            .O(N__40296),
            .I(N__40258));
    Span4Mux_v I__6315 (
            .O(N__40287),
            .I(N__40251));
    LocalMux I__6314 (
            .O(N__40284),
            .I(N__40251));
    LocalMux I__6313 (
            .O(N__40271),
            .I(N__40251));
    InMux I__6312 (
            .O(N__40270),
            .I(N__40248));
    InMux I__6311 (
            .O(N__40269),
            .I(N__40237));
    InMux I__6310 (
            .O(N__40266),
            .I(N__40237));
    InMux I__6309 (
            .O(N__40265),
            .I(N__40237));
    InMux I__6308 (
            .O(N__40262),
            .I(N__40237));
    InMux I__6307 (
            .O(N__40261),
            .I(N__40237));
    Odrv4 I__6306 (
            .O(N__40258),
            .I(\foc.u_Park_Transform.n592 ));
    Odrv4 I__6305 (
            .O(N__40251),
            .I(\foc.u_Park_Transform.n592 ));
    LocalMux I__6304 (
            .O(N__40248),
            .I(\foc.u_Park_Transform.n592 ));
    LocalMux I__6303 (
            .O(N__40237),
            .I(\foc.u_Park_Transform.n592 ));
    InMux I__6302 (
            .O(N__40228),
            .I(N__40225));
    LocalMux I__6301 (
            .O(N__40225),
            .I(N__40222));
    Odrv4 I__6300 (
            .O(N__40222),
            .I(\foc.qCurrent_3 ));
    InMux I__6299 (
            .O(N__40219),
            .I(N__40216));
    LocalMux I__6298 (
            .O(N__40216),
            .I(\foc.qCurrent_18 ));
    InMux I__6297 (
            .O(N__40213),
            .I(N__40210));
    LocalMux I__6296 (
            .O(N__40210),
            .I(\foc.qCurrent_19 ));
    InMux I__6295 (
            .O(N__40207),
            .I(N__40204));
    LocalMux I__6294 (
            .O(N__40204),
            .I(\foc.qCurrent_13 ));
    InMux I__6293 (
            .O(N__40201),
            .I(\foc.u_Park_Transform.n17059 ));
    InMux I__6292 (
            .O(N__40198),
            .I(N__40195));
    LocalMux I__6291 (
            .O(N__40195),
            .I(\foc.u_Park_Transform.n446 ));
    InMux I__6290 (
            .O(N__40192),
            .I(bfn_15_16_0_));
    InMux I__6289 (
            .O(N__40189),
            .I(N__40186));
    LocalMux I__6288 (
            .O(N__40186),
            .I(\foc.u_Park_Transform.n495 ));
    InMux I__6287 (
            .O(N__40183),
            .I(\foc.u_Park_Transform.n17061 ));
    InMux I__6286 (
            .O(N__40180),
            .I(N__40177));
    LocalMux I__6285 (
            .O(N__40177),
            .I(\foc.u_Park_Transform.n544 ));
    InMux I__6284 (
            .O(N__40174),
            .I(\foc.u_Park_Transform.n17062 ));
    InMux I__6283 (
            .O(N__40171),
            .I(N__40168));
    LocalMux I__6282 (
            .O(N__40168),
            .I(\foc.u_Park_Transform.n593 ));
    InMux I__6281 (
            .O(N__40165),
            .I(\foc.u_Park_Transform.n17063 ));
    InMux I__6280 (
            .O(N__40162),
            .I(N__40159));
    LocalMux I__6279 (
            .O(N__40159),
            .I(\foc.u_Park_Transform.n642 ));
    InMux I__6278 (
            .O(N__40156),
            .I(\foc.u_Park_Transform.n17064 ));
    CascadeMux I__6277 (
            .O(N__40153),
            .I(N__40150));
    InMux I__6276 (
            .O(N__40150),
            .I(N__40147));
    LocalMux I__6275 (
            .O(N__40147),
            .I(\foc.u_Park_Transform.n691 ));
    InMux I__6274 (
            .O(N__40144),
            .I(\foc.u_Park_Transform.n17065 ));
    InMux I__6273 (
            .O(N__40141),
            .I(N__40138));
    LocalMux I__6272 (
            .O(N__40138),
            .I(N__40135));
    Span4Mux_v I__6271 (
            .O(N__40135),
            .I(N__40132));
    Odrv4 I__6270 (
            .O(N__40132),
            .I(\foc.u_Park_Transform.n742_adj_2086 ));
    InMux I__6269 (
            .O(N__40129),
            .I(\foc.u_Park_Transform.n17066 ));
    InMux I__6268 (
            .O(N__40126),
            .I(\foc.u_Park_Transform.n743_adj_2096 ));
    CascadeMux I__6267 (
            .O(N__40123),
            .I(N__40120));
    InMux I__6266 (
            .O(N__40120),
            .I(N__40117));
    LocalMux I__6265 (
            .O(N__40117),
            .I(N__40114));
    Span4Mux_v I__6264 (
            .O(N__40114),
            .I(N__40111));
    Odrv4 I__6263 (
            .O(N__40111),
            .I(\foc.u_Park_Transform.n743_adj_2096_THRU_CO ));
    InMux I__6262 (
            .O(N__40108),
            .I(\foc.u_Park_Transform.n751 ));
    CascadeMux I__6261 (
            .O(N__40105),
            .I(N__40102));
    InMux I__6260 (
            .O(N__40102),
            .I(N__40099));
    LocalMux I__6259 (
            .O(N__40099),
            .I(N__40096));
    Span4Mux_v I__6258 (
            .O(N__40096),
            .I(N__40093));
    Odrv4 I__6257 (
            .O(N__40093),
            .I(\foc.u_Park_Transform.n751_THRU_CO ));
    CascadeMux I__6256 (
            .O(N__40090),
            .I(N__40087));
    InMux I__6255 (
            .O(N__40087),
            .I(N__40084));
    LocalMux I__6254 (
            .O(N__40084),
            .I(\foc.u_Park_Transform.n54 ));
    InMux I__6253 (
            .O(N__40081),
            .I(N__40078));
    LocalMux I__6252 (
            .O(N__40078),
            .I(\foc.u_Park_Transform.n103 ));
    InMux I__6251 (
            .O(N__40075),
            .I(\foc.u_Park_Transform.n17053 ));
    CascadeMux I__6250 (
            .O(N__40072),
            .I(N__40069));
    InMux I__6249 (
            .O(N__40069),
            .I(N__40066));
    LocalMux I__6248 (
            .O(N__40066),
            .I(\foc.u_Park_Transform.n152 ));
    InMux I__6247 (
            .O(N__40063),
            .I(\foc.u_Park_Transform.n17054 ));
    InMux I__6246 (
            .O(N__40060),
            .I(N__40057));
    LocalMux I__6245 (
            .O(N__40057),
            .I(\foc.u_Park_Transform.n201 ));
    InMux I__6244 (
            .O(N__40054),
            .I(\foc.u_Park_Transform.n17055 ));
    CascadeMux I__6243 (
            .O(N__40051),
            .I(N__40048));
    InMux I__6242 (
            .O(N__40048),
            .I(N__40045));
    LocalMux I__6241 (
            .O(N__40045),
            .I(\foc.u_Park_Transform.n250 ));
    InMux I__6240 (
            .O(N__40042),
            .I(\foc.u_Park_Transform.n17056 ));
    InMux I__6239 (
            .O(N__40039),
            .I(N__40036));
    LocalMux I__6238 (
            .O(N__40036),
            .I(\foc.u_Park_Transform.n299 ));
    InMux I__6237 (
            .O(N__40033),
            .I(\foc.u_Park_Transform.n17057 ));
    CascadeMux I__6236 (
            .O(N__40030),
            .I(N__40027));
    InMux I__6235 (
            .O(N__40027),
            .I(N__40024));
    LocalMux I__6234 (
            .O(N__40024),
            .I(\foc.u_Park_Transform.n348 ));
    InMux I__6233 (
            .O(N__40021),
            .I(\foc.u_Park_Transform.n17058 ));
    InMux I__6232 (
            .O(N__40018),
            .I(N__40015));
    LocalMux I__6231 (
            .O(N__40015),
            .I(\foc.u_Park_Transform.n397 ));
    InMux I__6230 (
            .O(N__40012),
            .I(N__40009));
    LocalMux I__6229 (
            .O(N__40009),
            .I(\foc.u_Park_Transform.n357 ));
    InMux I__6228 (
            .O(N__40006),
            .I(\foc.u_Park_Transform.n17029 ));
    CascadeMux I__6227 (
            .O(N__40003),
            .I(N__40000));
    InMux I__6226 (
            .O(N__40000),
            .I(N__39997));
    LocalMux I__6225 (
            .O(N__39997),
            .I(\foc.u_Park_Transform.n406 ));
    InMux I__6224 (
            .O(N__39994),
            .I(bfn_15_14_0_));
    InMux I__6223 (
            .O(N__39991),
            .I(N__39988));
    LocalMux I__6222 (
            .O(N__39988),
            .I(\foc.u_Park_Transform.n455 ));
    InMux I__6221 (
            .O(N__39985),
            .I(\foc.u_Park_Transform.n17031 ));
    CascadeMux I__6220 (
            .O(N__39982),
            .I(N__39979));
    InMux I__6219 (
            .O(N__39979),
            .I(N__39976));
    LocalMux I__6218 (
            .O(N__39976),
            .I(\foc.u_Park_Transform.n504 ));
    InMux I__6217 (
            .O(N__39973),
            .I(\foc.u_Park_Transform.n17032 ));
    InMux I__6216 (
            .O(N__39970),
            .I(N__39967));
    LocalMux I__6215 (
            .O(N__39967),
            .I(\foc.u_Park_Transform.n553 ));
    InMux I__6214 (
            .O(N__39964),
            .I(\foc.u_Park_Transform.n17033 ));
    CascadeMux I__6213 (
            .O(N__39961),
            .I(N__39958));
    InMux I__6212 (
            .O(N__39958),
            .I(N__39955));
    LocalMux I__6211 (
            .O(N__39955),
            .I(\foc.u_Park_Transform.n602 ));
    InMux I__6210 (
            .O(N__39952),
            .I(\foc.u_Park_Transform.n17034 ));
    InMux I__6209 (
            .O(N__39949),
            .I(N__39946));
    LocalMux I__6208 (
            .O(N__39946),
            .I(\foc.u_Park_Transform.n651 ));
    InMux I__6207 (
            .O(N__39943),
            .I(\foc.u_Park_Transform.n17035 ));
    CascadeMux I__6206 (
            .O(N__39940),
            .I(N__39937));
    InMux I__6205 (
            .O(N__39937),
            .I(N__39934));
    LocalMux I__6204 (
            .O(N__39934),
            .I(\foc.u_Park_Transform.n700 ));
    InMux I__6203 (
            .O(N__39931),
            .I(N__39928));
    LocalMux I__6202 (
            .O(N__39928),
            .I(N__39925));
    Span4Mux_h I__6201 (
            .O(N__39925),
            .I(N__39922));
    Odrv4 I__6200 (
            .O(N__39922),
            .I(\foc.u_Park_Transform.n750_adj_2117 ));
    InMux I__6199 (
            .O(N__39919),
            .I(\foc.u_Park_Transform.n17036 ));
    CascadeMux I__6198 (
            .O(N__39916),
            .I(N__39913));
    InMux I__6197 (
            .O(N__39913),
            .I(N__39910));
    LocalMux I__6196 (
            .O(N__39910),
            .I(\foc.u_Park_Transform.n694_adj_2097 ));
    InMux I__6195 (
            .O(N__39907),
            .I(N__39904));
    LocalMux I__6194 (
            .O(N__39904),
            .I(N__39901));
    Span4Mux_h I__6193 (
            .O(N__39901),
            .I(N__39898));
    Odrv4 I__6192 (
            .O(N__39898),
            .I(\foc.u_Park_Transform.n742 ));
    InMux I__6191 (
            .O(N__39895),
            .I(\foc.u_Park_Transform.n17249 ));
    InMux I__6190 (
            .O(N__39892),
            .I(\foc.u_Park_Transform.n743 ));
    CascadeMux I__6189 (
            .O(N__39889),
            .I(N__39886));
    InMux I__6188 (
            .O(N__39886),
            .I(N__39883));
    LocalMux I__6187 (
            .O(N__39883),
            .I(N__39880));
    Span4Mux_v I__6186 (
            .O(N__39880),
            .I(N__39877));
    Odrv4 I__6185 (
            .O(N__39877),
            .I(\foc.u_Park_Transform.n743_THRU_CO ));
    InMux I__6184 (
            .O(N__39874),
            .I(N__39871));
    LocalMux I__6183 (
            .O(N__39871),
            .I(\foc.u_Park_Transform.n63 ));
    InMux I__6182 (
            .O(N__39868),
            .I(\foc.u_Park_Transform.n17023 ));
    CascadeMux I__6181 (
            .O(N__39865),
            .I(N__39862));
    InMux I__6180 (
            .O(N__39862),
            .I(N__39859));
    LocalMux I__6179 (
            .O(N__39859),
            .I(\foc.u_Park_Transform.n112 ));
    InMux I__6178 (
            .O(N__39856),
            .I(\foc.u_Park_Transform.n17024 ));
    InMux I__6177 (
            .O(N__39853),
            .I(N__39850));
    LocalMux I__6176 (
            .O(N__39850),
            .I(\foc.u_Park_Transform.n161 ));
    InMux I__6175 (
            .O(N__39847),
            .I(\foc.u_Park_Transform.n17025 ));
    CascadeMux I__6174 (
            .O(N__39844),
            .I(N__39841));
    InMux I__6173 (
            .O(N__39841),
            .I(N__39838));
    LocalMux I__6172 (
            .O(N__39838),
            .I(\foc.u_Park_Transform.n210 ));
    InMux I__6171 (
            .O(N__39835),
            .I(\foc.u_Park_Transform.n17026 ));
    InMux I__6170 (
            .O(N__39832),
            .I(N__39829));
    LocalMux I__6169 (
            .O(N__39829),
            .I(\foc.u_Park_Transform.n259 ));
    InMux I__6168 (
            .O(N__39826),
            .I(\foc.u_Park_Transform.n17027 ));
    CascadeMux I__6167 (
            .O(N__39823),
            .I(N__39820));
    InMux I__6166 (
            .O(N__39820),
            .I(N__39817));
    LocalMux I__6165 (
            .O(N__39817),
            .I(N__39814));
    Odrv4 I__6164 (
            .O(N__39814),
            .I(\foc.u_Park_Transform.n308 ));
    InMux I__6163 (
            .O(N__39811),
            .I(\foc.u_Park_Transform.n17028 ));
    CascadeMux I__6162 (
            .O(N__39808),
            .I(N__39805));
    InMux I__6161 (
            .O(N__39805),
            .I(N__39802));
    LocalMux I__6160 (
            .O(N__39802),
            .I(N__39799));
    Odrv4 I__6159 (
            .O(N__39799),
            .I(\foc.u_Park_Transform.n348_adj_2082 ));
    InMux I__6158 (
            .O(N__39796),
            .I(\foc.u_Park_Transform.n17241 ));
    InMux I__6157 (
            .O(N__39793),
            .I(N__39790));
    LocalMux I__6156 (
            .O(N__39790),
            .I(\foc.u_Park_Transform.n351_adj_2108 ));
    InMux I__6155 (
            .O(N__39787),
            .I(N__39784));
    LocalMux I__6154 (
            .O(N__39784),
            .I(\foc.u_Park_Transform.n397_adj_2081 ));
    InMux I__6153 (
            .O(N__39781),
            .I(\foc.u_Park_Transform.n17242 ));
    CascadeMux I__6152 (
            .O(N__39778),
            .I(N__39775));
    InMux I__6151 (
            .O(N__39775),
            .I(N__39772));
    LocalMux I__6150 (
            .O(N__39772),
            .I(\foc.u_Park_Transform.n400_adj_2106 ));
    CascadeMux I__6149 (
            .O(N__39769),
            .I(N__39766));
    InMux I__6148 (
            .O(N__39766),
            .I(N__39763));
    LocalMux I__6147 (
            .O(N__39763),
            .I(N__39760));
    Odrv4 I__6146 (
            .O(N__39760),
            .I(\foc.u_Park_Transform.n446_adj_2079 ));
    InMux I__6145 (
            .O(N__39757),
            .I(bfn_15_12_0_));
    InMux I__6144 (
            .O(N__39754),
            .I(N__39751));
    LocalMux I__6143 (
            .O(N__39751),
            .I(\foc.u_Park_Transform.n449_adj_2103 ));
    InMux I__6142 (
            .O(N__39748),
            .I(N__39745));
    LocalMux I__6141 (
            .O(N__39745),
            .I(N__39742));
    Odrv4 I__6140 (
            .O(N__39742),
            .I(\foc.u_Park_Transform.n495_adj_2077 ));
    InMux I__6139 (
            .O(N__39739),
            .I(\foc.u_Park_Transform.n17244 ));
    CascadeMux I__6138 (
            .O(N__39736),
            .I(N__39733));
    InMux I__6137 (
            .O(N__39733),
            .I(N__39730));
    LocalMux I__6136 (
            .O(N__39730),
            .I(\foc.u_Park_Transform.n498_adj_2102 ));
    CascadeMux I__6135 (
            .O(N__39727),
            .I(N__39724));
    InMux I__6134 (
            .O(N__39724),
            .I(N__39721));
    LocalMux I__6133 (
            .O(N__39721),
            .I(N__39718));
    Odrv4 I__6132 (
            .O(N__39718),
            .I(\foc.u_Park_Transform.n544_adj_2074 ));
    InMux I__6131 (
            .O(N__39715),
            .I(\foc.u_Park_Transform.n17245 ));
    InMux I__6130 (
            .O(N__39712),
            .I(N__39709));
    LocalMux I__6129 (
            .O(N__39709),
            .I(\foc.u_Park_Transform.n547_adj_2100 ));
    InMux I__6128 (
            .O(N__39706),
            .I(N__39703));
    LocalMux I__6127 (
            .O(N__39703),
            .I(N__39700));
    Odrv4 I__6126 (
            .O(N__39700),
            .I(\foc.u_Park_Transform.n593_adj_2073 ));
    InMux I__6125 (
            .O(N__39697),
            .I(\foc.u_Park_Transform.n17246 ));
    CascadeMux I__6124 (
            .O(N__39694),
            .I(N__39691));
    InMux I__6123 (
            .O(N__39691),
            .I(N__39688));
    LocalMux I__6122 (
            .O(N__39688),
            .I(\foc.u_Park_Transform.n596_adj_2099 ));
    CascadeMux I__6121 (
            .O(N__39685),
            .I(N__39682));
    InMux I__6120 (
            .O(N__39682),
            .I(N__39679));
    LocalMux I__6119 (
            .O(N__39679),
            .I(N__39676));
    Odrv4 I__6118 (
            .O(N__39676),
            .I(\foc.u_Park_Transform.n642_adj_2072 ));
    InMux I__6117 (
            .O(N__39673),
            .I(\foc.u_Park_Transform.n17247 ));
    InMux I__6116 (
            .O(N__39670),
            .I(N__39667));
    LocalMux I__6115 (
            .O(N__39667),
            .I(\foc.u_Park_Transform.n645_adj_2098 ));
    CascadeMux I__6114 (
            .O(N__39664),
            .I(N__39661));
    InMux I__6113 (
            .O(N__39661),
            .I(N__39658));
    LocalMux I__6112 (
            .O(N__39658),
            .I(N__39655));
    Odrv4 I__6111 (
            .O(N__39655),
            .I(\foc.u_Park_Transform.n691_adj_2071 ));
    InMux I__6110 (
            .O(N__39652),
            .I(\foc.u_Park_Transform.n17248 ));
    CascadeMux I__6109 (
            .O(N__39649),
            .I(N__39646));
    InMux I__6108 (
            .O(N__39646),
            .I(N__39642));
    InMux I__6107 (
            .O(N__39645),
            .I(N__39639));
    LocalMux I__6106 (
            .O(N__39642),
            .I(N__39634));
    LocalMux I__6105 (
            .O(N__39639),
            .I(N__39634));
    Span4Mux_v I__6104 (
            .O(N__39634),
            .I(N__39631));
    Odrv4 I__6103 (
            .O(N__39631),
            .I(\foc.u_Park_Transform.n738 ));
    InMux I__6102 (
            .O(N__39628),
            .I(\foc.u_Park_Transform.n17264 ));
    InMux I__6101 (
            .O(N__39625),
            .I(\foc.u_Park_Transform.n739 ));
    CascadeMux I__6100 (
            .O(N__39622),
            .I(N__39619));
    InMux I__6099 (
            .O(N__39619),
            .I(N__39616));
    LocalMux I__6098 (
            .O(N__39616),
            .I(N__39613));
    Span4Mux_h I__6097 (
            .O(N__39613),
            .I(N__39610));
    Odrv4 I__6096 (
            .O(N__39610),
            .I(\foc.u_Park_Transform.n739_THRU_CO ));
    InMux I__6095 (
            .O(N__39607),
            .I(N__39604));
    LocalMux I__6094 (
            .O(N__39604),
            .I(N__39601));
    Odrv4 I__6093 (
            .O(N__39601),
            .I(\foc.u_Park_Transform.n54_adj_2095 ));
    CascadeMux I__6092 (
            .O(N__39598),
            .I(N__39595));
    InMux I__6091 (
            .O(N__39595),
            .I(N__39592));
    LocalMux I__6090 (
            .O(N__39592),
            .I(\foc.u_Park_Transform.n57_adj_2116 ));
    InMux I__6089 (
            .O(N__39589),
            .I(N__39586));
    LocalMux I__6088 (
            .O(N__39586),
            .I(N__39583));
    Odrv4 I__6087 (
            .O(N__39583),
            .I(\foc.u_Park_Transform.n103_adj_2092 ));
    InMux I__6086 (
            .O(N__39580),
            .I(\foc.u_Park_Transform.n17236 ));
    CascadeMux I__6085 (
            .O(N__39577),
            .I(N__39574));
    InMux I__6084 (
            .O(N__39574),
            .I(N__39571));
    LocalMux I__6083 (
            .O(N__39571),
            .I(\foc.u_Park_Transform.n106_adj_2115 ));
    CascadeMux I__6082 (
            .O(N__39568),
            .I(N__39565));
    InMux I__6081 (
            .O(N__39565),
            .I(N__39562));
    LocalMux I__6080 (
            .O(N__39562),
            .I(N__39559));
    Odrv12 I__6079 (
            .O(N__39559),
            .I(\foc.u_Park_Transform.n152_adj_2088 ));
    InMux I__6078 (
            .O(N__39556),
            .I(\foc.u_Park_Transform.n17237 ));
    InMux I__6077 (
            .O(N__39553),
            .I(N__39550));
    LocalMux I__6076 (
            .O(N__39550),
            .I(\foc.u_Park_Transform.n155_adj_2114 ));
    InMux I__6075 (
            .O(N__39547),
            .I(N__39544));
    LocalMux I__6074 (
            .O(N__39544),
            .I(N__39541));
    Odrv12 I__6073 (
            .O(N__39541),
            .I(\foc.u_Park_Transform.n201_adj_2085 ));
    InMux I__6072 (
            .O(N__39538),
            .I(\foc.u_Park_Transform.n17238 ));
    CascadeMux I__6071 (
            .O(N__39535),
            .I(N__39532));
    InMux I__6070 (
            .O(N__39532),
            .I(N__39529));
    LocalMux I__6069 (
            .O(N__39529),
            .I(\foc.u_Park_Transform.n204_adj_2113 ));
    CascadeMux I__6068 (
            .O(N__39526),
            .I(N__39523));
    InMux I__6067 (
            .O(N__39523),
            .I(N__39520));
    LocalMux I__6066 (
            .O(N__39520),
            .I(N__39517));
    Odrv4 I__6065 (
            .O(N__39517),
            .I(\foc.u_Park_Transform.n250_adj_2084 ));
    InMux I__6064 (
            .O(N__39514),
            .I(\foc.u_Park_Transform.n17239 ));
    InMux I__6063 (
            .O(N__39511),
            .I(N__39508));
    LocalMux I__6062 (
            .O(N__39508),
            .I(\foc.u_Park_Transform.n253_adj_2112 ));
    InMux I__6061 (
            .O(N__39505),
            .I(N__39502));
    LocalMux I__6060 (
            .O(N__39502),
            .I(N__39499));
    Odrv4 I__6059 (
            .O(N__39499),
            .I(\foc.u_Park_Transform.n299_adj_2083 ));
    InMux I__6058 (
            .O(N__39496),
            .I(\foc.u_Park_Transform.n17240 ));
    CascadeMux I__6057 (
            .O(N__39493),
            .I(N__39490));
    InMux I__6056 (
            .O(N__39490),
            .I(N__39487));
    LocalMux I__6055 (
            .O(N__39487),
            .I(\foc.u_Park_Transform.n302_adj_2111 ));
    InMux I__6054 (
            .O(N__39484),
            .I(N__39481));
    LocalMux I__6053 (
            .O(N__39481),
            .I(N__39478));
    Odrv4 I__6052 (
            .O(N__39478),
            .I(\foc.u_Park_Transform.Product1_mul_temp_7 ));
    InMux I__6051 (
            .O(N__39475),
            .I(\foc.u_Park_Transform.n17256 ));
    InMux I__6050 (
            .O(N__39472),
            .I(N__39469));
    LocalMux I__6049 (
            .O(N__39469),
            .I(N__39466));
    Span4Mux_h I__6048 (
            .O(N__39466),
            .I(N__39463));
    Odrv4 I__6047 (
            .O(N__39463),
            .I(\foc.u_Park_Transform.Product1_mul_temp_8 ));
    InMux I__6046 (
            .O(N__39460),
            .I(\foc.u_Park_Transform.n17257 ));
    InMux I__6045 (
            .O(N__39457),
            .I(N__39454));
    LocalMux I__6044 (
            .O(N__39454),
            .I(N__39451));
    Sp12to4 I__6043 (
            .O(N__39451),
            .I(N__39448));
    Odrv12 I__6042 (
            .O(N__39448),
            .I(\foc.u_Park_Transform.Product1_mul_temp_9 ));
    InMux I__6041 (
            .O(N__39445),
            .I(bfn_15_10_0_));
    InMux I__6040 (
            .O(N__39442),
            .I(N__39439));
    LocalMux I__6039 (
            .O(N__39439),
            .I(N__39436));
    Span4Mux_h I__6038 (
            .O(N__39436),
            .I(N__39433));
    Odrv4 I__6037 (
            .O(N__39433),
            .I(\foc.u_Park_Transform.Product1_mul_temp_10 ));
    InMux I__6036 (
            .O(N__39430),
            .I(\foc.u_Park_Transform.n17259 ));
    InMux I__6035 (
            .O(N__39427),
            .I(N__39424));
    LocalMux I__6034 (
            .O(N__39424),
            .I(N__39421));
    Odrv4 I__6033 (
            .O(N__39421),
            .I(\foc.u_Park_Transform.Product1_mul_temp_11 ));
    InMux I__6032 (
            .O(N__39418),
            .I(\foc.u_Park_Transform.n17260 ));
    InMux I__6031 (
            .O(N__39415),
            .I(N__39412));
    LocalMux I__6030 (
            .O(N__39412),
            .I(N__39409));
    Odrv4 I__6029 (
            .O(N__39409),
            .I(\foc.u_Park_Transform.Product1_mul_temp_12 ));
    InMux I__6028 (
            .O(N__39406),
            .I(\foc.u_Park_Transform.n17261 ));
    InMux I__6027 (
            .O(N__39403),
            .I(N__39400));
    LocalMux I__6026 (
            .O(N__39400),
            .I(N__39397));
    Odrv4 I__6025 (
            .O(N__39397),
            .I(\foc.u_Park_Transform.Product1_mul_temp_13 ));
    InMux I__6024 (
            .O(N__39394),
            .I(\foc.u_Park_Transform.n17262 ));
    CascadeMux I__6023 (
            .O(N__39391),
            .I(N__39381));
    CascadeMux I__6022 (
            .O(N__39390),
            .I(N__39377));
    CascadeMux I__6021 (
            .O(N__39389),
            .I(N__39373));
    CascadeMux I__6020 (
            .O(N__39388),
            .I(N__39369));
    CascadeMux I__6019 (
            .O(N__39387),
            .I(N__39366));
    CascadeMux I__6018 (
            .O(N__39386),
            .I(N__39362));
    CascadeMux I__6017 (
            .O(N__39385),
            .I(N__39358));
    CascadeMux I__6016 (
            .O(N__39384),
            .I(N__39354));
    InMux I__6015 (
            .O(N__39381),
            .I(N__39345));
    InMux I__6014 (
            .O(N__39380),
            .I(N__39330));
    InMux I__6013 (
            .O(N__39377),
            .I(N__39330));
    InMux I__6012 (
            .O(N__39376),
            .I(N__39330));
    InMux I__6011 (
            .O(N__39373),
            .I(N__39330));
    InMux I__6010 (
            .O(N__39372),
            .I(N__39330));
    InMux I__6009 (
            .O(N__39369),
            .I(N__39330));
    InMux I__6008 (
            .O(N__39366),
            .I(N__39330));
    InMux I__6007 (
            .O(N__39365),
            .I(N__39317));
    InMux I__6006 (
            .O(N__39362),
            .I(N__39317));
    InMux I__6005 (
            .O(N__39361),
            .I(N__39317));
    InMux I__6004 (
            .O(N__39358),
            .I(N__39317));
    InMux I__6003 (
            .O(N__39357),
            .I(N__39317));
    InMux I__6002 (
            .O(N__39354),
            .I(N__39317));
    CascadeMux I__6001 (
            .O(N__39353),
            .I(N__39310));
    CascadeMux I__6000 (
            .O(N__39352),
            .I(N__39307));
    CascadeMux I__5999 (
            .O(N__39351),
            .I(N__39304));
    CascadeMux I__5998 (
            .O(N__39350),
            .I(N__39301));
    CascadeMux I__5997 (
            .O(N__39349),
            .I(N__39298));
    CascadeMux I__5996 (
            .O(N__39348),
            .I(N__39295));
    LocalMux I__5995 (
            .O(N__39345),
            .I(N__39292));
    LocalMux I__5994 (
            .O(N__39330),
            .I(N__39287));
    LocalMux I__5993 (
            .O(N__39317),
            .I(N__39287));
    CascadeMux I__5992 (
            .O(N__39316),
            .I(N__39283));
    CascadeMux I__5991 (
            .O(N__39315),
            .I(N__39279));
    CascadeMux I__5990 (
            .O(N__39314),
            .I(N__39275));
    CascadeMux I__5989 (
            .O(N__39313),
            .I(N__39271));
    InMux I__5988 (
            .O(N__39310),
            .I(N__39264));
    InMux I__5987 (
            .O(N__39307),
            .I(N__39264));
    InMux I__5986 (
            .O(N__39304),
            .I(N__39264));
    InMux I__5985 (
            .O(N__39301),
            .I(N__39257));
    InMux I__5984 (
            .O(N__39298),
            .I(N__39257));
    InMux I__5983 (
            .O(N__39295),
            .I(N__39257));
    Span4Mux_v I__5982 (
            .O(N__39292),
            .I(N__39252));
    Span4Mux_v I__5981 (
            .O(N__39287),
            .I(N__39252));
    InMux I__5980 (
            .O(N__39286),
            .I(N__39235));
    InMux I__5979 (
            .O(N__39283),
            .I(N__39235));
    InMux I__5978 (
            .O(N__39282),
            .I(N__39235));
    InMux I__5977 (
            .O(N__39279),
            .I(N__39235));
    InMux I__5976 (
            .O(N__39278),
            .I(N__39235));
    InMux I__5975 (
            .O(N__39275),
            .I(N__39235));
    InMux I__5974 (
            .O(N__39274),
            .I(N__39235));
    InMux I__5973 (
            .O(N__39271),
            .I(N__39235));
    LocalMux I__5972 (
            .O(N__39264),
            .I(N__39232));
    LocalMux I__5971 (
            .O(N__39257),
            .I(N__39229));
    Span4Mux_v I__5970 (
            .O(N__39252),
            .I(N__39224));
    LocalMux I__5969 (
            .O(N__39235),
            .I(N__39224));
    Span4Mux_v I__5968 (
            .O(N__39232),
            .I(N__39219));
    Span4Mux_v I__5967 (
            .O(N__39229),
            .I(N__39219));
    Span4Mux_h I__5966 (
            .O(N__39224),
            .I(N__39216));
    Odrv4 I__5965 (
            .O(N__39219),
            .I(\foc.u_Park_Transform.dCurrent_2 ));
    Odrv4 I__5964 (
            .O(N__39216),
            .I(\foc.u_Park_Transform.dCurrent_2 ));
    InMux I__5963 (
            .O(N__39211),
            .I(N__39208));
    LocalMux I__5962 (
            .O(N__39208),
            .I(N__39205));
    Odrv4 I__5961 (
            .O(N__39205),
            .I(\foc.u_Park_Transform.Product1_mul_temp_14 ));
    InMux I__5960 (
            .O(N__39202),
            .I(\foc.u_Park_Transform.n17263 ));
    InMux I__5959 (
            .O(N__39199),
            .I(N__39196));
    LocalMux I__5958 (
            .O(N__39196),
            .I(N__39192));
    InMux I__5957 (
            .O(N__39195),
            .I(N__39189));
    Span4Mux_v I__5956 (
            .O(N__39192),
            .I(N__39186));
    LocalMux I__5955 (
            .O(N__39189),
            .I(N__39183));
    Span4Mux_h I__5954 (
            .O(N__39186),
            .I(N__39178));
    Span4Mux_h I__5953 (
            .O(N__39183),
            .I(N__39178));
    Odrv4 I__5952 (
            .O(N__39178),
            .I(\foc.u_Park_Transform.n737 ));
    InMux I__5951 (
            .O(N__39175),
            .I(N__39172));
    LocalMux I__5950 (
            .O(N__39172),
            .I(N__39169));
    Odrv4 I__5949 (
            .O(N__39169),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n2 ));
    InMux I__5948 (
            .O(N__39166),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15804 ));
    InMux I__5947 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__5946 (
            .O(N__39160),
            .I(\foc.dCurrent_26 ));
    InMux I__5945 (
            .O(N__39157),
            .I(N__39154));
    LocalMux I__5944 (
            .O(N__39154),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n7 ));
    InMux I__5943 (
            .O(N__39151),
            .I(N__39148));
    LocalMux I__5942 (
            .O(N__39148),
            .I(N__39145));
    Span4Mux_v I__5941 (
            .O(N__39145),
            .I(N__39142));
    Odrv4 I__5940 (
            .O(N__39142),
            .I(\foc.dCurrent_3 ));
    InMux I__5939 (
            .O(N__39139),
            .I(N__39136));
    LocalMux I__5938 (
            .O(N__39136),
            .I(N__39133));
    Odrv4 I__5937 (
            .O(N__39133),
            .I(\foc.u_Park_Transform.Product1_mul_temp_2 ));
    InMux I__5936 (
            .O(N__39130),
            .I(\foc.u_Park_Transform.n17251 ));
    InMux I__5935 (
            .O(N__39127),
            .I(N__39124));
    LocalMux I__5934 (
            .O(N__39124),
            .I(N__39121));
    Odrv4 I__5933 (
            .O(N__39121),
            .I(\foc.u_Park_Transform.Product1_mul_temp_3 ));
    InMux I__5932 (
            .O(N__39118),
            .I(\foc.u_Park_Transform.n17252 ));
    InMux I__5931 (
            .O(N__39115),
            .I(N__39112));
    LocalMux I__5930 (
            .O(N__39112),
            .I(N__39109));
    Odrv4 I__5929 (
            .O(N__39109),
            .I(\foc.u_Park_Transform.Product1_mul_temp_4 ));
    InMux I__5928 (
            .O(N__39106),
            .I(\foc.u_Park_Transform.n17253 ));
    InMux I__5927 (
            .O(N__39103),
            .I(N__39100));
    LocalMux I__5926 (
            .O(N__39100),
            .I(N__39097));
    Odrv4 I__5925 (
            .O(N__39097),
            .I(\foc.u_Park_Transform.Product1_mul_temp_5 ));
    InMux I__5924 (
            .O(N__39094),
            .I(\foc.u_Park_Transform.n17254 ));
    InMux I__5923 (
            .O(N__39091),
            .I(N__39088));
    LocalMux I__5922 (
            .O(N__39088),
            .I(N__39085));
    Odrv4 I__5921 (
            .O(N__39085),
            .I(\foc.u_Park_Transform.Product1_mul_temp_6 ));
    InMux I__5920 (
            .O(N__39082),
            .I(\foc.u_Park_Transform.n17255 ));
    InMux I__5919 (
            .O(N__39079),
            .I(N__39076));
    LocalMux I__5918 (
            .O(N__39076),
            .I(N__39073));
    Span4Mux_v I__5917 (
            .O(N__39073),
            .I(N__39070));
    Odrv4 I__5916 (
            .O(N__39070),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n11 ));
    InMux I__5915 (
            .O(N__39067),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15795 ));
    InMux I__5914 (
            .O(N__39064),
            .I(N__39061));
    LocalMux I__5913 (
            .O(N__39061),
            .I(N__39058));
    Span4Mux_h I__5912 (
            .O(N__39058),
            .I(N__39055));
    Odrv4 I__5911 (
            .O(N__39055),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n10 ));
    InMux I__5910 (
            .O(N__39052),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15796 ));
    InMux I__5909 (
            .O(N__39049),
            .I(N__39046));
    LocalMux I__5908 (
            .O(N__39046),
            .I(N__39043));
    Span4Mux_h I__5907 (
            .O(N__39043),
            .I(N__39040));
    Odrv4 I__5906 (
            .O(N__39040),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n9 ));
    InMux I__5905 (
            .O(N__39037),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15797 ));
    InMux I__5904 (
            .O(N__39034),
            .I(N__39031));
    LocalMux I__5903 (
            .O(N__39031),
            .I(N__39028));
    Odrv4 I__5902 (
            .O(N__39028),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n8 ));
    InMux I__5901 (
            .O(N__39025),
            .I(bfn_15_8_0_));
    InMux I__5900 (
            .O(N__39022),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15799 ));
    InMux I__5899 (
            .O(N__39019),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15800 ));
    InMux I__5898 (
            .O(N__39016),
            .I(N__39013));
    LocalMux I__5897 (
            .O(N__39013),
            .I(N__39010));
    Odrv4 I__5896 (
            .O(N__39010),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n5 ));
    InMux I__5895 (
            .O(N__39007),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15801 ));
    InMux I__5894 (
            .O(N__39004),
            .I(N__39001));
    LocalMux I__5893 (
            .O(N__39001),
            .I(N__38998));
    Odrv4 I__5892 (
            .O(N__38998),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515 ));
    InMux I__5891 (
            .O(N__38995),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15802 ));
    InMux I__5890 (
            .O(N__38992),
            .I(N__38989));
    LocalMux I__5889 (
            .O(N__38989),
            .I(N__38986));
    Odrv4 I__5888 (
            .O(N__38986),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n3 ));
    InMux I__5887 (
            .O(N__38983),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15803 ));
    InMux I__5886 (
            .O(N__38980),
            .I(N__38977));
    LocalMux I__5885 (
            .O(N__38977),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n19 ));
    InMux I__5884 (
            .O(N__38974),
            .I(N__38971));
    LocalMux I__5883 (
            .O(N__38971),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n18 ));
    InMux I__5882 (
            .O(N__38968),
            .I(N__38965));
    LocalMux I__5881 (
            .O(N__38965),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n17 ));
    InMux I__5880 (
            .O(N__38962),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15789 ));
    InMux I__5879 (
            .O(N__38959),
            .I(N__38956));
    LocalMux I__5878 (
            .O(N__38956),
            .I(N__38953));
    Span4Mux_h I__5877 (
            .O(N__38953),
            .I(N__38950));
    Odrv4 I__5876 (
            .O(N__38950),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n16 ));
    InMux I__5875 (
            .O(N__38947),
            .I(bfn_15_7_0_));
    InMux I__5874 (
            .O(N__38944),
            .I(N__38941));
    LocalMux I__5873 (
            .O(N__38941),
            .I(N__38938));
    Odrv4 I__5872 (
            .O(N__38938),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518 ));
    InMux I__5871 (
            .O(N__38935),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15791 ));
    InMux I__5870 (
            .O(N__38932),
            .I(N__38929));
    LocalMux I__5869 (
            .O(N__38929),
            .I(N__38926));
    Span4Mux_h I__5868 (
            .O(N__38926),
            .I(N__38923));
    Odrv4 I__5867 (
            .O(N__38923),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517 ));
    InMux I__5866 (
            .O(N__38920),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15792 ));
    InMux I__5865 (
            .O(N__38917),
            .I(N__38914));
    LocalMux I__5864 (
            .O(N__38914),
            .I(N__38911));
    Span4Mux_h I__5863 (
            .O(N__38911),
            .I(N__38908));
    Odrv4 I__5862 (
            .O(N__38908),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n13 ));
    InMux I__5861 (
            .O(N__38905),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15793 ));
    InMux I__5860 (
            .O(N__38902),
            .I(N__38899));
    LocalMux I__5859 (
            .O(N__38899),
            .I(N__38896));
    Span4Mux_v I__5858 (
            .O(N__38896),
            .I(N__38893));
    Odrv4 I__5857 (
            .O(N__38893),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516 ));
    InMux I__5856 (
            .O(N__38890),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n15794 ));
    InMux I__5855 (
            .O(N__38887),
            .I(N__38884));
    LocalMux I__5854 (
            .O(N__38884),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n28 ));
    InMux I__5853 (
            .O(N__38881),
            .I(N__38878));
    LocalMux I__5852 (
            .O(N__38878),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n27 ));
    InMux I__5851 (
            .O(N__38875),
            .I(N__38872));
    LocalMux I__5850 (
            .O(N__38872),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n26 ));
    InMux I__5849 (
            .O(N__38869),
            .I(N__38866));
    LocalMux I__5848 (
            .O(N__38866),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n25 ));
    InMux I__5847 (
            .O(N__38863),
            .I(N__38860));
    LocalMux I__5846 (
            .O(N__38860),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n24 ));
    InMux I__5845 (
            .O(N__38857),
            .I(N__38854));
    LocalMux I__5844 (
            .O(N__38854),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n23 ));
    InMux I__5843 (
            .O(N__38851),
            .I(N__38848));
    LocalMux I__5842 (
            .O(N__38848),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n22 ));
    InMux I__5841 (
            .O(N__38845),
            .I(N__38842));
    LocalMux I__5840 (
            .O(N__38842),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n21 ));
    InMux I__5839 (
            .O(N__38839),
            .I(N__38836));
    LocalMux I__5838 (
            .O(N__38836),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n20 ));
    InMux I__5837 (
            .O(N__38833),
            .I(N__38830));
    LocalMux I__5836 (
            .O(N__38830),
            .I(N__38827));
    Odrv4 I__5835 (
            .O(N__38827),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671 ));
    InMux I__5834 (
            .O(N__38824),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18043 ));
    CascadeMux I__5833 (
            .O(N__38821),
            .I(N__38818));
    InMux I__5832 (
            .O(N__38818),
            .I(N__38815));
    LocalMux I__5831 (
            .O(N__38815),
            .I(N__38812));
    Odrv12 I__5830 (
            .O(N__38812),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670 ));
    InMux I__5829 (
            .O(N__38809),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18044 ));
    CascadeMux I__5828 (
            .O(N__38806),
            .I(N__38803));
    InMux I__5827 (
            .O(N__38803),
            .I(N__38800));
    LocalMux I__5826 (
            .O(N__38800),
            .I(N__38797));
    Odrv4 I__5825 (
            .O(N__38797),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669 ));
    InMux I__5824 (
            .O(N__38794),
            .I(N__38791));
    LocalMux I__5823 (
            .O(N__38791),
            .I(N__38788));
    Span4Mux_v I__5822 (
            .O(N__38788),
            .I(N__38785));
    Odrv4 I__5821 (
            .O(N__38785),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683 ));
    InMux I__5820 (
            .O(N__38782),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18045 ));
    InMux I__5819 (
            .O(N__38779),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684 ));
    CascadeMux I__5818 (
            .O(N__38776),
            .I(N__38773));
    InMux I__5817 (
            .O(N__38773),
            .I(N__38770));
    LocalMux I__5816 (
            .O(N__38770),
            .I(N__38767));
    Span4Mux_v I__5815 (
            .O(N__38767),
            .I(N__38764));
    Odrv4 I__5814 (
            .O(N__38764),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO ));
    InMux I__5813 (
            .O(N__38761),
            .I(N__38758));
    LocalMux I__5812 (
            .O(N__38758),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n30 ));
    InMux I__5811 (
            .O(N__38755),
            .I(N__38752));
    LocalMux I__5810 (
            .O(N__38752),
            .I(\foc.u_DQ_Current_Control.u_D_Current_Control.n29 ));
    InMux I__5809 (
            .O(N__38749),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18034 ));
    InMux I__5808 (
            .O(N__38746),
            .I(N__38743));
    LocalMux I__5807 (
            .O(N__38743),
            .I(N__38740));
    Odrv12 I__5806 (
            .O(N__38740),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679 ));
    InMux I__5805 (
            .O(N__38737),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18035 ));
    CascadeMux I__5804 (
            .O(N__38734),
            .I(N__38731));
    InMux I__5803 (
            .O(N__38731),
            .I(N__38728));
    LocalMux I__5802 (
            .O(N__38728),
            .I(N__38725));
    Odrv4 I__5801 (
            .O(N__38725),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678 ));
    InMux I__5800 (
            .O(N__38722),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18036 ));
    InMux I__5799 (
            .O(N__38719),
            .I(N__38716));
    LocalMux I__5798 (
            .O(N__38716),
            .I(N__38713));
    Odrv12 I__5797 (
            .O(N__38713),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677 ));
    InMux I__5796 (
            .O(N__38710),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18037 ));
    CascadeMux I__5795 (
            .O(N__38707),
            .I(N__38704));
    InMux I__5794 (
            .O(N__38704),
            .I(N__38701));
    LocalMux I__5793 (
            .O(N__38701),
            .I(N__38698));
    Odrv4 I__5792 (
            .O(N__38698),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676 ));
    InMux I__5791 (
            .O(N__38695),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18038 ));
    InMux I__5790 (
            .O(N__38692),
            .I(N__38689));
    LocalMux I__5789 (
            .O(N__38689),
            .I(N__38686));
    Odrv12 I__5788 (
            .O(N__38686),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675 ));
    InMux I__5787 (
            .O(N__38683),
            .I(bfn_14_26_0_));
    CascadeMux I__5786 (
            .O(N__38680),
            .I(N__38677));
    InMux I__5785 (
            .O(N__38677),
            .I(N__38674));
    LocalMux I__5784 (
            .O(N__38674),
            .I(N__38671));
    Odrv4 I__5783 (
            .O(N__38671),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674 ));
    InMux I__5782 (
            .O(N__38668),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18040 ));
    InMux I__5781 (
            .O(N__38665),
            .I(N__38662));
    LocalMux I__5780 (
            .O(N__38662),
            .I(N__38659));
    Odrv4 I__5779 (
            .O(N__38659),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673 ));
    InMux I__5778 (
            .O(N__38656),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18041 ));
    CascadeMux I__5777 (
            .O(N__38653),
            .I(N__38650));
    InMux I__5776 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__5775 (
            .O(N__38647),
            .I(N__38644));
    Odrv12 I__5774 (
            .O(N__38644),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672 ));
    InMux I__5773 (
            .O(N__38641),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18042 ));
    InMux I__5772 (
            .O(N__38638),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18057 ));
    InMux I__5771 (
            .O(N__38635),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18058 ));
    InMux I__5770 (
            .O(N__38632),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18059 ));
    InMux I__5769 (
            .O(N__38629),
            .I(N__38626));
    LocalMux I__5768 (
            .O(N__38626),
            .I(N__38623));
    Odrv4 I__5767 (
            .O(N__38623),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667 ));
    InMux I__5766 (
            .O(N__38620),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18060 ));
    InMux I__5765 (
            .O(N__38617),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668 ));
    CascadeMux I__5764 (
            .O(N__38614),
            .I(N__38611));
    InMux I__5763 (
            .O(N__38611),
            .I(N__38608));
    LocalMux I__5762 (
            .O(N__38608),
            .I(N__38605));
    Odrv4 I__5761 (
            .O(N__38605),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO ));
    CascadeMux I__5760 (
            .O(N__38602),
            .I(N__38599));
    InMux I__5759 (
            .O(N__38599),
            .I(N__38596));
    LocalMux I__5758 (
            .O(N__38596),
            .I(N__38593));
    Odrv4 I__5757 (
            .O(N__38593),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682 ));
    InMux I__5756 (
            .O(N__38590),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18032 ));
    InMux I__5755 (
            .O(N__38587),
            .I(N__38584));
    LocalMux I__5754 (
            .O(N__38584),
            .I(N__38581));
    Odrv4 I__5753 (
            .O(N__38581),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681 ));
    InMux I__5752 (
            .O(N__38578),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18033 ));
    CascadeMux I__5751 (
            .O(N__38575),
            .I(N__38572));
    InMux I__5750 (
            .O(N__38572),
            .I(N__38569));
    LocalMux I__5749 (
            .O(N__38569),
            .I(N__38566));
    Odrv12 I__5748 (
            .O(N__38566),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680 ));
    InMux I__5747 (
            .O(N__38563),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18048 ));
    InMux I__5746 (
            .O(N__38560),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18049 ));
    InMux I__5745 (
            .O(N__38557),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18050 ));
    InMux I__5744 (
            .O(N__38554),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18051 ));
    InMux I__5743 (
            .O(N__38551),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18052 ));
    InMux I__5742 (
            .O(N__38548),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18053 ));
    InMux I__5741 (
            .O(N__38545),
            .I(bfn_14_24_0_));
    InMux I__5740 (
            .O(N__38542),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18055 ));
    InMux I__5739 (
            .O(N__38539),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18056 ));
    CascadeMux I__5738 (
            .O(N__38536),
            .I(N__38533));
    InMux I__5737 (
            .O(N__38533),
            .I(N__38530));
    LocalMux I__5736 (
            .O(N__38530),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743 ));
    InMux I__5735 (
            .O(N__38527),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17730 ));
    InMux I__5734 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__5733 (
            .O(N__38521),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740 ));
    InMux I__5732 (
            .O(N__38518),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17731 ));
    CascadeMux I__5731 (
            .O(N__38515),
            .I(N__38512));
    InMux I__5730 (
            .O(N__38512),
            .I(N__38509));
    LocalMux I__5729 (
            .O(N__38509),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739 ));
    InMux I__5728 (
            .O(N__38506),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17732 ));
    CascadeMux I__5727 (
            .O(N__38503),
            .I(N__38499));
    CascadeMux I__5726 (
            .O(N__38502),
            .I(N__38496));
    InMux I__5725 (
            .O(N__38499),
            .I(N__38492));
    InMux I__5724 (
            .O(N__38496),
            .I(N__38487));
    InMux I__5723 (
            .O(N__38495),
            .I(N__38487));
    LocalMux I__5722 (
            .O(N__38492),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738 ));
    LocalMux I__5721 (
            .O(N__38487),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738 ));
    InMux I__5720 (
            .O(N__38482),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17733 ));
    InMux I__5719 (
            .O(N__38479),
            .I(N__38476));
    LocalMux I__5718 (
            .O(N__38476),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735 ));
    InMux I__5717 (
            .O(N__38473),
            .I(bfn_14_22_0_));
    InMux I__5716 (
            .O(N__38470),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734 ));
    CascadeMux I__5715 (
            .O(N__38467),
            .I(N__38464));
    InMux I__5714 (
            .O(N__38464),
            .I(N__38461));
    LocalMux I__5713 (
            .O(N__38461),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO ));
    InMux I__5712 (
            .O(N__38458),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18047 ));
    InMux I__5711 (
            .O(N__38455),
            .I(N__38452));
    LocalMux I__5710 (
            .O(N__38452),
            .I(N__38449));
    Span4Mux_v I__5709 (
            .O(N__38449),
            .I(N__38446));
    Odrv4 I__5708 (
            .O(N__38446),
            .I(\foc.u_Park_Transform.Product4_mul_temp_29 ));
    InMux I__5707 (
            .O(N__38443),
            .I(\foc.u_Park_Transform.n15774 ));
    InMux I__5706 (
            .O(N__38440),
            .I(N__38437));
    LocalMux I__5705 (
            .O(N__38437),
            .I(\foc.qCurrent_21 ));
    InMux I__5704 (
            .O(N__38434),
            .I(N__38431));
    LocalMux I__5703 (
            .O(N__38431),
            .I(\foc.qCurrent_29 ));
    InMux I__5702 (
            .O(N__38428),
            .I(N__38425));
    LocalMux I__5701 (
            .O(N__38425),
            .I(\foc.qCurrent_23 ));
    InMux I__5700 (
            .O(N__38422),
            .I(N__38419));
    LocalMux I__5699 (
            .O(N__38419),
            .I(\foc.qCurrent_30 ));
    CascadeMux I__5698 (
            .O(N__38416),
            .I(N__38413));
    InMux I__5697 (
            .O(N__38413),
            .I(N__38410));
    LocalMux I__5696 (
            .O(N__38410),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749 ));
    InMux I__5695 (
            .O(N__38407),
            .I(N__38404));
    LocalMux I__5694 (
            .O(N__38404),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747 ));
    InMux I__5693 (
            .O(N__38401),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17727 ));
    CascadeMux I__5692 (
            .O(N__38398),
            .I(N__38395));
    InMux I__5691 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__5690 (
            .O(N__38392),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745 ));
    InMux I__5689 (
            .O(N__38389),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17728 ));
    InMux I__5688 (
            .O(N__38386),
            .I(N__38383));
    LocalMux I__5687 (
            .O(N__38383),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744 ));
    InMux I__5686 (
            .O(N__38380),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17729 ));
    CascadeMux I__5685 (
            .O(N__38377),
            .I(N__38374));
    InMux I__5684 (
            .O(N__38374),
            .I(N__38371));
    LocalMux I__5683 (
            .O(N__38371),
            .I(N__38368));
    Span4Mux_h I__5682 (
            .O(N__38368),
            .I(N__38365));
    Odrv4 I__5681 (
            .O(N__38365),
            .I(\foc.u_Park_Transform.Product4_mul_temp_21 ));
    InMux I__5680 (
            .O(N__38362),
            .I(\foc.u_Park_Transform.n15766 ));
    InMux I__5679 (
            .O(N__38359),
            .I(N__38356));
    LocalMux I__5678 (
            .O(N__38356),
            .I(N__38353));
    Span4Mux_v I__5677 (
            .O(N__38353),
            .I(N__38350));
    Odrv4 I__5676 (
            .O(N__38350),
            .I(\foc.u_Park_Transform.Product4_mul_temp_22 ));
    InMux I__5675 (
            .O(N__38347),
            .I(\foc.u_Park_Transform.n15767 ));
    CascadeMux I__5674 (
            .O(N__38344),
            .I(N__38341));
    InMux I__5673 (
            .O(N__38341),
            .I(N__38338));
    LocalMux I__5672 (
            .O(N__38338),
            .I(N__38335));
    Span4Mux_h I__5671 (
            .O(N__38335),
            .I(N__38332));
    Odrv4 I__5670 (
            .O(N__38332),
            .I(\foc.u_Park_Transform.Product4_mul_temp_23 ));
    InMux I__5669 (
            .O(N__38329),
            .I(\foc.u_Park_Transform.n15768 ));
    InMux I__5668 (
            .O(N__38326),
            .I(N__38323));
    LocalMux I__5667 (
            .O(N__38323),
            .I(N__38320));
    Span4Mux_h I__5666 (
            .O(N__38320),
            .I(N__38317));
    Odrv4 I__5665 (
            .O(N__38317),
            .I(\foc.u_Park_Transform.Product4_mul_temp_24 ));
    InMux I__5664 (
            .O(N__38314),
            .I(\foc.u_Park_Transform.n15769 ));
    CascadeMux I__5663 (
            .O(N__38311),
            .I(N__38308));
    InMux I__5662 (
            .O(N__38308),
            .I(N__38305));
    LocalMux I__5661 (
            .O(N__38305),
            .I(N__38302));
    Span4Mux_v I__5660 (
            .O(N__38302),
            .I(N__38299));
    Odrv4 I__5659 (
            .O(N__38299),
            .I(\foc.u_Park_Transform.Product4_mul_temp_25 ));
    InMux I__5658 (
            .O(N__38296),
            .I(\foc.u_Park_Transform.n15770 ));
    InMux I__5657 (
            .O(N__38293),
            .I(N__38290));
    LocalMux I__5656 (
            .O(N__38290),
            .I(N__38287));
    Span4Mux_h I__5655 (
            .O(N__38287),
            .I(N__38284));
    Odrv4 I__5654 (
            .O(N__38284),
            .I(\foc.u_Park_Transform.Product4_mul_temp_26 ));
    InMux I__5653 (
            .O(N__38281),
            .I(bfn_14_20_0_));
    CascadeMux I__5652 (
            .O(N__38278),
            .I(N__38275));
    InMux I__5651 (
            .O(N__38275),
            .I(N__38272));
    LocalMux I__5650 (
            .O(N__38272),
            .I(N__38269));
    Span4Mux_v I__5649 (
            .O(N__38269),
            .I(N__38266));
    Odrv4 I__5648 (
            .O(N__38266),
            .I(\foc.u_Park_Transform.Product4_mul_temp_27 ));
    InMux I__5647 (
            .O(N__38263),
            .I(\foc.u_Park_Transform.n15772 ));
    InMux I__5646 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__5645 (
            .O(N__38257),
            .I(N__38254));
    Span4Mux_h I__5644 (
            .O(N__38254),
            .I(N__38251));
    Odrv4 I__5643 (
            .O(N__38251),
            .I(\foc.u_Park_Transform.Product4_mul_temp_28 ));
    InMux I__5642 (
            .O(N__38248),
            .I(\foc.u_Park_Transform.n15773 ));
    InMux I__5641 (
            .O(N__38245),
            .I(N__38242));
    LocalMux I__5640 (
            .O(N__38242),
            .I(N__38239));
    Odrv12 I__5639 (
            .O(N__38239),
            .I(\foc.u_Park_Transform.Product4_mul_temp_12 ));
    InMux I__5638 (
            .O(N__38236),
            .I(\foc.u_Park_Transform.n15757 ));
    CascadeMux I__5637 (
            .O(N__38233),
            .I(N__38230));
    InMux I__5636 (
            .O(N__38230),
            .I(N__38227));
    LocalMux I__5635 (
            .O(N__38227),
            .I(N__38224));
    Odrv4 I__5634 (
            .O(N__38224),
            .I(\foc.u_Park_Transform.Product4_mul_temp_13 ));
    InMux I__5633 (
            .O(N__38221),
            .I(\foc.u_Park_Transform.n15758 ));
    InMux I__5632 (
            .O(N__38218),
            .I(N__38215));
    LocalMux I__5631 (
            .O(N__38215),
            .I(N__38212));
    Odrv4 I__5630 (
            .O(N__38212),
            .I(\foc.u_Park_Transform.Product4_mul_temp_14 ));
    InMux I__5629 (
            .O(N__38209),
            .I(\foc.u_Park_Transform.n15759 ));
    CascadeMux I__5628 (
            .O(N__38206),
            .I(N__38203));
    InMux I__5627 (
            .O(N__38203),
            .I(N__38200));
    LocalMux I__5626 (
            .O(N__38200),
            .I(N__38197));
    Span4Mux_v I__5625 (
            .O(N__38197),
            .I(N__38194));
    Odrv4 I__5624 (
            .O(N__38194),
            .I(\foc.u_Park_Transform.Product4_mul_temp_15 ));
    InMux I__5623 (
            .O(N__38191),
            .I(\foc.u_Park_Transform.n15760 ));
    InMux I__5622 (
            .O(N__38188),
            .I(N__38185));
    LocalMux I__5621 (
            .O(N__38185),
            .I(N__38182));
    Span4Mux_h I__5620 (
            .O(N__38182),
            .I(N__38179));
    Odrv4 I__5619 (
            .O(N__38179),
            .I(\foc.u_Park_Transform.Product4_mul_temp_16 ));
    InMux I__5618 (
            .O(N__38176),
            .I(\foc.u_Park_Transform.n15761 ));
    CascadeMux I__5617 (
            .O(N__38173),
            .I(N__38170));
    InMux I__5616 (
            .O(N__38170),
            .I(N__38167));
    LocalMux I__5615 (
            .O(N__38167),
            .I(N__38164));
    Span4Mux_h I__5614 (
            .O(N__38164),
            .I(N__38161));
    Odrv4 I__5613 (
            .O(N__38161),
            .I(\foc.u_Park_Transform.Product4_mul_temp_17 ));
    InMux I__5612 (
            .O(N__38158),
            .I(\foc.u_Park_Transform.n15762 ));
    InMux I__5611 (
            .O(N__38155),
            .I(N__38152));
    LocalMux I__5610 (
            .O(N__38152),
            .I(N__38149));
    Span4Mux_h I__5609 (
            .O(N__38149),
            .I(N__38146));
    Odrv4 I__5608 (
            .O(N__38146),
            .I(\foc.u_Park_Transform.Product4_mul_temp_18 ));
    InMux I__5607 (
            .O(N__38143),
            .I(bfn_14_19_0_));
    CascadeMux I__5606 (
            .O(N__38140),
            .I(N__38137));
    InMux I__5605 (
            .O(N__38137),
            .I(N__38134));
    LocalMux I__5604 (
            .O(N__38134),
            .I(N__38131));
    Span4Mux_v I__5603 (
            .O(N__38131),
            .I(N__38128));
    Odrv4 I__5602 (
            .O(N__38128),
            .I(\foc.u_Park_Transform.Product4_mul_temp_19 ));
    InMux I__5601 (
            .O(N__38125),
            .I(\foc.u_Park_Transform.n15764 ));
    InMux I__5600 (
            .O(N__38122),
            .I(N__38119));
    LocalMux I__5599 (
            .O(N__38119),
            .I(N__38116));
    Span4Mux_h I__5598 (
            .O(N__38116),
            .I(N__38113));
    Odrv4 I__5597 (
            .O(N__38113),
            .I(\foc.u_Park_Transform.Product4_mul_temp_20 ));
    InMux I__5596 (
            .O(N__38110),
            .I(\foc.u_Park_Transform.n15765 ));
    InMux I__5595 (
            .O(N__38107),
            .I(N__38104));
    LocalMux I__5594 (
            .O(N__38104),
            .I(N__38101));
    Odrv4 I__5593 (
            .O(N__38101),
            .I(\foc.u_Park_Transform.Product4_mul_temp_4 ));
    InMux I__5592 (
            .O(N__38098),
            .I(\foc.u_Park_Transform.n15749 ));
    InMux I__5591 (
            .O(N__38095),
            .I(N__38092));
    LocalMux I__5590 (
            .O(N__38092),
            .I(N__38089));
    Odrv4 I__5589 (
            .O(N__38089),
            .I(\foc.u_Park_Transform.Product4_mul_temp_5 ));
    InMux I__5588 (
            .O(N__38086),
            .I(\foc.u_Park_Transform.n15750 ));
    InMux I__5587 (
            .O(N__38083),
            .I(N__38080));
    LocalMux I__5586 (
            .O(N__38080),
            .I(N__38077));
    Odrv4 I__5585 (
            .O(N__38077),
            .I(\foc.u_Park_Transform.Product4_mul_temp_6 ));
    InMux I__5584 (
            .O(N__38074),
            .I(\foc.u_Park_Transform.n15751 ));
    InMux I__5583 (
            .O(N__38071),
            .I(N__38068));
    LocalMux I__5582 (
            .O(N__38068),
            .I(N__38065));
    Odrv4 I__5581 (
            .O(N__38065),
            .I(\foc.u_Park_Transform.Product4_mul_temp_7 ));
    InMux I__5580 (
            .O(N__38062),
            .I(\foc.u_Park_Transform.n15752 ));
    InMux I__5579 (
            .O(N__38059),
            .I(N__38056));
    LocalMux I__5578 (
            .O(N__38056),
            .I(N__38053));
    Odrv12 I__5577 (
            .O(N__38053),
            .I(\foc.u_Park_Transform.Product4_mul_temp_8 ));
    InMux I__5576 (
            .O(N__38050),
            .I(\foc.u_Park_Transform.n15753 ));
    CascadeMux I__5575 (
            .O(N__38047),
            .I(N__38044));
    InMux I__5574 (
            .O(N__38044),
            .I(N__38041));
    LocalMux I__5573 (
            .O(N__38041),
            .I(\foc.u_Park_Transform.Product4_mul_temp_9 ));
    InMux I__5572 (
            .O(N__38038),
            .I(\foc.u_Park_Transform.n15754 ));
    InMux I__5571 (
            .O(N__38035),
            .I(N__38032));
    LocalMux I__5570 (
            .O(N__38032),
            .I(N__38029));
    Odrv4 I__5569 (
            .O(N__38029),
            .I(\foc.u_Park_Transform.Product4_mul_temp_10 ));
    InMux I__5568 (
            .O(N__38026),
            .I(bfn_14_18_0_));
    CascadeMux I__5567 (
            .O(N__38023),
            .I(N__38020));
    InMux I__5566 (
            .O(N__38020),
            .I(N__38017));
    LocalMux I__5565 (
            .O(N__38017),
            .I(N__38014));
    Odrv12 I__5564 (
            .O(N__38014),
            .I(\foc.u_Park_Transform.Product4_mul_temp_11 ));
    InMux I__5563 (
            .O(N__38011),
            .I(\foc.u_Park_Transform.n15756 ));
    InMux I__5562 (
            .O(N__38008),
            .I(\foc.u_Park_Transform.n17076 ));
    InMux I__5561 (
            .O(N__38005),
            .I(\foc.u_Park_Transform.n17077 ));
    InMux I__5560 (
            .O(N__38002),
            .I(\foc.u_Park_Transform.n17078 ));
    InMux I__5559 (
            .O(N__37999),
            .I(\foc.u_Park_Transform.n17079 ));
    InMux I__5558 (
            .O(N__37996),
            .I(\foc.u_Park_Transform.n17080 ));
    CascadeMux I__5557 (
            .O(N__37993),
            .I(N__37990));
    InMux I__5556 (
            .O(N__37990),
            .I(N__37986));
    InMux I__5555 (
            .O(N__37989),
            .I(N__37983));
    LocalMux I__5554 (
            .O(N__37986),
            .I(N__37978));
    LocalMux I__5553 (
            .O(N__37983),
            .I(N__37978));
    Span4Mux_v I__5552 (
            .O(N__37978),
            .I(N__37975));
    Odrv4 I__5551 (
            .O(N__37975),
            .I(\foc.u_Park_Transform.n738_adj_2003 ));
    InMux I__5550 (
            .O(N__37972),
            .I(\foc.u_Park_Transform.n17081 ));
    InMux I__5549 (
            .O(N__37969),
            .I(\foc.u_Park_Transform.n739_adj_2006 ));
    CascadeMux I__5548 (
            .O(N__37966),
            .I(N__37963));
    InMux I__5547 (
            .O(N__37963),
            .I(N__37960));
    LocalMux I__5546 (
            .O(N__37960),
            .I(N__37957));
    Span4Mux_v I__5545 (
            .O(N__37957),
            .I(N__37954));
    Odrv4 I__5544 (
            .O(N__37954),
            .I(\foc.u_Park_Transform.n739_adj_2006_THRU_CO ));
    InMux I__5543 (
            .O(N__37951),
            .I(N__37948));
    LocalMux I__5542 (
            .O(N__37948),
            .I(N__37945));
    Odrv4 I__5541 (
            .O(N__37945),
            .I(\foc.u_Park_Transform.Product4_mul_temp_2 ));
    InMux I__5540 (
            .O(N__37942),
            .I(bfn_14_17_0_));
    InMux I__5539 (
            .O(N__37939),
            .I(N__37936));
    LocalMux I__5538 (
            .O(N__37936),
            .I(N__37933));
    Odrv4 I__5537 (
            .O(N__37933),
            .I(\foc.u_Park_Transform.Product4_mul_temp_3 ));
    InMux I__5536 (
            .O(N__37930),
            .I(\foc.u_Park_Transform.n15748 ));
    InMux I__5535 (
            .O(N__37927),
            .I(\foc.u_Park_Transform.n17068 ));
    InMux I__5534 (
            .O(N__37924),
            .I(\foc.u_Park_Transform.n17069 ));
    InMux I__5533 (
            .O(N__37921),
            .I(\foc.u_Park_Transform.n17070 ));
    InMux I__5532 (
            .O(N__37918),
            .I(\foc.u_Park_Transform.n17071 ));
    InMux I__5531 (
            .O(N__37915),
            .I(\foc.u_Park_Transform.n17072 ));
    InMux I__5530 (
            .O(N__37912),
            .I(\foc.u_Park_Transform.n17073 ));
    InMux I__5529 (
            .O(N__37909),
            .I(\foc.u_Park_Transform.n17074 ));
    InMux I__5528 (
            .O(N__37906),
            .I(bfn_14_16_0_));
    CascadeMux I__5527 (
            .O(N__37903),
            .I(N__37900));
    InMux I__5526 (
            .O(N__37900),
            .I(N__37897));
    LocalMux I__5525 (
            .O(N__37897),
            .I(\foc.u_Park_Transform.n409_adj_1997 ));
    InMux I__5524 (
            .O(N__37894),
            .I(bfn_14_14_0_));
    InMux I__5523 (
            .O(N__37891),
            .I(N__37888));
    LocalMux I__5522 (
            .O(N__37888),
            .I(\foc.u_Park_Transform.n458_adj_2093 ));
    InMux I__5521 (
            .O(N__37885),
            .I(\foc.u_Park_Transform.n17016 ));
    CascadeMux I__5520 (
            .O(N__37882),
            .I(N__37879));
    InMux I__5519 (
            .O(N__37879),
            .I(N__37876));
    LocalMux I__5518 (
            .O(N__37876),
            .I(\foc.u_Park_Transform.n507 ));
    InMux I__5517 (
            .O(N__37873),
            .I(\foc.u_Park_Transform.n17017 ));
    InMux I__5516 (
            .O(N__37870),
            .I(N__37867));
    LocalMux I__5515 (
            .O(N__37867),
            .I(\foc.u_Park_Transform.n556 ));
    InMux I__5514 (
            .O(N__37864),
            .I(\foc.u_Park_Transform.n17018 ));
    CascadeMux I__5513 (
            .O(N__37861),
            .I(N__37858));
    InMux I__5512 (
            .O(N__37858),
            .I(N__37855));
    LocalMux I__5511 (
            .O(N__37855),
            .I(\foc.u_Park_Transform.n605 ));
    InMux I__5510 (
            .O(N__37852),
            .I(\foc.u_Park_Transform.n17019 ));
    InMux I__5509 (
            .O(N__37849),
            .I(N__37846));
    LocalMux I__5508 (
            .O(N__37846),
            .I(\foc.u_Park_Transform.n654 ));
    InMux I__5507 (
            .O(N__37843),
            .I(\foc.u_Park_Transform.n17020 ));
    InMux I__5506 (
            .O(N__37840),
            .I(N__37837));
    LocalMux I__5505 (
            .O(N__37837),
            .I(N__37834));
    Span4Mux_v I__5504 (
            .O(N__37834),
            .I(N__37830));
    InMux I__5503 (
            .O(N__37833),
            .I(N__37827));
    Odrv4 I__5502 (
            .O(N__37830),
            .I(\foc.u_Park_Transform.n753 ));
    LocalMux I__5501 (
            .O(N__37827),
            .I(\foc.u_Park_Transform.n753 ));
    CascadeMux I__5500 (
            .O(N__37822),
            .I(N__37819));
    InMux I__5499 (
            .O(N__37819),
            .I(N__37816));
    LocalMux I__5498 (
            .O(N__37816),
            .I(\foc.u_Park_Transform.n703 ));
    InMux I__5497 (
            .O(N__37813),
            .I(N__37810));
    LocalMux I__5496 (
            .O(N__37810),
            .I(N__37807));
    Span4Mux_h I__5495 (
            .O(N__37807),
            .I(N__37804));
    Odrv4 I__5494 (
            .O(N__37804),
            .I(\foc.u_Park_Transform.n754 ));
    InMux I__5493 (
            .O(N__37801),
            .I(\foc.u_Park_Transform.n17021 ));
    InMux I__5492 (
            .O(N__37798),
            .I(\foc.u_Park_Transform.n755 ));
    CascadeMux I__5491 (
            .O(N__37795),
            .I(N__37792));
    InMux I__5490 (
            .O(N__37792),
            .I(N__37789));
    LocalMux I__5489 (
            .O(N__37789),
            .I(N__37786));
    Span4Mux_h I__5488 (
            .O(N__37786),
            .I(N__37783));
    Odrv4 I__5487 (
            .O(N__37783),
            .I(\foc.u_Park_Transform.n755_THRU_CO ));
    InMux I__5486 (
            .O(N__37780),
            .I(\foc.u_Park_Transform.n747 ));
    CascadeMux I__5485 (
            .O(N__37777),
            .I(N__37774));
    InMux I__5484 (
            .O(N__37774),
            .I(N__37771));
    LocalMux I__5483 (
            .O(N__37771),
            .I(N__37768));
    Span4Mux_v I__5482 (
            .O(N__37768),
            .I(N__37765));
    Odrv4 I__5481 (
            .O(N__37765),
            .I(\foc.u_Park_Transform.n747_THRU_CO ));
    CascadeMux I__5480 (
            .O(N__37762),
            .I(N__37746));
    CascadeMux I__5479 (
            .O(N__37761),
            .I(N__37742));
    CascadeMux I__5478 (
            .O(N__37760),
            .I(N__37738));
    CascadeMux I__5477 (
            .O(N__37759),
            .I(N__37733));
    CascadeMux I__5476 (
            .O(N__37758),
            .I(N__37730));
    CascadeMux I__5475 (
            .O(N__37757),
            .I(N__37726));
    CascadeMux I__5474 (
            .O(N__37756),
            .I(N__37722));
    CascadeMux I__5473 (
            .O(N__37755),
            .I(N__37717));
    InMux I__5472 (
            .O(N__37754),
            .I(N__37710));
    CascadeMux I__5471 (
            .O(N__37753),
            .I(N__37707));
    CascadeMux I__5470 (
            .O(N__37752),
            .I(N__37704));
    CascadeMux I__5469 (
            .O(N__37751),
            .I(N__37701));
    CascadeMux I__5468 (
            .O(N__37750),
            .I(N__37697));
    InMux I__5467 (
            .O(N__37749),
            .I(N__37693));
    InMux I__5466 (
            .O(N__37746),
            .I(N__37680));
    InMux I__5465 (
            .O(N__37745),
            .I(N__37680));
    InMux I__5464 (
            .O(N__37742),
            .I(N__37680));
    InMux I__5463 (
            .O(N__37741),
            .I(N__37680));
    InMux I__5462 (
            .O(N__37738),
            .I(N__37680));
    InMux I__5461 (
            .O(N__37737),
            .I(N__37680));
    InMux I__5460 (
            .O(N__37736),
            .I(N__37675));
    InMux I__5459 (
            .O(N__37733),
            .I(N__37675));
    InMux I__5458 (
            .O(N__37730),
            .I(N__37662));
    InMux I__5457 (
            .O(N__37729),
            .I(N__37662));
    InMux I__5456 (
            .O(N__37726),
            .I(N__37662));
    InMux I__5455 (
            .O(N__37725),
            .I(N__37662));
    InMux I__5454 (
            .O(N__37722),
            .I(N__37662));
    InMux I__5453 (
            .O(N__37721),
            .I(N__37662));
    InMux I__5452 (
            .O(N__37720),
            .I(N__37657));
    InMux I__5451 (
            .O(N__37717),
            .I(N__37657));
    CascadeMux I__5450 (
            .O(N__37716),
            .I(N__37654));
    CascadeMux I__5449 (
            .O(N__37715),
            .I(N__37651));
    CascadeMux I__5448 (
            .O(N__37714),
            .I(N__37648));
    CascadeMux I__5447 (
            .O(N__37713),
            .I(N__37644));
    LocalMux I__5446 (
            .O(N__37710),
            .I(N__37640));
    InMux I__5445 (
            .O(N__37707),
            .I(N__37637));
    InMux I__5444 (
            .O(N__37704),
            .I(N__37626));
    InMux I__5443 (
            .O(N__37701),
            .I(N__37626));
    InMux I__5442 (
            .O(N__37700),
            .I(N__37626));
    InMux I__5441 (
            .O(N__37697),
            .I(N__37626));
    InMux I__5440 (
            .O(N__37696),
            .I(N__37626));
    LocalMux I__5439 (
            .O(N__37693),
            .I(N__37623));
    LocalMux I__5438 (
            .O(N__37680),
            .I(N__37618));
    LocalMux I__5437 (
            .O(N__37675),
            .I(N__37618));
    LocalMux I__5436 (
            .O(N__37662),
            .I(N__37613));
    LocalMux I__5435 (
            .O(N__37657),
            .I(N__37613));
    InMux I__5434 (
            .O(N__37654),
            .I(N__37610));
    InMux I__5433 (
            .O(N__37651),
            .I(N__37599));
    InMux I__5432 (
            .O(N__37648),
            .I(N__37599));
    InMux I__5431 (
            .O(N__37647),
            .I(N__37599));
    InMux I__5430 (
            .O(N__37644),
            .I(N__37599));
    InMux I__5429 (
            .O(N__37643),
            .I(N__37599));
    Odrv4 I__5428 (
            .O(N__37640),
            .I(\foc.u_Park_Transform.n604 ));
    LocalMux I__5427 (
            .O(N__37637),
            .I(\foc.u_Park_Transform.n604 ));
    LocalMux I__5426 (
            .O(N__37626),
            .I(\foc.u_Park_Transform.n604 ));
    Odrv4 I__5425 (
            .O(N__37623),
            .I(\foc.u_Park_Transform.n604 ));
    Odrv12 I__5424 (
            .O(N__37618),
            .I(\foc.u_Park_Transform.n604 ));
    Odrv4 I__5423 (
            .O(N__37613),
            .I(\foc.u_Park_Transform.n604 ));
    LocalMux I__5422 (
            .O(N__37610),
            .I(\foc.u_Park_Transform.n604 ));
    LocalMux I__5421 (
            .O(N__37599),
            .I(\foc.u_Park_Transform.n604 ));
    CascadeMux I__5420 (
            .O(N__37582),
            .I(N__37579));
    InMux I__5419 (
            .O(N__37579),
            .I(N__37576));
    LocalMux I__5418 (
            .O(N__37576),
            .I(\foc.u_Park_Transform.n66_adj_2033 ));
    InMux I__5417 (
            .O(N__37573),
            .I(\foc.u_Park_Transform.n17008 ));
    CascadeMux I__5416 (
            .O(N__37570),
            .I(N__37567));
    InMux I__5415 (
            .O(N__37567),
            .I(N__37564));
    LocalMux I__5414 (
            .O(N__37564),
            .I(\foc.u_Park_Transform.n115_adj_2028 ));
    InMux I__5413 (
            .O(N__37561),
            .I(\foc.u_Park_Transform.n17009 ));
    InMux I__5412 (
            .O(N__37558),
            .I(N__37555));
    LocalMux I__5411 (
            .O(N__37555),
            .I(\foc.u_Park_Transform.n164_adj_2014 ));
    InMux I__5410 (
            .O(N__37552),
            .I(\foc.u_Park_Transform.n17010 ));
    CascadeMux I__5409 (
            .O(N__37549),
            .I(N__37546));
    InMux I__5408 (
            .O(N__37546),
            .I(N__37543));
    LocalMux I__5407 (
            .O(N__37543),
            .I(\foc.u_Park_Transform.n213_adj_1999 ));
    InMux I__5406 (
            .O(N__37540),
            .I(\foc.u_Park_Transform.n17011 ));
    InMux I__5405 (
            .O(N__37537),
            .I(N__37534));
    LocalMux I__5404 (
            .O(N__37534),
            .I(\foc.u_Park_Transform.n262 ));
    InMux I__5403 (
            .O(N__37531),
            .I(\foc.u_Park_Transform.n17012 ));
    CascadeMux I__5402 (
            .O(N__37528),
            .I(N__37525));
    InMux I__5401 (
            .O(N__37525),
            .I(N__37522));
    LocalMux I__5400 (
            .O(N__37522),
            .I(\foc.u_Park_Transform.n311_adj_2022 ));
    InMux I__5399 (
            .O(N__37519),
            .I(\foc.u_Park_Transform.n17013 ));
    InMux I__5398 (
            .O(N__37516),
            .I(N__37513));
    LocalMux I__5397 (
            .O(N__37513),
            .I(\foc.u_Park_Transform.n360_adj_2009 ));
    InMux I__5396 (
            .O(N__37510),
            .I(\foc.u_Park_Transform.n17014 ));
    InMux I__5395 (
            .O(N__37507),
            .I(\foc.u_Park_Transform.n17226 ));
    InMux I__5394 (
            .O(N__37504),
            .I(\foc.u_Park_Transform.n17227 ));
    InMux I__5393 (
            .O(N__37501),
            .I(bfn_14_12_0_));
    InMux I__5392 (
            .O(N__37498),
            .I(\foc.u_Park_Transform.n17229 ));
    InMux I__5391 (
            .O(N__37495),
            .I(\foc.u_Park_Transform.n17230 ));
    InMux I__5390 (
            .O(N__37492),
            .I(\foc.u_Park_Transform.n17231 ));
    InMux I__5389 (
            .O(N__37489),
            .I(\foc.u_Park_Transform.n17232 ));
    InMux I__5388 (
            .O(N__37486),
            .I(\foc.u_Park_Transform.n17233 ));
    InMux I__5387 (
            .O(N__37483),
            .I(N__37480));
    LocalMux I__5386 (
            .O(N__37480),
            .I(N__37477));
    Span4Mux_v I__5385 (
            .O(N__37477),
            .I(N__37474));
    Odrv4 I__5384 (
            .O(N__37474),
            .I(\foc.u_Park_Transform.n746 ));
    InMux I__5383 (
            .O(N__37471),
            .I(\foc.u_Park_Transform.n17234 ));
    InMux I__5382 (
            .O(N__37468),
            .I(N__37465));
    LocalMux I__5381 (
            .O(N__37465),
            .I(\foc.dCurrent_29 ));
    InMux I__5380 (
            .O(N__37462),
            .I(N__37459));
    LocalMux I__5379 (
            .O(N__37459),
            .I(\foc.dCurrent_28 ));
    InMux I__5378 (
            .O(N__37456),
            .I(N__37453));
    LocalMux I__5377 (
            .O(N__37453),
            .I(\foc.dCurrent_30 ));
    InMux I__5376 (
            .O(N__37450),
            .I(\foc.u_Park_Transform.n17221 ));
    InMux I__5375 (
            .O(N__37447),
            .I(\foc.u_Park_Transform.n17222 ));
    InMux I__5374 (
            .O(N__37444),
            .I(\foc.u_Park_Transform.n17223 ));
    InMux I__5373 (
            .O(N__37441),
            .I(\foc.u_Park_Transform.n17224 ));
    InMux I__5372 (
            .O(N__37438),
            .I(\foc.u_Park_Transform.n17225 ));
    InMux I__5371 (
            .O(N__37435),
            .I(N__37432));
    LocalMux I__5370 (
            .O(N__37432),
            .I(\foc.u_Park_Transform.Product1_mul_temp_23 ));
    InMux I__5369 (
            .O(N__37429),
            .I(N__37426));
    LocalMux I__5368 (
            .O(N__37426),
            .I(N__37423));
    Odrv12 I__5367 (
            .O(N__37423),
            .I(\foc.dCurrent_25 ));
    InMux I__5366 (
            .O(N__37420),
            .I(\foc.u_Park_Transform.n17297 ));
    InMux I__5365 (
            .O(N__37417),
            .I(N__37414));
    LocalMux I__5364 (
            .O(N__37414),
            .I(\foc.u_Park_Transform.Product1_mul_temp_24 ));
    InMux I__5363 (
            .O(N__37411),
            .I(\foc.u_Park_Transform.n17298 ));
    InMux I__5362 (
            .O(N__37408),
            .I(N__37405));
    LocalMux I__5361 (
            .O(N__37405),
            .I(\foc.u_Park_Transform.Product1_mul_temp_25 ));
    InMux I__5360 (
            .O(N__37402),
            .I(\foc.u_Park_Transform.n17299 ));
    InMux I__5359 (
            .O(N__37399),
            .I(N__37396));
    LocalMux I__5358 (
            .O(N__37396),
            .I(\foc.u_Park_Transform.Product1_mul_temp_26 ));
    InMux I__5357 (
            .O(N__37393),
            .I(bfn_14_10_0_));
    InMux I__5356 (
            .O(N__37390),
            .I(N__37387));
    LocalMux I__5355 (
            .O(N__37387),
            .I(\foc.u_Park_Transform.Product1_mul_temp_27 ));
    InMux I__5354 (
            .O(N__37384),
            .I(\foc.u_Park_Transform.n17301 ));
    InMux I__5353 (
            .O(N__37381),
            .I(N__37378));
    LocalMux I__5352 (
            .O(N__37378),
            .I(\foc.u_Park_Transform.Product1_mul_temp_28 ));
    InMux I__5351 (
            .O(N__37375),
            .I(\foc.u_Park_Transform.n17302 ));
    InMux I__5350 (
            .O(N__37372),
            .I(N__37369));
    LocalMux I__5349 (
            .O(N__37369),
            .I(\foc.u_Park_Transform.Product1_mul_temp_29 ));
    InMux I__5348 (
            .O(N__37366),
            .I(\foc.u_Park_Transform.n17303 ));
    CascadeMux I__5347 (
            .O(N__37363),
            .I(\foc.dCurrent_31_cascade_ ));
    InMux I__5346 (
            .O(N__37360),
            .I(N__37357));
    LocalMux I__5345 (
            .O(N__37357),
            .I(\foc.u_Park_Transform.Product1_mul_temp_15 ));
    InMux I__5344 (
            .O(N__37354),
            .I(N__37351));
    LocalMux I__5343 (
            .O(N__37351),
            .I(N__37348));
    Odrv4 I__5342 (
            .O(N__37348),
            .I(\foc.dCurrent_17 ));
    InMux I__5341 (
            .O(N__37345),
            .I(\foc.u_Park_Transform.n17289 ));
    InMux I__5340 (
            .O(N__37342),
            .I(N__37339));
    LocalMux I__5339 (
            .O(N__37339),
            .I(\foc.u_Park_Transform.Product1_mul_temp_16 ));
    InMux I__5338 (
            .O(N__37336),
            .I(N__37333));
    LocalMux I__5337 (
            .O(N__37333),
            .I(N__37330));
    Odrv12 I__5336 (
            .O(N__37330),
            .I(\foc.dCurrent_18 ));
    InMux I__5335 (
            .O(N__37327),
            .I(\foc.u_Park_Transform.n17290 ));
    InMux I__5334 (
            .O(N__37324),
            .I(N__37321));
    LocalMux I__5333 (
            .O(N__37321),
            .I(\foc.u_Park_Transform.Product1_mul_temp_17 ));
    InMux I__5332 (
            .O(N__37318),
            .I(N__37315));
    LocalMux I__5331 (
            .O(N__37315),
            .I(N__37312));
    Odrv4 I__5330 (
            .O(N__37312),
            .I(\foc.dCurrent_19 ));
    InMux I__5329 (
            .O(N__37309),
            .I(\foc.u_Park_Transform.n17291 ));
    InMux I__5328 (
            .O(N__37306),
            .I(N__37303));
    LocalMux I__5327 (
            .O(N__37303),
            .I(\foc.u_Park_Transform.Product1_mul_temp_18 ));
    InMux I__5326 (
            .O(N__37300),
            .I(N__37297));
    LocalMux I__5325 (
            .O(N__37297),
            .I(N__37294));
    Odrv4 I__5324 (
            .O(N__37294),
            .I(\foc.dCurrent_20 ));
    InMux I__5323 (
            .O(N__37291),
            .I(bfn_14_9_0_));
    InMux I__5322 (
            .O(N__37288),
            .I(N__37285));
    LocalMux I__5321 (
            .O(N__37285),
            .I(\foc.u_Park_Transform.Product1_mul_temp_19 ));
    InMux I__5320 (
            .O(N__37282),
            .I(N__37279));
    LocalMux I__5319 (
            .O(N__37279),
            .I(N__37276));
    Odrv4 I__5318 (
            .O(N__37276),
            .I(\foc.dCurrent_21 ));
    InMux I__5317 (
            .O(N__37273),
            .I(\foc.u_Park_Transform.n17293 ));
    InMux I__5316 (
            .O(N__37270),
            .I(N__37267));
    LocalMux I__5315 (
            .O(N__37267),
            .I(\foc.u_Park_Transform.Product1_mul_temp_20 ));
    InMux I__5314 (
            .O(N__37264),
            .I(N__37261));
    LocalMux I__5313 (
            .O(N__37261),
            .I(N__37258));
    Odrv4 I__5312 (
            .O(N__37258),
            .I(\foc.dCurrent_22 ));
    InMux I__5311 (
            .O(N__37255),
            .I(\foc.u_Park_Transform.n17294 ));
    InMux I__5310 (
            .O(N__37252),
            .I(N__37249));
    LocalMux I__5309 (
            .O(N__37249),
            .I(\foc.u_Park_Transform.Product1_mul_temp_21 ));
    InMux I__5308 (
            .O(N__37246),
            .I(N__37243));
    LocalMux I__5307 (
            .O(N__37243),
            .I(N__37240));
    Odrv4 I__5306 (
            .O(N__37240),
            .I(\foc.dCurrent_23 ));
    InMux I__5305 (
            .O(N__37237),
            .I(\foc.u_Park_Transform.n17295 ));
    InMux I__5304 (
            .O(N__37234),
            .I(N__37231));
    LocalMux I__5303 (
            .O(N__37231),
            .I(\foc.u_Park_Transform.Product1_mul_temp_22 ));
    InMux I__5302 (
            .O(N__37228),
            .I(N__37225));
    LocalMux I__5301 (
            .O(N__37225),
            .I(N__37222));
    Odrv4 I__5300 (
            .O(N__37222),
            .I(\foc.dCurrent_24 ));
    InMux I__5299 (
            .O(N__37219),
            .I(\foc.u_Park_Transform.n17296 ));
    InMux I__5298 (
            .O(N__37216),
            .I(N__37213));
    LocalMux I__5297 (
            .O(N__37213),
            .I(\foc.dCurrent_9 ));
    InMux I__5296 (
            .O(N__37210),
            .I(\foc.u_Park_Transform.n17281 ));
    InMux I__5295 (
            .O(N__37207),
            .I(N__37204));
    LocalMux I__5294 (
            .O(N__37204),
            .I(\foc.dCurrent_10 ));
    InMux I__5293 (
            .O(N__37201),
            .I(\foc.u_Park_Transform.n17282 ));
    InMux I__5292 (
            .O(N__37198),
            .I(N__37195));
    LocalMux I__5291 (
            .O(N__37195),
            .I(\foc.dCurrent_11 ));
    InMux I__5290 (
            .O(N__37192),
            .I(\foc.u_Park_Transform.n17283 ));
    InMux I__5289 (
            .O(N__37189),
            .I(N__37186));
    LocalMux I__5288 (
            .O(N__37186),
            .I(N__37183));
    Odrv12 I__5287 (
            .O(N__37183),
            .I(\foc.dCurrent_12 ));
    InMux I__5286 (
            .O(N__37180),
            .I(bfn_14_8_0_));
    InMux I__5285 (
            .O(N__37177),
            .I(N__37174));
    LocalMux I__5284 (
            .O(N__37174),
            .I(N__37171));
    Odrv4 I__5283 (
            .O(N__37171),
            .I(\foc.dCurrent_13 ));
    InMux I__5282 (
            .O(N__37168),
            .I(\foc.u_Park_Transform.n17285 ));
    InMux I__5281 (
            .O(N__37165),
            .I(N__37162));
    LocalMux I__5280 (
            .O(N__37162),
            .I(N__37159));
    Odrv12 I__5279 (
            .O(N__37159),
            .I(\foc.dCurrent_14 ));
    InMux I__5278 (
            .O(N__37156),
            .I(\foc.u_Park_Transform.n17286 ));
    InMux I__5277 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__5276 (
            .O(N__37150),
            .I(N__37147));
    Odrv12 I__5275 (
            .O(N__37147),
            .I(\foc.dCurrent_15 ));
    InMux I__5274 (
            .O(N__37144),
            .I(\foc.u_Park_Transform.n17287 ));
    InMux I__5273 (
            .O(N__37141),
            .I(N__37138));
    LocalMux I__5272 (
            .O(N__37138),
            .I(N__37135));
    Odrv4 I__5271 (
            .O(N__37135),
            .I(\foc.dCurrent_16 ));
    InMux I__5270 (
            .O(N__37132),
            .I(\foc.u_Park_Transform.n17288 ));
    InMux I__5269 (
            .O(N__37129),
            .I(N__37126));
    LocalMux I__5268 (
            .O(N__37126),
            .I(N__37123));
    Odrv4 I__5267 (
            .O(N__37123),
            .I(\foc.dCurrent_4 ));
    InMux I__5266 (
            .O(N__37120),
            .I(N__37117));
    LocalMux I__5265 (
            .O(N__37117),
            .I(N__37114));
    Odrv4 I__5264 (
            .O(N__37114),
            .I(\foc.dCurrent_5 ));
    InMux I__5263 (
            .O(N__37111),
            .I(\foc.u_Park_Transform.n17277 ));
    InMux I__5262 (
            .O(N__37108),
            .I(N__37105));
    LocalMux I__5261 (
            .O(N__37105),
            .I(N__37102));
    Odrv4 I__5260 (
            .O(N__37102),
            .I(\foc.dCurrent_6 ));
    InMux I__5259 (
            .O(N__37099),
            .I(\foc.u_Park_Transform.n17278 ));
    InMux I__5258 (
            .O(N__37096),
            .I(N__37093));
    LocalMux I__5257 (
            .O(N__37093),
            .I(N__37090));
    Odrv4 I__5256 (
            .O(N__37090),
            .I(\foc.dCurrent_7 ));
    InMux I__5255 (
            .O(N__37087),
            .I(\foc.u_Park_Transform.n17279 ));
    InMux I__5254 (
            .O(N__37084),
            .I(N__37081));
    LocalMux I__5253 (
            .O(N__37081),
            .I(N__37078));
    Odrv4 I__5252 (
            .O(N__37078),
            .I(\foc.dCurrent_8 ));
    InMux I__5251 (
            .O(N__37075),
            .I(\foc.u_Park_Transform.n17280 ));
    CascadeMux I__5250 (
            .O(N__37072),
            .I(N__37069));
    InMux I__5249 (
            .O(N__37069),
            .I(N__37066));
    LocalMux I__5248 (
            .O(N__37066),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604 ));
    InMux I__5247 (
            .O(N__37063),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18100 ));
    InMux I__5246 (
            .O(N__37060),
            .I(N__37057));
    LocalMux I__5245 (
            .O(N__37057),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603 ));
    InMux I__5244 (
            .O(N__37054),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18101 ));
    CascadeMux I__5243 (
            .O(N__37051),
            .I(N__37048));
    InMux I__5242 (
            .O(N__37048),
            .I(N__37045));
    LocalMux I__5241 (
            .O(N__37045),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602 ));
    InMux I__5240 (
            .O(N__37042),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18102 ));
    InMux I__5239 (
            .O(N__37039),
            .I(N__37036));
    LocalMux I__5238 (
            .O(N__37036),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601 ));
    InMux I__5237 (
            .O(N__37033),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18103 ));
    CascadeMux I__5236 (
            .O(N__37030),
            .I(N__37027));
    InMux I__5235 (
            .O(N__37027),
            .I(N__37024));
    LocalMux I__5234 (
            .O(N__37024),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600 ));
    InMux I__5233 (
            .O(N__37021),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18104 ));
    CascadeMux I__5232 (
            .O(N__37018),
            .I(N__37015));
    InMux I__5231 (
            .O(N__37015),
            .I(N__37012));
    LocalMux I__5230 (
            .O(N__37012),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599 ));
    InMux I__5229 (
            .O(N__37009),
            .I(N__37006));
    LocalMux I__5228 (
            .O(N__37006),
            .I(N__37003));
    Odrv12 I__5227 (
            .O(N__37003),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619 ));
    InMux I__5226 (
            .O(N__37000),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18105 ));
    InMux I__5225 (
            .O(N__36997),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620 ));
    InMux I__5224 (
            .O(N__36994),
            .I(N__36991));
    LocalMux I__5223 (
            .O(N__36991),
            .I(N__36988));
    Odrv12 I__5222 (
            .O(N__36988),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO ));
    InMux I__5221 (
            .O(N__36985),
            .I(N__36982));
    LocalMux I__5220 (
            .O(N__36982),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618 ));
    InMux I__5219 (
            .O(N__36979),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18092 ));
    InMux I__5218 (
            .O(N__36976),
            .I(N__36973));
    LocalMux I__5217 (
            .O(N__36973),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616 ));
    InMux I__5216 (
            .O(N__36970),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18093 ));
    InMux I__5215 (
            .O(N__36967),
            .I(N__36964));
    LocalMux I__5214 (
            .O(N__36964),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614 ));
    InMux I__5213 (
            .O(N__36961),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18094 ));
    InMux I__5212 (
            .O(N__36958),
            .I(N__36955));
    LocalMux I__5211 (
            .O(N__36955),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612 ));
    InMux I__5210 (
            .O(N__36952),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18095 ));
    InMux I__5209 (
            .O(N__36949),
            .I(N__36946));
    LocalMux I__5208 (
            .O(N__36946),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610 ));
    InMux I__5207 (
            .O(N__36943),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18096 ));
    InMux I__5206 (
            .O(N__36940),
            .I(N__36937));
    LocalMux I__5205 (
            .O(N__36937),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608 ));
    InMux I__5204 (
            .O(N__36934),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18097 ));
    InMux I__5203 (
            .O(N__36931),
            .I(N__36928));
    LocalMux I__5202 (
            .O(N__36928),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606 ));
    InMux I__5201 (
            .O(N__36925),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18098 ));
    InMux I__5200 (
            .O(N__36922),
            .I(N__36919));
    LocalMux I__5199 (
            .O(N__36919),
            .I(N__36916));
    Odrv4 I__5198 (
            .O(N__36916),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605 ));
    InMux I__5197 (
            .O(N__36913),
            .I(bfn_13_26_0_));
    CascadeMux I__5196 (
            .O(N__36910),
            .I(N__36907));
    InMux I__5195 (
            .O(N__36907),
            .I(N__36904));
    LocalMux I__5194 (
            .O(N__36904),
            .I(N__36901));
    Odrv4 I__5193 (
            .O(N__36901),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597 ));
    InMux I__5192 (
            .O(N__36898),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17965 ));
    InMux I__5191 (
            .O(N__36895),
            .I(N__36892));
    LocalMux I__5190 (
            .O(N__36892),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n774 ));
    CascadeMux I__5189 (
            .O(N__36889),
            .I(N__36886));
    InMux I__5188 (
            .O(N__36886),
            .I(N__36883));
    LocalMux I__5187 (
            .O(N__36883),
            .I(N__36880));
    Odrv4 I__5186 (
            .O(N__36880),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO ));
    InMux I__5185 (
            .O(N__36877),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17966 ));
    InMux I__5184 (
            .O(N__36874),
            .I(N__36871));
    LocalMux I__5183 (
            .O(N__36871),
            .I(N__36868));
    Odrv12 I__5182 (
            .O(N__36868),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737 ));
    CascadeMux I__5181 (
            .O(N__36865),
            .I(N__36862));
    InMux I__5180 (
            .O(N__36862),
            .I(N__36859));
    LocalMux I__5179 (
            .O(N__36859),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO ));
    InMux I__5178 (
            .O(N__36856),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17967 ));
    CascadeMux I__5177 (
            .O(N__36853),
            .I(N__36850));
    InMux I__5176 (
            .O(N__36850),
            .I(N__36847));
    LocalMux I__5175 (
            .O(N__36847),
            .I(N__36844));
    Odrv12 I__5174 (
            .O(N__36844),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO ));
    InMux I__5173 (
            .O(N__36841),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17968 ));
    InMux I__5172 (
            .O(N__36838),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17969 ));
    InMux I__5171 (
            .O(N__36835),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17970 ));
    InMux I__5170 (
            .O(N__36832),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17971 ));
    InMux I__5169 (
            .O(N__36829),
            .I(bfn_13_24_0_));
    InMux I__5168 (
            .O(N__36826),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17957 ));
    InMux I__5167 (
            .O(N__36823),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17958 ));
    InMux I__5166 (
            .O(N__36820),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17959 ));
    InMux I__5165 (
            .O(N__36817),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17960 ));
    InMux I__5164 (
            .O(N__36814),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17961 ));
    InMux I__5163 (
            .O(N__36811),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17962 ));
    InMux I__5162 (
            .O(N__36808),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17963 ));
    InMux I__5161 (
            .O(N__36805),
            .I(bfn_13_23_0_));
    CascadeMux I__5160 (
            .O(N__36802),
            .I(N__36799));
    InMux I__5159 (
            .O(N__36799),
            .I(N__36796));
    LocalMux I__5158 (
            .O(N__36796),
            .I(N__36793));
    Odrv4 I__5157 (
            .O(N__36793),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742 ));
    InMux I__5156 (
            .O(N__36790),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17858 ));
    InMux I__5155 (
            .O(N__36787),
            .I(N__36784));
    LocalMux I__5154 (
            .O(N__36784),
            .I(N__36781));
    Span4Mux_h I__5153 (
            .O(N__36781),
            .I(N__36778));
    Odrv4 I__5152 (
            .O(N__36778),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741 ));
    InMux I__5151 (
            .O(N__36775),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17859 ));
    InMux I__5150 (
            .O(N__36772),
            .I(N__36769));
    LocalMux I__5149 (
            .O(N__36769),
            .I(N__36766));
    Odrv4 I__5148 (
            .O(N__36766),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n326 ));
    InMux I__5147 (
            .O(N__36763),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17860 ));
    InMux I__5146 (
            .O(N__36760),
            .I(N__36757));
    LocalMux I__5145 (
            .O(N__36757),
            .I(N__36754));
    Span4Mux_h I__5144 (
            .O(N__36754),
            .I(N__36751));
    Odrv4 I__5143 (
            .O(N__36751),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n375 ));
    InMux I__5142 (
            .O(N__36748),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17861 ));
    InMux I__5141 (
            .O(N__36745),
            .I(N__36742));
    LocalMux I__5140 (
            .O(N__36742),
            .I(N__36739));
    Odrv4 I__5139 (
            .O(N__36739),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n424 ));
    InMux I__5138 (
            .O(N__36736),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17862 ));
    InMux I__5137 (
            .O(N__36733),
            .I(N__36730));
    LocalMux I__5136 (
            .O(N__36730),
            .I(N__36727));
    Odrv4 I__5135 (
            .O(N__36727),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n473 ));
    InMux I__5134 (
            .O(N__36724),
            .I(bfn_13_21_0_));
    CascadeMux I__5133 (
            .O(N__36721),
            .I(N__36717));
    CascadeMux I__5132 (
            .O(N__36720),
            .I(N__36713));
    InMux I__5131 (
            .O(N__36717),
            .I(N__36706));
    InMux I__5130 (
            .O(N__36716),
            .I(N__36706));
    InMux I__5129 (
            .O(N__36713),
            .I(N__36706));
    LocalMux I__5128 (
            .O(N__36706),
            .I(N__36703));
    Odrv4 I__5127 (
            .O(N__36703),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n522 ));
    InMux I__5126 (
            .O(N__36700),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17864 ));
    InMux I__5125 (
            .O(N__36697),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17865 ));
    InMux I__5124 (
            .O(N__36694),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736 ));
    InMux I__5123 (
            .O(N__36691),
            .I(N__36688));
    LocalMux I__5122 (
            .O(N__36688),
            .I(N__36685));
    Odrv4 I__5121 (
            .O(N__36685),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014 ));
    CascadeMux I__5120 (
            .O(N__36682),
            .I(N__36675));
    CascadeMux I__5119 (
            .O(N__36681),
            .I(N__36672));
    CascadeMux I__5118 (
            .O(N__36680),
            .I(N__36669));
    CascadeMux I__5117 (
            .O(N__36679),
            .I(N__36666));
    CascadeMux I__5116 (
            .O(N__36678),
            .I(N__36662));
    InMux I__5115 (
            .O(N__36675),
            .I(N__36655));
    InMux I__5114 (
            .O(N__36672),
            .I(N__36655));
    InMux I__5113 (
            .O(N__36669),
            .I(N__36644));
    InMux I__5112 (
            .O(N__36666),
            .I(N__36644));
    InMux I__5111 (
            .O(N__36665),
            .I(N__36644));
    InMux I__5110 (
            .O(N__36662),
            .I(N__36644));
    InMux I__5109 (
            .O(N__36661),
            .I(N__36644));
    InMux I__5108 (
            .O(N__36660),
            .I(N__36641));
    LocalMux I__5107 (
            .O(N__36655),
            .I(N__36636));
    LocalMux I__5106 (
            .O(N__36644),
            .I(N__36636));
    LocalMux I__5105 (
            .O(N__36641),
            .I(N__36633));
    Span4Mux_h I__5104 (
            .O(N__36636),
            .I(N__36630));
    Span4Mux_v I__5103 (
            .O(N__36633),
            .I(N__36627));
    Odrv4 I__5102 (
            .O(N__36630),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810 ));
    Odrv4 I__5101 (
            .O(N__36627),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810 ));
    InMux I__5100 (
            .O(N__36622),
            .I(N__36619));
    LocalMux I__5099 (
            .O(N__36619),
            .I(N__36616));
    Span4Mux_h I__5098 (
            .O(N__36616),
            .I(N__36613));
    Odrv4 I__5097 (
            .O(N__36613),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111 ));
    InMux I__5096 (
            .O(N__36610),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373 ));
    InMux I__5095 (
            .O(N__36607),
            .I(N__36604));
    LocalMux I__5094 (
            .O(N__36604),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114 ));
    InMux I__5093 (
            .O(N__36601),
            .I(N__36598));
    LocalMux I__5092 (
            .O(N__36598),
            .I(N__36595));
    Span4Mux_h I__5091 (
            .O(N__36595),
            .I(N__36592));
    Odrv4 I__5090 (
            .O(N__36592),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215 ));
    InMux I__5089 (
            .O(N__36589),
            .I(bfn_13_18_0_));
    InMux I__5088 (
            .O(N__36586),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216 ));
    CascadeMux I__5087 (
            .O(N__36583),
            .I(N__36580));
    InMux I__5086 (
            .O(N__36580),
            .I(N__36577));
    LocalMux I__5085 (
            .O(N__36577),
            .I(N__36574));
    Span4Mux_h I__5084 (
            .O(N__36574),
            .I(N__36571));
    Odrv4 I__5083 (
            .O(N__36571),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO ));
    InMux I__5082 (
            .O(N__36568),
            .I(N__36562));
    InMux I__5081 (
            .O(N__36567),
            .I(N__36562));
    LocalMux I__5080 (
            .O(N__36562),
            .I(N__36558));
    InMux I__5079 (
            .O(N__36561),
            .I(N__36555));
    Span4Mux_v I__5078 (
            .O(N__36558),
            .I(N__36550));
    LocalMux I__5077 (
            .O(N__36555),
            .I(N__36550));
    Span4Mux_v I__5076 (
            .O(N__36550),
            .I(N__36547));
    Odrv4 I__5075 (
            .O(N__36547),
            .I(\foc.Look_Up_Table_out1_1_0 ));
    InMux I__5074 (
            .O(N__36544),
            .I(N__36541));
    LocalMux I__5073 (
            .O(N__36541),
            .I(N__36538));
    Span12Mux_v I__5072 (
            .O(N__36538),
            .I(N__36534));
    InMux I__5071 (
            .O(N__36537),
            .I(N__36531));
    Odrv12 I__5070 (
            .O(N__36534),
            .I(n794));
    LocalMux I__5069 (
            .O(N__36531),
            .I(n794));
    InMux I__5068 (
            .O(N__36526),
            .I(N__36523));
    LocalMux I__5067 (
            .O(N__36523),
            .I(N__36520));
    Odrv4 I__5066 (
            .O(N__36520),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750 ));
    CascadeMux I__5065 (
            .O(N__36517),
            .I(N__36514));
    InMux I__5064 (
            .O(N__36514),
            .I(N__36511));
    LocalMux I__5063 (
            .O(N__36511),
            .I(N__36508));
    Odrv4 I__5062 (
            .O(N__36508),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748 ));
    InMux I__5061 (
            .O(N__36505),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17856 ));
    InMux I__5060 (
            .O(N__36502),
            .I(N__36499));
    LocalMux I__5059 (
            .O(N__36499),
            .I(N__36496));
    Odrv4 I__5058 (
            .O(N__36496),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746 ));
    InMux I__5057 (
            .O(N__36493),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17857 ));
    InMux I__5056 (
            .O(N__36490),
            .I(\foc.u_Park_Transform.n763_adj_2054 ));
    CascadeMux I__5055 (
            .O(N__36487),
            .I(N__36484));
    InMux I__5054 (
            .O(N__36484),
            .I(N__36481));
    LocalMux I__5053 (
            .O(N__36481),
            .I(N__36478));
    Span4Mux_v I__5052 (
            .O(N__36478),
            .I(N__36475));
    Odrv4 I__5051 (
            .O(N__36475),
            .I(\foc.u_Park_Transform.n763_adj_2054_THRU_CO ));
    InMux I__5050 (
            .O(N__36472),
            .I(N__36464));
    CascadeMux I__5049 (
            .O(N__36471),
            .I(N__36461));
    CascadeMux I__5048 (
            .O(N__36470),
            .I(N__36458));
    CascadeMux I__5047 (
            .O(N__36469),
            .I(N__36455));
    CascadeMux I__5046 (
            .O(N__36468),
            .I(N__36452));
    CascadeMux I__5045 (
            .O(N__36467),
            .I(N__36448));
    LocalMux I__5044 (
            .O(N__36464),
            .I(N__36444));
    InMux I__5043 (
            .O(N__36461),
            .I(N__36439));
    InMux I__5042 (
            .O(N__36458),
            .I(N__36439));
    InMux I__5041 (
            .O(N__36455),
            .I(N__36428));
    InMux I__5040 (
            .O(N__36452),
            .I(N__36428));
    InMux I__5039 (
            .O(N__36451),
            .I(N__36428));
    InMux I__5038 (
            .O(N__36448),
            .I(N__36428));
    InMux I__5037 (
            .O(N__36447),
            .I(N__36428));
    Span4Mux_v I__5036 (
            .O(N__36444),
            .I(N__36425));
    LocalMux I__5035 (
            .O(N__36439),
            .I(N__36420));
    LocalMux I__5034 (
            .O(N__36428),
            .I(N__36420));
    Odrv4 I__5033 (
            .O(N__36425),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813 ));
    Odrv12 I__5032 (
            .O(N__36420),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813 ));
    CascadeMux I__5031 (
            .O(N__36415),
            .I(N__36412));
    InMux I__5030 (
            .O(N__36412),
            .I(N__36409));
    LocalMux I__5029 (
            .O(N__36409),
            .I(N__36406));
    Span4Mux_v I__5028 (
            .O(N__36406),
            .I(N__36403));
    Odrv4 I__5027 (
            .O(N__36403),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411 ));
    CascadeMux I__5026 (
            .O(N__36400),
            .I(N__36397));
    InMux I__5025 (
            .O(N__36397),
            .I(N__36394));
    LocalMux I__5024 (
            .O(N__36394),
            .I(N__36391));
    Odrv4 I__5023 (
            .O(N__36391),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414 ));
    InMux I__5022 (
            .O(N__36388),
            .I(N__36385));
    LocalMux I__5021 (
            .O(N__36385),
            .I(N__36382));
    Odrv12 I__5020 (
            .O(N__36382),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511 ));
    InMux I__5019 (
            .O(N__36379),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367 ));
    InMux I__5018 (
            .O(N__36376),
            .I(N__36373));
    LocalMux I__5017 (
            .O(N__36373),
            .I(N__36370));
    Span4Mux_h I__5016 (
            .O(N__36370),
            .I(N__36367));
    Odrv4 I__5015 (
            .O(N__36367),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514 ));
    CascadeMux I__5014 (
            .O(N__36364),
            .I(N__36361));
    InMux I__5013 (
            .O(N__36361),
            .I(N__36358));
    LocalMux I__5012 (
            .O(N__36358),
            .I(N__36355));
    Span4Mux_h I__5011 (
            .O(N__36355),
            .I(N__36352));
    Odrv4 I__5010 (
            .O(N__36352),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611 ));
    InMux I__5009 (
            .O(N__36349),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368 ));
    CascadeMux I__5008 (
            .O(N__36346),
            .I(N__36343));
    InMux I__5007 (
            .O(N__36343),
            .I(N__36340));
    LocalMux I__5006 (
            .O(N__36340),
            .I(N__36337));
    Odrv4 I__5005 (
            .O(N__36337),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614 ));
    InMux I__5004 (
            .O(N__36334),
            .I(N__36331));
    LocalMux I__5003 (
            .O(N__36331),
            .I(N__36328));
    Span4Mux_h I__5002 (
            .O(N__36328),
            .I(N__36325));
    Odrv4 I__5001 (
            .O(N__36325),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711 ));
    InMux I__5000 (
            .O(N__36322),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369 ));
    InMux I__4999 (
            .O(N__36319),
            .I(N__36316));
    LocalMux I__4998 (
            .O(N__36316),
            .I(N__36313));
    Odrv4 I__4997 (
            .O(N__36313),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714 ));
    CascadeMux I__4996 (
            .O(N__36310),
            .I(N__36307));
    InMux I__4995 (
            .O(N__36307),
            .I(N__36304));
    LocalMux I__4994 (
            .O(N__36304),
            .I(N__36301));
    Odrv12 I__4993 (
            .O(N__36301),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811 ));
    InMux I__4992 (
            .O(N__36298),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370 ));
    InMux I__4991 (
            .O(N__36295),
            .I(N__36292));
    LocalMux I__4990 (
            .O(N__36292),
            .I(N__36289));
    Odrv4 I__4989 (
            .O(N__36289),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814 ));
    InMux I__4988 (
            .O(N__36286),
            .I(N__36283));
    LocalMux I__4987 (
            .O(N__36283),
            .I(N__36280));
    Odrv4 I__4986 (
            .O(N__36280),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911 ));
    InMux I__4985 (
            .O(N__36277),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371 ));
    InMux I__4984 (
            .O(N__36274),
            .I(N__36271));
    LocalMux I__4983 (
            .O(N__36271),
            .I(N__36268));
    Odrv4 I__4982 (
            .O(N__36268),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914 ));
    CascadeMux I__4981 (
            .O(N__36265),
            .I(N__36262));
    InMux I__4980 (
            .O(N__36262),
            .I(N__36259));
    LocalMux I__4979 (
            .O(N__36259),
            .I(N__36256));
    Odrv12 I__4978 (
            .O(N__36256),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011 ));
    InMux I__4977 (
            .O(N__36253),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372 ));
    CascadeMux I__4976 (
            .O(N__36250),
            .I(N__36247));
    InMux I__4975 (
            .O(N__36247),
            .I(N__36244));
    LocalMux I__4974 (
            .O(N__36244),
            .I(\foc.u_Park_Transform.n412_adj_1995 ));
    InMux I__4973 (
            .O(N__36241),
            .I(\foc.u_Park_Transform.n16984 ));
    CascadeMux I__4972 (
            .O(N__36238),
            .I(N__36235));
    InMux I__4971 (
            .O(N__36235),
            .I(N__36232));
    LocalMux I__4970 (
            .O(N__36232),
            .I(\foc.u_Park_Transform.n415 ));
    InMux I__4969 (
            .O(N__36229),
            .I(N__36226));
    LocalMux I__4968 (
            .O(N__36226),
            .I(N__36223));
    Odrv4 I__4967 (
            .O(N__36223),
            .I(\foc.u_Park_Transform.n461_adj_2007 ));
    InMux I__4966 (
            .O(N__36220),
            .I(bfn_13_16_0_));
    InMux I__4965 (
            .O(N__36217),
            .I(N__36214));
    LocalMux I__4964 (
            .O(N__36214),
            .I(\foc.u_Park_Transform.n464 ));
    CascadeMux I__4963 (
            .O(N__36211),
            .I(N__36208));
    InMux I__4962 (
            .O(N__36208),
            .I(N__36205));
    LocalMux I__4961 (
            .O(N__36205),
            .I(N__36202));
    Odrv4 I__4960 (
            .O(N__36202),
            .I(\foc.u_Park_Transform.n510 ));
    InMux I__4959 (
            .O(N__36199),
            .I(\foc.u_Park_Transform.n16986 ));
    CascadeMux I__4958 (
            .O(N__36196),
            .I(N__36193));
    InMux I__4957 (
            .O(N__36193),
            .I(N__36190));
    LocalMux I__4956 (
            .O(N__36190),
            .I(\foc.u_Park_Transform.n513 ));
    InMux I__4955 (
            .O(N__36187),
            .I(N__36184));
    LocalMux I__4954 (
            .O(N__36184),
            .I(N__36181));
    Odrv4 I__4953 (
            .O(N__36181),
            .I(\foc.u_Park_Transform.n559 ));
    InMux I__4952 (
            .O(N__36178),
            .I(\foc.u_Park_Transform.n16987 ));
    InMux I__4951 (
            .O(N__36175),
            .I(N__36172));
    LocalMux I__4950 (
            .O(N__36172),
            .I(\foc.u_Park_Transform.n562 ));
    InMux I__4949 (
            .O(N__36169),
            .I(N__36166));
    LocalMux I__4948 (
            .O(N__36166),
            .I(N__36163));
    Odrv4 I__4947 (
            .O(N__36163),
            .I(\foc.u_Park_Transform.n608_adj_2067 ));
    InMux I__4946 (
            .O(N__36160),
            .I(\foc.u_Park_Transform.n16988 ));
    InMux I__4945 (
            .O(N__36157),
            .I(N__36154));
    LocalMux I__4944 (
            .O(N__36154),
            .I(\foc.u_Park_Transform.n611_adj_2107 ));
    InMux I__4943 (
            .O(N__36151),
            .I(N__36148));
    LocalMux I__4942 (
            .O(N__36148),
            .I(N__36145));
    Odrv4 I__4941 (
            .O(N__36145),
            .I(\foc.u_Park_Transform.n657_adj_2064 ));
    InMux I__4940 (
            .O(N__36142),
            .I(\foc.u_Park_Transform.n16989 ));
    InMux I__4939 (
            .O(N__36139),
            .I(N__36136));
    LocalMux I__4938 (
            .O(N__36136),
            .I(\foc.u_Park_Transform.n660_adj_2091 ));
    CascadeMux I__4937 (
            .O(N__36133),
            .I(N__36121));
    CascadeMux I__4936 (
            .O(N__36132),
            .I(N__36118));
    CascadeMux I__4935 (
            .O(N__36131),
            .I(N__36115));
    CascadeMux I__4934 (
            .O(N__36130),
            .I(N__36112));
    CascadeMux I__4933 (
            .O(N__36129),
            .I(N__36108));
    CascadeMux I__4932 (
            .O(N__36128),
            .I(N__36104));
    CascadeMux I__4931 (
            .O(N__36127),
            .I(N__36100));
    CascadeMux I__4930 (
            .O(N__36126),
            .I(N__36096));
    CascadeMux I__4929 (
            .O(N__36125),
            .I(N__36092));
    InMux I__4928 (
            .O(N__36124),
            .I(N__36086));
    InMux I__4927 (
            .O(N__36121),
            .I(N__36086));
    InMux I__4926 (
            .O(N__36118),
            .I(N__36075));
    InMux I__4925 (
            .O(N__36115),
            .I(N__36064));
    InMux I__4924 (
            .O(N__36112),
            .I(N__36064));
    InMux I__4923 (
            .O(N__36111),
            .I(N__36064));
    InMux I__4922 (
            .O(N__36108),
            .I(N__36064));
    InMux I__4921 (
            .O(N__36107),
            .I(N__36064));
    InMux I__4920 (
            .O(N__36104),
            .I(N__36047));
    InMux I__4919 (
            .O(N__36103),
            .I(N__36047));
    InMux I__4918 (
            .O(N__36100),
            .I(N__36047));
    InMux I__4917 (
            .O(N__36099),
            .I(N__36047));
    InMux I__4916 (
            .O(N__36096),
            .I(N__36047));
    InMux I__4915 (
            .O(N__36095),
            .I(N__36047));
    InMux I__4914 (
            .O(N__36092),
            .I(N__36047));
    InMux I__4913 (
            .O(N__36091),
            .I(N__36047));
    LocalMux I__4912 (
            .O(N__36086),
            .I(N__36044));
    InMux I__4911 (
            .O(N__36085),
            .I(N__36041));
    CascadeMux I__4910 (
            .O(N__36084),
            .I(N__36038));
    CascadeMux I__4909 (
            .O(N__36083),
            .I(N__36034));
    CascadeMux I__4908 (
            .O(N__36082),
            .I(N__36030));
    CascadeMux I__4907 (
            .O(N__36081),
            .I(N__36026));
    CascadeMux I__4906 (
            .O(N__36080),
            .I(N__36023));
    CascadeMux I__4905 (
            .O(N__36079),
            .I(N__36019));
    CascadeMux I__4904 (
            .O(N__36078),
            .I(N__36015));
    LocalMux I__4903 (
            .O(N__36075),
            .I(N__36004));
    LocalMux I__4902 (
            .O(N__36064),
            .I(N__36004));
    LocalMux I__4901 (
            .O(N__36047),
            .I(N__36004));
    Span4Mux_v I__4900 (
            .O(N__36044),
            .I(N__36004));
    LocalMux I__4899 (
            .O(N__36041),
            .I(N__36004));
    InMux I__4898 (
            .O(N__36038),
            .I(N__35991));
    InMux I__4897 (
            .O(N__36037),
            .I(N__35991));
    InMux I__4896 (
            .O(N__36034),
            .I(N__35991));
    InMux I__4895 (
            .O(N__36033),
            .I(N__35991));
    InMux I__4894 (
            .O(N__36030),
            .I(N__35991));
    InMux I__4893 (
            .O(N__36029),
            .I(N__35991));
    InMux I__4892 (
            .O(N__36026),
            .I(N__35988));
    InMux I__4891 (
            .O(N__36023),
            .I(N__35977));
    InMux I__4890 (
            .O(N__36022),
            .I(N__35977));
    InMux I__4889 (
            .O(N__36019),
            .I(N__35977));
    InMux I__4888 (
            .O(N__36018),
            .I(N__35977));
    InMux I__4887 (
            .O(N__36015),
            .I(N__35977));
    Span4Mux_v I__4886 (
            .O(N__36004),
            .I(N__35973));
    LocalMux I__4885 (
            .O(N__35991),
            .I(N__35966));
    LocalMux I__4884 (
            .O(N__35988),
            .I(N__35966));
    LocalMux I__4883 (
            .O(N__35977),
            .I(N__35966));
    InMux I__4882 (
            .O(N__35976),
            .I(N__35963));
    Odrv4 I__4881 (
            .O(N__35973),
            .I(\foc.u_Park_Transform.n607 ));
    Odrv4 I__4880 (
            .O(N__35966),
            .I(\foc.u_Park_Transform.n607 ));
    LocalMux I__4879 (
            .O(N__35963),
            .I(\foc.u_Park_Transform.n607 ));
    CascadeMux I__4878 (
            .O(N__35956),
            .I(N__35953));
    InMux I__4877 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__4876 (
            .O(N__35950),
            .I(N__35947));
    Odrv4 I__4875 (
            .O(N__35947),
            .I(\foc.u_Park_Transform.n706_adj_2044 ));
    InMux I__4874 (
            .O(N__35944),
            .I(\foc.u_Park_Transform.n16990 ));
    InMux I__4873 (
            .O(N__35941),
            .I(N__35938));
    LocalMux I__4872 (
            .O(N__35938),
            .I(N__35935));
    Span4Mux_h I__4871 (
            .O(N__35935),
            .I(N__35931));
    InMux I__4870 (
            .O(N__35934),
            .I(N__35928));
    Span4Mux_v I__4869 (
            .O(N__35931),
            .I(N__35923));
    LocalMux I__4868 (
            .O(N__35928),
            .I(N__35923));
    Odrv4 I__4867 (
            .O(N__35923),
            .I(\foc.u_Park_Transform.n761 ));
    CascadeMux I__4866 (
            .O(N__35920),
            .I(N__35917));
    InMux I__4865 (
            .O(N__35917),
            .I(N__35914));
    LocalMux I__4864 (
            .O(N__35914),
            .I(N__35911));
    Odrv4 I__4863 (
            .O(N__35911),
            .I(\foc.u_Park_Transform.n709_adj_2066 ));
    CascadeMux I__4862 (
            .O(N__35908),
            .I(N__35905));
    InMux I__4861 (
            .O(N__35905),
            .I(N__35902));
    LocalMux I__4860 (
            .O(N__35902),
            .I(\foc.u_Park_Transform.n762_adj_2065 ));
    InMux I__4859 (
            .O(N__35899),
            .I(\foc.u_Park_Transform.n16991 ));
    CascadeMux I__4858 (
            .O(N__35896),
            .I(N__35880));
    CascadeMux I__4857 (
            .O(N__35895),
            .I(N__35876));
    CascadeMux I__4856 (
            .O(N__35894),
            .I(N__35872));
    CascadeMux I__4855 (
            .O(N__35893),
            .I(N__35867));
    CascadeMux I__4854 (
            .O(N__35892),
            .I(N__35864));
    CascadeMux I__4853 (
            .O(N__35891),
            .I(N__35861));
    CascadeMux I__4852 (
            .O(N__35890),
            .I(N__35858));
    CascadeMux I__4851 (
            .O(N__35889),
            .I(N__35855));
    CascadeMux I__4850 (
            .O(N__35888),
            .I(N__35851));
    CascadeMux I__4849 (
            .O(N__35887),
            .I(N__35847));
    CascadeMux I__4848 (
            .O(N__35886),
            .I(N__35843));
    CascadeMux I__4847 (
            .O(N__35885),
            .I(N__35839));
    CascadeMux I__4846 (
            .O(N__35884),
            .I(N__35835));
    CascadeMux I__4845 (
            .O(N__35883),
            .I(N__35832));
    InMux I__4844 (
            .O(N__35880),
            .I(N__35819));
    InMux I__4843 (
            .O(N__35879),
            .I(N__35819));
    InMux I__4842 (
            .O(N__35876),
            .I(N__35819));
    InMux I__4841 (
            .O(N__35875),
            .I(N__35819));
    InMux I__4840 (
            .O(N__35872),
            .I(N__35819));
    InMux I__4839 (
            .O(N__35871),
            .I(N__35819));
    InMux I__4838 (
            .O(N__35870),
            .I(N__35814));
    InMux I__4837 (
            .O(N__35867),
            .I(N__35814));
    InMux I__4836 (
            .O(N__35864),
            .I(N__35807));
    InMux I__4835 (
            .O(N__35861),
            .I(N__35804));
    InMux I__4834 (
            .O(N__35858),
            .I(N__35793));
    InMux I__4833 (
            .O(N__35855),
            .I(N__35793));
    InMux I__4832 (
            .O(N__35854),
            .I(N__35793));
    InMux I__4831 (
            .O(N__35851),
            .I(N__35793));
    InMux I__4830 (
            .O(N__35850),
            .I(N__35793));
    InMux I__4829 (
            .O(N__35847),
            .I(N__35778));
    InMux I__4828 (
            .O(N__35846),
            .I(N__35778));
    InMux I__4827 (
            .O(N__35843),
            .I(N__35778));
    InMux I__4826 (
            .O(N__35842),
            .I(N__35778));
    InMux I__4825 (
            .O(N__35839),
            .I(N__35778));
    InMux I__4824 (
            .O(N__35838),
            .I(N__35778));
    InMux I__4823 (
            .O(N__35835),
            .I(N__35778));
    InMux I__4822 (
            .O(N__35832),
            .I(N__35775));
    LocalMux I__4821 (
            .O(N__35819),
            .I(N__35770));
    LocalMux I__4820 (
            .O(N__35814),
            .I(N__35770));
    InMux I__4819 (
            .O(N__35813),
            .I(N__35767));
    CascadeMux I__4818 (
            .O(N__35812),
            .I(N__35763));
    CascadeMux I__4817 (
            .O(N__35811),
            .I(N__35759));
    CascadeMux I__4816 (
            .O(N__35810),
            .I(N__35755));
    LocalMux I__4815 (
            .O(N__35807),
            .I(N__35752));
    LocalMux I__4814 (
            .O(N__35804),
            .I(N__35743));
    LocalMux I__4813 (
            .O(N__35793),
            .I(N__35743));
    LocalMux I__4812 (
            .O(N__35778),
            .I(N__35743));
    LocalMux I__4811 (
            .O(N__35775),
            .I(N__35743));
    Span4Mux_h I__4810 (
            .O(N__35770),
            .I(N__35738));
    LocalMux I__4809 (
            .O(N__35767),
            .I(N__35738));
    InMux I__4808 (
            .O(N__35766),
            .I(N__35725));
    InMux I__4807 (
            .O(N__35763),
            .I(N__35725));
    InMux I__4806 (
            .O(N__35762),
            .I(N__35725));
    InMux I__4805 (
            .O(N__35759),
            .I(N__35725));
    InMux I__4804 (
            .O(N__35758),
            .I(N__35725));
    InMux I__4803 (
            .O(N__35755),
            .I(N__35725));
    Span4Mux_v I__4802 (
            .O(N__35752),
            .I(N__35722));
    Span12Mux_v I__4801 (
            .O(N__35743),
            .I(N__35719));
    Span4Mux_h I__4800 (
            .O(N__35738),
            .I(N__35714));
    LocalMux I__4799 (
            .O(N__35725),
            .I(N__35714));
    Odrv4 I__4798 (
            .O(N__35722),
            .I(\foc.u_Park_Transform.n610 ));
    Odrv12 I__4797 (
            .O(N__35719),
            .I(\foc.u_Park_Transform.n610 ));
    Odrv4 I__4796 (
            .O(N__35714),
            .I(\foc.u_Park_Transform.n610 ));
    CascadeMux I__4795 (
            .O(N__35707),
            .I(N__35704));
    InMux I__4794 (
            .O(N__35704),
            .I(N__35701));
    LocalMux I__4793 (
            .O(N__35701),
            .I(N__35698));
    Odrv12 I__4792 (
            .O(N__35698),
            .I(\foc.u_Park_Transform.n69_adj_2059 ));
    InMux I__4791 (
            .O(N__35695),
            .I(N__35692));
    LocalMux I__4790 (
            .O(N__35692),
            .I(\foc.u_Park_Transform.n72_adj_2062 ));
    CascadeMux I__4789 (
            .O(N__35689),
            .I(N__35686));
    InMux I__4788 (
            .O(N__35686),
            .I(N__35683));
    LocalMux I__4787 (
            .O(N__35683),
            .I(N__35680));
    Odrv4 I__4786 (
            .O(N__35680),
            .I(\foc.u_Park_Transform.n118_adj_2037 ));
    InMux I__4785 (
            .O(N__35677),
            .I(\foc.u_Park_Transform.n16978 ));
    CascadeMux I__4784 (
            .O(N__35674),
            .I(N__35671));
    InMux I__4783 (
            .O(N__35671),
            .I(N__35668));
    LocalMux I__4782 (
            .O(N__35668),
            .I(\foc.u_Park_Transform.n121_adj_2051 ));
    InMux I__4781 (
            .O(N__35665),
            .I(N__35662));
    LocalMux I__4780 (
            .O(N__35662),
            .I(N__35659));
    Odrv4 I__4779 (
            .O(N__35659),
            .I(\foc.u_Park_Transform.n167_adj_2029 ));
    InMux I__4778 (
            .O(N__35656),
            .I(\foc.u_Park_Transform.n16979 ));
    InMux I__4777 (
            .O(N__35653),
            .I(N__35650));
    LocalMux I__4776 (
            .O(N__35650),
            .I(\foc.u_Park_Transform.n170_adj_2048 ));
    CascadeMux I__4775 (
            .O(N__35647),
            .I(N__35644));
    InMux I__4774 (
            .O(N__35644),
            .I(N__35641));
    LocalMux I__4773 (
            .O(N__35641),
            .I(N__35638));
    Odrv12 I__4772 (
            .O(N__35638),
            .I(\foc.u_Park_Transform.n216_adj_2025 ));
    InMux I__4771 (
            .O(N__35635),
            .I(\foc.u_Park_Transform.n16980 ));
    CascadeMux I__4770 (
            .O(N__35632),
            .I(N__35629));
    InMux I__4769 (
            .O(N__35629),
            .I(N__35626));
    LocalMux I__4768 (
            .O(N__35626),
            .I(\foc.u_Park_Transform.n219_adj_2040 ));
    InMux I__4767 (
            .O(N__35623),
            .I(N__35620));
    LocalMux I__4766 (
            .O(N__35620),
            .I(N__35617));
    Odrv4 I__4765 (
            .O(N__35617),
            .I(\foc.u_Park_Transform.n265_adj_2023 ));
    InMux I__4764 (
            .O(N__35614),
            .I(\foc.u_Park_Transform.n16981 ));
    InMux I__4763 (
            .O(N__35611),
            .I(N__35608));
    LocalMux I__4762 (
            .O(N__35608),
            .I(\foc.u_Park_Transform.n268_adj_2027 ));
    CascadeMux I__4761 (
            .O(N__35605),
            .I(N__35602));
    InMux I__4760 (
            .O(N__35602),
            .I(N__35599));
    LocalMux I__4759 (
            .O(N__35599),
            .I(N__35596));
    Odrv4 I__4758 (
            .O(N__35596),
            .I(\foc.u_Park_Transform.n314_adj_2010 ));
    InMux I__4757 (
            .O(N__35593),
            .I(\foc.u_Park_Transform.n16982 ));
    CascadeMux I__4756 (
            .O(N__35590),
            .I(N__35587));
    InMux I__4755 (
            .O(N__35587),
            .I(N__35584));
    LocalMux I__4754 (
            .O(N__35584),
            .I(\foc.u_Park_Transform.n317_adj_2021 ));
    InMux I__4753 (
            .O(N__35581),
            .I(N__35578));
    LocalMux I__4752 (
            .O(N__35578),
            .I(N__35575));
    Odrv12 I__4751 (
            .O(N__35575),
            .I(\foc.u_Park_Transform.n363_adj_1998 ));
    InMux I__4750 (
            .O(N__35572),
            .I(\foc.u_Park_Transform.n16983 ));
    InMux I__4749 (
            .O(N__35569),
            .I(N__35566));
    LocalMux I__4748 (
            .O(N__35566),
            .I(\foc.u_Park_Transform.n366_adj_2013 ));
    InMux I__4747 (
            .O(N__35563),
            .I(\foc.u_Park_Transform.n16999 ));
    InMux I__4746 (
            .O(N__35560),
            .I(bfn_13_14_0_));
    InMux I__4745 (
            .O(N__35557),
            .I(\foc.u_Park_Transform.n17001 ));
    InMux I__4744 (
            .O(N__35554),
            .I(\foc.u_Park_Transform.n17002 ));
    InMux I__4743 (
            .O(N__35551),
            .I(\foc.u_Park_Transform.n17003 ));
    InMux I__4742 (
            .O(N__35548),
            .I(\foc.u_Park_Transform.n17004 ));
    InMux I__4741 (
            .O(N__35545),
            .I(\foc.u_Park_Transform.n17005 ));
    InMux I__4740 (
            .O(N__35542),
            .I(N__35538));
    InMux I__4739 (
            .O(N__35541),
            .I(N__35535));
    LocalMux I__4738 (
            .O(N__35538),
            .I(\foc.u_Park_Transform.n757 ));
    LocalMux I__4737 (
            .O(N__35535),
            .I(\foc.u_Park_Transform.n757 ));
    InMux I__4736 (
            .O(N__35530),
            .I(N__35527));
    LocalMux I__4735 (
            .O(N__35527),
            .I(N__35524));
    Odrv4 I__4734 (
            .O(N__35524),
            .I(\foc.u_Park_Transform.n758 ));
    InMux I__4733 (
            .O(N__35521),
            .I(\foc.u_Park_Transform.n17006 ));
    InMux I__4732 (
            .O(N__35518),
            .I(\foc.u_Park_Transform.n759 ));
    InMux I__4731 (
            .O(N__35515),
            .I(N__35512));
    LocalMux I__4730 (
            .O(N__35512),
            .I(N__35509));
    Span4Mux_v I__4729 (
            .O(N__35509),
            .I(N__35506));
    Odrv4 I__4728 (
            .O(N__35506),
            .I(\foc.u_Park_Transform.n759_THRU_CO ));
    CascadeMux I__4727 (
            .O(N__35503),
            .I(N__35500));
    InMux I__4726 (
            .O(N__35500),
            .I(N__35497));
    LocalMux I__4725 (
            .O(N__35497),
            .I(\foc.u_Park_Transform.n703_adj_2160 ));
    InMux I__4724 (
            .O(N__35494),
            .I(N__35491));
    LocalMux I__4723 (
            .O(N__35491),
            .I(N__35488));
    Odrv12 I__4722 (
            .O(N__35488),
            .I(\foc.u_Park_Transform.n754_adj_2159 ));
    InMux I__4721 (
            .O(N__35485),
            .I(\foc.u_Park_Transform.n17204 ));
    InMux I__4720 (
            .O(N__35482),
            .I(\foc.u_Park_Transform.n755_adj_2161 ));
    CascadeMux I__4719 (
            .O(N__35479),
            .I(N__35476));
    InMux I__4718 (
            .O(N__35476),
            .I(N__35473));
    LocalMux I__4717 (
            .O(N__35473),
            .I(N__35470));
    Odrv12 I__4716 (
            .O(N__35470),
            .I(\foc.u_Park_Transform.n755_adj_2161_THRU_CO ));
    InMux I__4715 (
            .O(N__35467),
            .I(\foc.u_Park_Transform.n16993 ));
    InMux I__4714 (
            .O(N__35464),
            .I(\foc.u_Park_Transform.n16994 ));
    InMux I__4713 (
            .O(N__35461),
            .I(\foc.u_Park_Transform.n16995 ));
    InMux I__4712 (
            .O(N__35458),
            .I(\foc.u_Park_Transform.n16996 ));
    InMux I__4711 (
            .O(N__35455),
            .I(\foc.u_Park_Transform.n16997 ));
    InMux I__4710 (
            .O(N__35452),
            .I(\foc.u_Park_Transform.n16998 ));
    CascadeMux I__4709 (
            .O(N__35449),
            .I(N__35446));
    InMux I__4708 (
            .O(N__35446),
            .I(N__35443));
    LocalMux I__4707 (
            .O(N__35443),
            .I(\foc.u_Park_Transform.n262_adj_1996 ));
    InMux I__4706 (
            .O(N__35440),
            .I(\foc.u_Park_Transform.n17195 ));
    CascadeMux I__4705 (
            .O(N__35437),
            .I(N__35434));
    InMux I__4704 (
            .O(N__35434),
            .I(N__35431));
    LocalMux I__4703 (
            .O(N__35431),
            .I(\foc.u_Park_Transform.n311 ));
    InMux I__4702 (
            .O(N__35428),
            .I(\foc.u_Park_Transform.n17196 ));
    CascadeMux I__4701 (
            .O(N__35425),
            .I(N__35422));
    InMux I__4700 (
            .O(N__35422),
            .I(N__35419));
    LocalMux I__4699 (
            .O(N__35419),
            .I(\foc.u_Park_Transform.n360 ));
    InMux I__4698 (
            .O(N__35416),
            .I(\foc.u_Park_Transform.n17197 ));
    InMux I__4697 (
            .O(N__35413),
            .I(N__35410));
    LocalMux I__4696 (
            .O(N__35410),
            .I(\foc.u_Park_Transform.n409 ));
    InMux I__4695 (
            .O(N__35407),
            .I(bfn_13_12_0_));
    CascadeMux I__4694 (
            .O(N__35404),
            .I(N__35401));
    InMux I__4693 (
            .O(N__35401),
            .I(N__35398));
    LocalMux I__4692 (
            .O(N__35398),
            .I(\foc.u_Park_Transform.n458 ));
    InMux I__4691 (
            .O(N__35395),
            .I(\foc.u_Park_Transform.n17199 ));
    InMux I__4690 (
            .O(N__35392),
            .I(N__35389));
    LocalMux I__4689 (
            .O(N__35389),
            .I(\foc.u_Park_Transform.n507_adj_2165 ));
    InMux I__4688 (
            .O(N__35386),
            .I(\foc.u_Park_Transform.n17200 ));
    CascadeMux I__4687 (
            .O(N__35383),
            .I(N__35380));
    InMux I__4686 (
            .O(N__35380),
            .I(N__35377));
    LocalMux I__4685 (
            .O(N__35377),
            .I(\foc.u_Park_Transform.n556_adj_2164 ));
    InMux I__4684 (
            .O(N__35374),
            .I(\foc.u_Park_Transform.n17201 ));
    InMux I__4683 (
            .O(N__35371),
            .I(N__35368));
    LocalMux I__4682 (
            .O(N__35368),
            .I(\foc.u_Park_Transform.n605_adj_2163 ));
    InMux I__4681 (
            .O(N__35365),
            .I(\foc.u_Park_Transform.n17202 ));
    CascadeMux I__4680 (
            .O(N__35362),
            .I(N__35359));
    InMux I__4679 (
            .O(N__35359),
            .I(N__35356));
    LocalMux I__4678 (
            .O(N__35356),
            .I(\foc.u_Park_Transform.n654_adj_2162 ));
    InMux I__4677 (
            .O(N__35353),
            .I(\foc.u_Park_Transform.n17203 ));
    InMux I__4676 (
            .O(N__35350),
            .I(N__35347));
    LocalMux I__4675 (
            .O(N__35347),
            .I(N__35344));
    Span4Mux_h I__4674 (
            .O(N__35344),
            .I(N__35341));
    Odrv4 I__4673 (
            .O(N__35341),
            .I(\foc.u_Park_Transform.n786_adj_2152 ));
    CascadeMux I__4672 (
            .O(N__35338),
            .I(N__35335));
    InMux I__4671 (
            .O(N__35335),
            .I(N__35332));
    LocalMux I__4670 (
            .O(N__35332),
            .I(N__35329));
    Odrv4 I__4669 (
            .O(N__35329),
            .I(\foc.u_Park_Transform.n783_THRU_CO ));
    InMux I__4668 (
            .O(N__35326),
            .I(\foc.u_Park_Transform.n17095 ));
    InMux I__4667 (
            .O(N__35323),
            .I(N__35320));
    LocalMux I__4666 (
            .O(N__35320),
            .I(N__35317));
    Span4Mux_h I__4665 (
            .O(N__35317),
            .I(N__35313));
    InMux I__4664 (
            .O(N__35316),
            .I(N__35310));
    Sp12to4 I__4663 (
            .O(N__35313),
            .I(N__35305));
    LocalMux I__4662 (
            .O(N__35310),
            .I(N__35305));
    Odrv12 I__4661 (
            .O(N__35305),
            .I(\foc.u_Park_Transform.n790 ));
    CascadeMux I__4660 (
            .O(N__35302),
            .I(N__35299));
    InMux I__4659 (
            .O(N__35299),
            .I(N__35296));
    LocalMux I__4658 (
            .O(N__35296),
            .I(N__35293));
    Span4Mux_v I__4657 (
            .O(N__35293),
            .I(N__35290));
    Odrv4 I__4656 (
            .O(N__35290),
            .I(\foc.u_Park_Transform.n787_adj_2149_THRU_CO ));
    InMux I__4655 (
            .O(N__35287),
            .I(\foc.u_Park_Transform.n17096 ));
    InMux I__4654 (
            .O(N__35284),
            .I(\foc.u_Park_Transform.n17097 ));
    InMux I__4653 (
            .O(N__35281),
            .I(N__35278));
    LocalMux I__4652 (
            .O(N__35278),
            .I(\foc.u_Park_Transform.n66 ));
    InMux I__4651 (
            .O(N__35275),
            .I(\foc.u_Park_Transform.n17191 ));
    CascadeMux I__4650 (
            .O(N__35272),
            .I(N__35269));
    InMux I__4649 (
            .O(N__35269),
            .I(N__35266));
    LocalMux I__4648 (
            .O(N__35266),
            .I(\foc.u_Park_Transform.n115 ));
    InMux I__4647 (
            .O(N__35263),
            .I(\foc.u_Park_Transform.n17192 ));
    CascadeMux I__4646 (
            .O(N__35260),
            .I(N__35257));
    InMux I__4645 (
            .O(N__35257),
            .I(N__35254));
    LocalMux I__4644 (
            .O(N__35254),
            .I(\foc.u_Park_Transform.n164 ));
    InMux I__4643 (
            .O(N__35251),
            .I(\foc.u_Park_Transform.n17193 ));
    CascadeMux I__4642 (
            .O(N__35248),
            .I(N__35245));
    InMux I__4641 (
            .O(N__35245),
            .I(N__35242));
    LocalMux I__4640 (
            .O(N__35242),
            .I(\foc.u_Park_Transform.n213 ));
    InMux I__4639 (
            .O(N__35239),
            .I(\foc.u_Park_Transform.n17194 ));
    InMux I__4638 (
            .O(N__35236),
            .I(\foc.u_Park_Transform.n17087 ));
    InMux I__4637 (
            .O(N__35233),
            .I(N__35230));
    LocalMux I__4636 (
            .O(N__35230),
            .I(N__35227));
    Span4Mux_v I__4635 (
            .O(N__35227),
            .I(N__35224));
    Odrv4 I__4634 (
            .O(N__35224),
            .I(\foc.u_Park_Transform.n758_adj_2168 ));
    InMux I__4633 (
            .O(N__35221),
            .I(\foc.u_Park_Transform.n17088 ));
    InMux I__4632 (
            .O(N__35218),
            .I(N__35215));
    LocalMux I__4631 (
            .O(N__35215),
            .I(N__35212));
    Span4Mux_v I__4630 (
            .O(N__35212),
            .I(N__35209));
    Odrv4 I__4629 (
            .O(N__35209),
            .I(\foc.u_Park_Transform.n759_adj_2166_THRU_CO ));
    CascadeMux I__4628 (
            .O(N__35206),
            .I(N__35203));
    InMux I__4627 (
            .O(N__35203),
            .I(N__35200));
    LocalMux I__4626 (
            .O(N__35200),
            .I(\foc.u_Park_Transform.n762 ));
    InMux I__4625 (
            .O(N__35197),
            .I(\foc.u_Park_Transform.n17089 ));
    InMux I__4624 (
            .O(N__35194),
            .I(N__35191));
    LocalMux I__4623 (
            .O(N__35191),
            .I(N__35188));
    Odrv12 I__4622 (
            .O(N__35188),
            .I(\foc.u_Park_Transform.n766 ));
    CascadeMux I__4621 (
            .O(N__35185),
            .I(N__35182));
    InMux I__4620 (
            .O(N__35182),
            .I(N__35179));
    LocalMux I__4619 (
            .O(N__35179),
            .I(\foc.u_Park_Transform.n763_THRU_CO ));
    InMux I__4618 (
            .O(N__35176),
            .I(bfn_13_10_0_));
    InMux I__4617 (
            .O(N__35173),
            .I(N__35170));
    LocalMux I__4616 (
            .O(N__35170),
            .I(N__35167));
    Span4Mux_h I__4615 (
            .O(N__35167),
            .I(N__35164));
    Odrv4 I__4614 (
            .O(N__35164),
            .I(\foc.u_Park_Transform.n770_adj_2030 ));
    CascadeMux I__4613 (
            .O(N__35161),
            .I(N__35158));
    InMux I__4612 (
            .O(N__35158),
            .I(N__35155));
    LocalMux I__4611 (
            .O(N__35155),
            .I(N__35152));
    Odrv12 I__4610 (
            .O(N__35152),
            .I(\foc.u_Park_Transform.n767_THRU_CO ));
    InMux I__4609 (
            .O(N__35149),
            .I(\foc.u_Park_Transform.n17091 ));
    InMux I__4608 (
            .O(N__35146),
            .I(N__35143));
    LocalMux I__4607 (
            .O(N__35143),
            .I(N__35140));
    Span4Mux_h I__4606 (
            .O(N__35140),
            .I(N__35137));
    Odrv4 I__4605 (
            .O(N__35137),
            .I(\foc.u_Park_Transform.n774_adj_2045 ));
    CascadeMux I__4604 (
            .O(N__35134),
            .I(N__35131));
    InMux I__4603 (
            .O(N__35131),
            .I(N__35128));
    LocalMux I__4602 (
            .O(N__35128),
            .I(N__35125));
    Span4Mux_h I__4601 (
            .O(N__35125),
            .I(N__35122));
    Odrv4 I__4600 (
            .O(N__35122),
            .I(\foc.u_Park_Transform.n771_adj_2032_THRU_CO ));
    InMux I__4599 (
            .O(N__35119),
            .I(\foc.u_Park_Transform.n17092 ));
    InMux I__4598 (
            .O(N__35116),
            .I(N__35113));
    LocalMux I__4597 (
            .O(N__35113),
            .I(N__35110));
    Odrv12 I__4596 (
            .O(N__35110),
            .I(\foc.u_Park_Transform.n778_adj_2068 ));
    CascadeMux I__4595 (
            .O(N__35107),
            .I(N__35104));
    InMux I__4594 (
            .O(N__35104),
            .I(N__35101));
    LocalMux I__4593 (
            .O(N__35101),
            .I(N__35098));
    Span4Mux_v I__4592 (
            .O(N__35098),
            .I(N__35095));
    Odrv4 I__4591 (
            .O(N__35095),
            .I(\foc.u_Park_Transform.n775_adj_2047_THRU_CO ));
    InMux I__4590 (
            .O(N__35092),
            .I(\foc.u_Park_Transform.n17093 ));
    InMux I__4589 (
            .O(N__35089),
            .I(N__35086));
    LocalMux I__4588 (
            .O(N__35086),
            .I(N__35083));
    Odrv4 I__4587 (
            .O(N__35083),
            .I(\foc.u_Park_Transform.n782_adj_2109 ));
    CascadeMux I__4586 (
            .O(N__35080),
            .I(N__35077));
    InMux I__4585 (
            .O(N__35077),
            .I(N__35074));
    LocalMux I__4584 (
            .O(N__35074),
            .I(N__35071));
    Odrv12 I__4583 (
            .O(N__35071),
            .I(\foc.u_Park_Transform.n779_adj_2070_THRU_CO ));
    InMux I__4582 (
            .O(N__35068),
            .I(\foc.u_Park_Transform.n17094 ));
    InMux I__4581 (
            .O(N__35065),
            .I(\foc.u_Park_Transform.n17083 ));
    InMux I__4580 (
            .O(N__35062),
            .I(\foc.u_Park_Transform.n17084 ));
    InMux I__4579 (
            .O(N__35059),
            .I(\foc.u_Park_Transform.n17085 ));
    InMux I__4578 (
            .O(N__35056),
            .I(\foc.u_Park_Transform.n17086 ));
    InMux I__4577 (
            .O(N__35053),
            .I(N__35050));
    LocalMux I__4576 (
            .O(N__35050),
            .I(N__35047));
    Odrv4 I__4575 (
            .O(N__35047),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n470 ));
    InMux I__4574 (
            .O(N__35044),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18115 ));
    InMux I__4573 (
            .O(N__35041),
            .I(N__35038));
    LocalMux I__4572 (
            .O(N__35038),
            .I(N__35035));
    Odrv4 I__4571 (
            .O(N__35035),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n519 ));
    InMux I__4570 (
            .O(N__35032),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18116 ));
    InMux I__4569 (
            .O(N__35029),
            .I(N__35026));
    LocalMux I__4568 (
            .O(N__35026),
            .I(N__35023));
    Odrv12 I__4567 (
            .O(N__35023),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n568 ));
    InMux I__4566 (
            .O(N__35020),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18117 ));
    InMux I__4565 (
            .O(N__35017),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18118 ));
    InMux I__4564 (
            .O(N__35014),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18119 ));
    CascadeMux I__4563 (
            .O(N__35011),
            .I(N__35007));
    CascadeMux I__4562 (
            .O(N__35010),
            .I(N__35004));
    InMux I__4561 (
            .O(N__35007),
            .I(N__35000));
    InMux I__4560 (
            .O(N__35004),
            .I(N__34995));
    InMux I__4559 (
            .O(N__35003),
            .I(N__34995));
    LocalMux I__4558 (
            .O(N__35000),
            .I(N__34990));
    LocalMux I__4557 (
            .O(N__34995),
            .I(N__34990));
    Odrv4 I__4556 (
            .O(N__34990),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n617 ));
    InMux I__4555 (
            .O(N__34987),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18120 ));
    InMux I__4554 (
            .O(N__34984),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598 ));
    InMux I__4553 (
            .O(N__34981),
            .I(N__34978));
    LocalMux I__4552 (
            .O(N__34978),
            .I(N__34975));
    Odrv12 I__4551 (
            .O(N__34975),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617 ));
    InMux I__4550 (
            .O(N__34972),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18107 ));
    InMux I__4549 (
            .O(N__34969),
            .I(N__34966));
    LocalMux I__4548 (
            .O(N__34966),
            .I(N__34963));
    Odrv4 I__4547 (
            .O(N__34963),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615 ));
    InMux I__4546 (
            .O(N__34960),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18108 ));
    InMux I__4545 (
            .O(N__34957),
            .I(N__34954));
    LocalMux I__4544 (
            .O(N__34954),
            .I(N__34951));
    Odrv12 I__4543 (
            .O(N__34951),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613 ));
    InMux I__4542 (
            .O(N__34948),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18109 ));
    InMux I__4541 (
            .O(N__34945),
            .I(N__34942));
    LocalMux I__4540 (
            .O(N__34942),
            .I(N__34939));
    Odrv12 I__4539 (
            .O(N__34939),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611 ));
    InMux I__4538 (
            .O(N__34936),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18110 ));
    InMux I__4537 (
            .O(N__34933),
            .I(N__34930));
    LocalMux I__4536 (
            .O(N__34930),
            .I(N__34927));
    Odrv4 I__4535 (
            .O(N__34927),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609 ));
    InMux I__4534 (
            .O(N__34924),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18111 ));
    InMux I__4533 (
            .O(N__34921),
            .I(N__34918));
    LocalMux I__4532 (
            .O(N__34918),
            .I(N__34915));
    Odrv4 I__4531 (
            .O(N__34915),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607 ));
    InMux I__4530 (
            .O(N__34912),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18112 ));
    InMux I__4529 (
            .O(N__34909),
            .I(N__34906));
    LocalMux I__4528 (
            .O(N__34906),
            .I(N__34903));
    Odrv4 I__4527 (
            .O(N__34903),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n372 ));
    InMux I__4526 (
            .O(N__34900),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18113 ));
    InMux I__4525 (
            .O(N__34897),
            .I(N__34894));
    LocalMux I__4524 (
            .O(N__34894),
            .I(N__34891));
    Odrv12 I__4523 (
            .O(N__34891),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n421 ));
    InMux I__4522 (
            .O(N__34888),
            .I(bfn_12_25_0_));
    InMux I__4521 (
            .O(N__34885),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17661 ));
    InMux I__4520 (
            .O(N__34882),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17662 ));
    InMux I__4519 (
            .O(N__34879),
            .I(bfn_12_23_0_));
    InMux I__4518 (
            .O(N__34876),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17664 ));
    InMux I__4517 (
            .O(N__34873),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17665 ));
    InMux I__4516 (
            .O(N__34870),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17666 ));
    InMux I__4515 (
            .O(N__34867),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17667 ));
    InMux I__4514 (
            .O(N__34864),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775 ));
    InMux I__4513 (
            .O(N__34861),
            .I(N__34858));
    LocalMux I__4512 (
            .O(N__34858),
            .I(N__34855));
    Odrv12 I__4511 (
            .O(N__34855),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017 ));
    InMux I__4510 (
            .O(N__34852),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382 ));
    InMux I__4509 (
            .O(N__34849),
            .I(N__34846));
    LocalMux I__4508 (
            .O(N__34846),
            .I(N__34843));
    Span4Mux_h I__4507 (
            .O(N__34843),
            .I(N__34840));
    Odrv4 I__4506 (
            .O(N__34840),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117 ));
    InMux I__4505 (
            .O(N__34837),
            .I(N__34834));
    LocalMux I__4504 (
            .O(N__34834),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219 ));
    InMux I__4503 (
            .O(N__34831),
            .I(bfn_12_20_0_));
    InMux I__4502 (
            .O(N__34828),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220 ));
    CascadeMux I__4501 (
            .O(N__34825),
            .I(N__34822));
    InMux I__4500 (
            .O(N__34822),
            .I(N__34819));
    LocalMux I__4499 (
            .O(N__34819),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO ));
    InMux I__4498 (
            .O(N__34816),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17656 ));
    InMux I__4497 (
            .O(N__34813),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17657 ));
    InMux I__4496 (
            .O(N__34810),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17658 ));
    InMux I__4495 (
            .O(N__34807),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17659 ));
    InMux I__4494 (
            .O(N__34804),
            .I(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17660 ));
    InMux I__4493 (
            .O(N__34801),
            .I(\foc.u_Park_Transform.n16914 ));
    InMux I__4492 (
            .O(N__34798),
            .I(N__34792));
    CascadeMux I__4491 (
            .O(N__34797),
            .I(N__34788));
    CascadeMux I__4490 (
            .O(N__34796),
            .I(N__34784));
    CascadeMux I__4489 (
            .O(N__34795),
            .I(N__34780));
    LocalMux I__4488 (
            .O(N__34792),
            .I(N__34776));
    InMux I__4487 (
            .O(N__34791),
            .I(N__34761));
    InMux I__4486 (
            .O(N__34788),
            .I(N__34761));
    InMux I__4485 (
            .O(N__34787),
            .I(N__34761));
    InMux I__4484 (
            .O(N__34784),
            .I(N__34761));
    InMux I__4483 (
            .O(N__34783),
            .I(N__34761));
    InMux I__4482 (
            .O(N__34780),
            .I(N__34761));
    InMux I__4481 (
            .O(N__34779),
            .I(N__34761));
    Odrv4 I__4480 (
            .O(N__34776),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816 ));
    LocalMux I__4479 (
            .O(N__34761),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816 ));
    CascadeMux I__4478 (
            .O(N__34756),
            .I(N__34753));
    InMux I__4477 (
            .O(N__34753),
            .I(N__34750));
    LocalMux I__4476 (
            .O(N__34750),
            .I(N__34747));
    Odrv4 I__4475 (
            .O(N__34747),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417 ));
    InMux I__4474 (
            .O(N__34744),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376 ));
    InMux I__4473 (
            .O(N__34741),
            .I(N__34738));
    LocalMux I__4472 (
            .O(N__34738),
            .I(N__34735));
    Odrv4 I__4471 (
            .O(N__34735),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517 ));
    InMux I__4470 (
            .O(N__34732),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377 ));
    CascadeMux I__4469 (
            .O(N__34729),
            .I(N__34726));
    InMux I__4468 (
            .O(N__34726),
            .I(N__34723));
    LocalMux I__4467 (
            .O(N__34723),
            .I(N__34720));
    Odrv12 I__4466 (
            .O(N__34720),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617 ));
    InMux I__4465 (
            .O(N__34717),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378 ));
    InMux I__4464 (
            .O(N__34714),
            .I(N__34711));
    LocalMux I__4463 (
            .O(N__34711),
            .I(N__34708));
    Odrv12 I__4462 (
            .O(N__34708),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717 ));
    InMux I__4461 (
            .O(N__34705),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379 ));
    InMux I__4460 (
            .O(N__34702),
            .I(N__34699));
    LocalMux I__4459 (
            .O(N__34699),
            .I(N__34696));
    Odrv4 I__4458 (
            .O(N__34696),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817 ));
    InMux I__4457 (
            .O(N__34693),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380 ));
    InMux I__4456 (
            .O(N__34690),
            .I(N__34687));
    LocalMux I__4455 (
            .O(N__34687),
            .I(N__34684));
    Odrv12 I__4454 (
            .O(N__34684),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917 ));
    InMux I__4453 (
            .O(N__34681),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381 ));
    InMux I__4452 (
            .O(N__34678),
            .I(\foc.u_Park_Transform.n16905 ));
    InMux I__4451 (
            .O(N__34675),
            .I(\foc.u_Park_Transform.n16906 ));
    InMux I__4450 (
            .O(N__34672),
            .I(N__34669));
    LocalMux I__4449 (
            .O(N__34669),
            .I(N__34666));
    Odrv12 I__4448 (
            .O(N__34666),
            .I(\foc.u_Park_Transform.n766_adj_2053 ));
    InMux I__4447 (
            .O(N__34663),
            .I(bfn_12_18_0_));
    InMux I__4446 (
            .O(N__34660),
            .I(N__34657));
    LocalMux I__4445 (
            .O(N__34657),
            .I(N__34654));
    Odrv4 I__4444 (
            .O(N__34654),
            .I(\foc.u_Park_Transform.n770 ));
    CascadeMux I__4443 (
            .O(N__34651),
            .I(N__34648));
    InMux I__4442 (
            .O(N__34648),
            .I(N__34645));
    LocalMux I__4441 (
            .O(N__34645),
            .I(N__34642));
    Odrv4 I__4440 (
            .O(N__34642),
            .I(\foc.u_Park_Transform.n767_adj_2041_THRU_CO ));
    InMux I__4439 (
            .O(N__34639),
            .I(\foc.u_Park_Transform.n16908 ));
    InMux I__4438 (
            .O(N__34636),
            .I(N__34633));
    LocalMux I__4437 (
            .O(N__34633),
            .I(N__34630));
    Span4Mux_h I__4436 (
            .O(N__34630),
            .I(N__34627));
    Odrv4 I__4435 (
            .O(N__34627),
            .I(\foc.u_Park_Transform.n774 ));
    CascadeMux I__4434 (
            .O(N__34624),
            .I(N__34621));
    InMux I__4433 (
            .O(N__34621),
            .I(N__34618));
    LocalMux I__4432 (
            .O(N__34618),
            .I(N__34615));
    Odrv4 I__4431 (
            .O(N__34615),
            .I(\foc.u_Park_Transform.n771_THRU_CO ));
    InMux I__4430 (
            .O(N__34612),
            .I(\foc.u_Park_Transform.n16909 ));
    InMux I__4429 (
            .O(N__34609),
            .I(N__34606));
    LocalMux I__4428 (
            .O(N__34606),
            .I(N__34603));
    Odrv12 I__4427 (
            .O(N__34603),
            .I(\foc.u_Park_Transform.n778 ));
    CascadeMux I__4426 (
            .O(N__34600),
            .I(N__34597));
    InMux I__4425 (
            .O(N__34597),
            .I(N__34594));
    LocalMux I__4424 (
            .O(N__34594),
            .I(N__34591));
    Span12Mux_v I__4423 (
            .O(N__34591),
            .I(N__34588));
    Odrv12 I__4422 (
            .O(N__34588),
            .I(\foc.u_Park_Transform.n775_THRU_CO ));
    InMux I__4421 (
            .O(N__34585),
            .I(\foc.u_Park_Transform.n16910 ));
    InMux I__4420 (
            .O(N__34582),
            .I(N__34579));
    LocalMux I__4419 (
            .O(N__34579),
            .I(N__34576));
    Span4Mux_h I__4418 (
            .O(N__34576),
            .I(N__34573));
    Odrv4 I__4417 (
            .O(N__34573),
            .I(\foc.u_Park_Transform.n782 ));
    CascadeMux I__4416 (
            .O(N__34570),
            .I(N__34567));
    InMux I__4415 (
            .O(N__34567),
            .I(N__34564));
    LocalMux I__4414 (
            .O(N__34564),
            .I(N__34561));
    Odrv12 I__4413 (
            .O(N__34561),
            .I(\foc.u_Park_Transform.n779_THRU_CO ));
    InMux I__4412 (
            .O(N__34558),
            .I(\foc.u_Park_Transform.n16911 ));
    InMux I__4411 (
            .O(N__34555),
            .I(N__34552));
    LocalMux I__4410 (
            .O(N__34552),
            .I(N__34549));
    Span12Mux_v I__4409 (
            .O(N__34549),
            .I(N__34546));
    Odrv12 I__4408 (
            .O(N__34546),
            .I(\foc.u_Park_Transform.n786 ));
    CascadeMux I__4407 (
            .O(N__34543),
            .I(N__34540));
    InMux I__4406 (
            .O(N__34540),
            .I(N__34537));
    LocalMux I__4405 (
            .O(N__34537),
            .I(N__34534));
    Span4Mux_v I__4404 (
            .O(N__34534),
            .I(N__34531));
    Odrv4 I__4403 (
            .O(N__34531),
            .I(\foc.u_Park_Transform.n783_adj_2167_THRU_CO ));
    InMux I__4402 (
            .O(N__34528),
            .I(\foc.u_Park_Transform.n16912 ));
    CascadeMux I__4401 (
            .O(N__34525),
            .I(N__34522));
    InMux I__4400 (
            .O(N__34522),
            .I(N__34519));
    LocalMux I__4399 (
            .O(N__34519),
            .I(N__34516));
    Span4Mux_v I__4398 (
            .O(N__34516),
            .I(N__34513));
    Odrv4 I__4397 (
            .O(N__34513),
            .I(\foc.u_Park_Transform.n787_THRU_CO ));
    InMux I__4396 (
            .O(N__34510),
            .I(\foc.u_Park_Transform.n16913 ));
    InMux I__4395 (
            .O(N__34507),
            .I(\foc.u_Park_Transform.n16975 ));
    InMux I__4394 (
            .O(N__34504),
            .I(N__34501));
    LocalMux I__4393 (
            .O(N__34501),
            .I(N__34497));
    InMux I__4392 (
            .O(N__34500),
            .I(N__34494));
    Span4Mux_v I__4391 (
            .O(N__34497),
            .I(N__34491));
    LocalMux I__4390 (
            .O(N__34494),
            .I(N__34488));
    Odrv4 I__4389 (
            .O(N__34491),
            .I(\foc.u_Park_Transform.n765 ));
    Odrv4 I__4388 (
            .O(N__34488),
            .I(\foc.u_Park_Transform.n765 ));
    CascadeMux I__4387 (
            .O(N__34483),
            .I(N__34480));
    InMux I__4386 (
            .O(N__34480),
            .I(N__34477));
    LocalMux I__4385 (
            .O(N__34477),
            .I(\foc.u_Park_Transform.n712 ));
    InMux I__4384 (
            .O(N__34474),
            .I(\foc.u_Park_Transform.n16976 ));
    InMux I__4383 (
            .O(N__34471),
            .I(\foc.u_Park_Transform.n767_adj_2041 ));
    InMux I__4382 (
            .O(N__34468),
            .I(\foc.u_Park_Transform.n16900 ));
    InMux I__4381 (
            .O(N__34465),
            .I(\foc.u_Park_Transform.n16901 ));
    InMux I__4380 (
            .O(N__34462),
            .I(\foc.u_Park_Transform.n16902 ));
    InMux I__4379 (
            .O(N__34459),
            .I(\foc.u_Park_Transform.n16903 ));
    InMux I__4378 (
            .O(N__34456),
            .I(\foc.u_Park_Transform.n16904 ));
    InMux I__4377 (
            .O(N__34453),
            .I(N__34450));
    LocalMux I__4376 (
            .O(N__34450),
            .I(\foc.u_Park_Transform.n271_adj_2043 ));
    InMux I__4375 (
            .O(N__34447),
            .I(\foc.u_Park_Transform.n16967 ));
    CascadeMux I__4374 (
            .O(N__34444),
            .I(N__34441));
    InMux I__4373 (
            .O(N__34441),
            .I(N__34438));
    LocalMux I__4372 (
            .O(N__34438),
            .I(\foc.u_Park_Transform.n320_adj_2036 ));
    InMux I__4371 (
            .O(N__34435),
            .I(\foc.u_Park_Transform.n16968 ));
    InMux I__4370 (
            .O(N__34432),
            .I(N__34429));
    LocalMux I__4369 (
            .O(N__34429),
            .I(\foc.u_Park_Transform.n369_adj_2026 ));
    InMux I__4368 (
            .O(N__34426),
            .I(\foc.u_Park_Transform.n16969 ));
    CascadeMux I__4367 (
            .O(N__34423),
            .I(N__34420));
    InMux I__4366 (
            .O(N__34420),
            .I(N__34417));
    LocalMux I__4365 (
            .O(N__34417),
            .I(\foc.u_Park_Transform.n418 ));
    InMux I__4364 (
            .O(N__34414),
            .I(bfn_12_16_0_));
    InMux I__4363 (
            .O(N__34411),
            .I(N__34408));
    LocalMux I__4362 (
            .O(N__34408),
            .I(\foc.u_Park_Transform.n467 ));
    InMux I__4361 (
            .O(N__34405),
            .I(\foc.u_Park_Transform.n16971 ));
    CascadeMux I__4360 (
            .O(N__34402),
            .I(N__34399));
    InMux I__4359 (
            .O(N__34399),
            .I(N__34396));
    LocalMux I__4358 (
            .O(N__34396),
            .I(\foc.u_Park_Transform.n516 ));
    InMux I__4357 (
            .O(N__34393),
            .I(\foc.u_Park_Transform.n16972 ));
    InMux I__4356 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__4355 (
            .O(N__34387),
            .I(\foc.u_Park_Transform.n565_adj_2020 ));
    InMux I__4354 (
            .O(N__34384),
            .I(\foc.u_Park_Transform.n16973 ));
    InMux I__4353 (
            .O(N__34381),
            .I(N__34378));
    LocalMux I__4352 (
            .O(N__34378),
            .I(\foc.u_Park_Transform.n614 ));
    InMux I__4351 (
            .O(N__34375),
            .I(\foc.u_Park_Transform.n16974 ));
    InMux I__4350 (
            .O(N__34372),
            .I(N__34369));
    LocalMux I__4349 (
            .O(N__34369),
            .I(\foc.u_Park_Transform.n663 ));
    CascadeMux I__4348 (
            .O(N__34366),
            .I(n4_cascade_));
    CascadeMux I__4347 (
            .O(N__34363),
            .I(N__34357));
    CascadeMux I__4346 (
            .O(N__34362),
            .I(N__34353));
    CascadeMux I__4345 (
            .O(N__34361),
            .I(N__34350));
    CascadeMux I__4344 (
            .O(N__34360),
            .I(N__34346));
    InMux I__4343 (
            .O(N__34357),
            .I(N__34339));
    InMux I__4342 (
            .O(N__34356),
            .I(N__34339));
    InMux I__4341 (
            .O(N__34353),
            .I(N__34339));
    InMux I__4340 (
            .O(N__34350),
            .I(N__34332));
    InMux I__4339 (
            .O(N__34349),
            .I(N__34332));
    InMux I__4338 (
            .O(N__34346),
            .I(N__34332));
    LocalMux I__4337 (
            .O(N__34339),
            .I(N__34329));
    LocalMux I__4336 (
            .O(N__34332),
            .I(N__34326));
    Odrv4 I__4335 (
            .O(N__34329),
            .I(\foc.u_Park_Transform.n237 ));
    Odrv12 I__4334 (
            .O(N__34326),
            .I(\foc.u_Park_Transform.n237 ));
    CascadeMux I__4333 (
            .O(N__34321),
            .I(N__34318));
    InMux I__4332 (
            .O(N__34318),
            .I(N__34314));
    CascadeMux I__4331 (
            .O(N__34317),
            .I(N__34311));
    LocalMux I__4330 (
            .O(N__34314),
            .I(N__34308));
    InMux I__4329 (
            .O(N__34311),
            .I(N__34305));
    Span4Mux_h I__4328 (
            .O(N__34308),
            .I(N__34302));
    LocalMux I__4327 (
            .O(N__34305),
            .I(N__34299));
    Odrv4 I__4326 (
            .O(N__34302),
            .I(\foc.u_Park_Transform.n188 ));
    Odrv12 I__4325 (
            .O(N__34299),
            .I(\foc.u_Park_Transform.n188 ));
    CascadeMux I__4324 (
            .O(N__34294),
            .I(N__34288));
    CascadeMux I__4323 (
            .O(N__34293),
            .I(N__34285));
    CascadeMux I__4322 (
            .O(N__34292),
            .I(N__34281));
    InMux I__4321 (
            .O(N__34291),
            .I(N__34267));
    InMux I__4320 (
            .O(N__34288),
            .I(N__34267));
    InMux I__4319 (
            .O(N__34285),
            .I(N__34258));
    InMux I__4318 (
            .O(N__34284),
            .I(N__34258));
    InMux I__4317 (
            .O(N__34281),
            .I(N__34258));
    InMux I__4316 (
            .O(N__34280),
            .I(N__34258));
    InMux I__4315 (
            .O(N__34279),
            .I(N__34255));
    InMux I__4314 (
            .O(N__34278),
            .I(N__34252));
    CascadeMux I__4313 (
            .O(N__34277),
            .I(N__34246));
    CascadeMux I__4312 (
            .O(N__34276),
            .I(N__34240));
    CascadeMux I__4311 (
            .O(N__34275),
            .I(N__34237));
    CascadeMux I__4310 (
            .O(N__34274),
            .I(N__34233));
    CascadeMux I__4309 (
            .O(N__34273),
            .I(N__34229));
    CascadeMux I__4308 (
            .O(N__34272),
            .I(N__34224));
    LocalMux I__4307 (
            .O(N__34267),
            .I(N__34216));
    LocalMux I__4306 (
            .O(N__34258),
            .I(N__34216));
    LocalMux I__4305 (
            .O(N__34255),
            .I(N__34213));
    LocalMux I__4304 (
            .O(N__34252),
            .I(N__34210));
    InMux I__4303 (
            .O(N__34251),
            .I(N__34201));
    InMux I__4302 (
            .O(N__34250),
            .I(N__34201));
    InMux I__4301 (
            .O(N__34249),
            .I(N__34201));
    InMux I__4300 (
            .O(N__34246),
            .I(N__34201));
    InMux I__4299 (
            .O(N__34245),
            .I(N__34192));
    InMux I__4298 (
            .O(N__34244),
            .I(N__34192));
    InMux I__4297 (
            .O(N__34243),
            .I(N__34192));
    InMux I__4296 (
            .O(N__34240),
            .I(N__34192));
    InMux I__4295 (
            .O(N__34237),
            .I(N__34179));
    InMux I__4294 (
            .O(N__34236),
            .I(N__34179));
    InMux I__4293 (
            .O(N__34233),
            .I(N__34179));
    InMux I__4292 (
            .O(N__34232),
            .I(N__34179));
    InMux I__4291 (
            .O(N__34229),
            .I(N__34179));
    InMux I__4290 (
            .O(N__34228),
            .I(N__34179));
    InMux I__4289 (
            .O(N__34227),
            .I(N__34174));
    InMux I__4288 (
            .O(N__34224),
            .I(N__34174));
    CascadeMux I__4287 (
            .O(N__34223),
            .I(N__34170));
    CascadeMux I__4286 (
            .O(N__34222),
            .I(N__34166));
    CascadeMux I__4285 (
            .O(N__34221),
            .I(N__34162));
    Span4Mux_v I__4284 (
            .O(N__34216),
            .I(N__34151));
    Span4Mux_h I__4283 (
            .O(N__34213),
            .I(N__34151));
    Span4Mux_v I__4282 (
            .O(N__34210),
            .I(N__34151));
    LocalMux I__4281 (
            .O(N__34201),
            .I(N__34151));
    LocalMux I__4280 (
            .O(N__34192),
            .I(N__34151));
    LocalMux I__4279 (
            .O(N__34179),
            .I(N__34146));
    LocalMux I__4278 (
            .O(N__34174),
            .I(N__34146));
    InMux I__4277 (
            .O(N__34173),
            .I(N__34133));
    InMux I__4276 (
            .O(N__34170),
            .I(N__34133));
    InMux I__4275 (
            .O(N__34169),
            .I(N__34133));
    InMux I__4274 (
            .O(N__34166),
            .I(N__34133));
    InMux I__4273 (
            .O(N__34165),
            .I(N__34133));
    InMux I__4272 (
            .O(N__34162),
            .I(N__34133));
    Odrv4 I__4271 (
            .O(N__34151),
            .I(\foc.u_Park_Transform.n613 ));
    Odrv4 I__4270 (
            .O(N__34146),
            .I(\foc.u_Park_Transform.n613 ));
    LocalMux I__4269 (
            .O(N__34133),
            .I(\foc.u_Park_Transform.n613 ));
    InMux I__4268 (
            .O(N__34126),
            .I(N__34123));
    LocalMux I__4267 (
            .O(N__34123),
            .I(\foc.u_Park_Transform.n75_adj_2123 ));
    InMux I__4266 (
            .O(N__34120),
            .I(\foc.u_Park_Transform.n16963 ));
    CascadeMux I__4265 (
            .O(N__34117),
            .I(N__34114));
    InMux I__4264 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__4263 (
            .O(N__34111),
            .I(\foc.u_Park_Transform.n124_adj_2090 ));
    InMux I__4262 (
            .O(N__34108),
            .I(\foc.u_Park_Transform.n16964 ));
    InMux I__4261 (
            .O(N__34105),
            .I(N__34102));
    LocalMux I__4260 (
            .O(N__34102),
            .I(\foc.u_Park_Transform.n173_adj_2061 ));
    InMux I__4259 (
            .O(N__34099),
            .I(\foc.u_Park_Transform.n16965 ));
    CascadeMux I__4258 (
            .O(N__34096),
            .I(N__34093));
    InMux I__4257 (
            .O(N__34093),
            .I(N__34090));
    LocalMux I__4256 (
            .O(N__34090),
            .I(\foc.u_Park_Transform.n222_adj_2049 ));
    InMux I__4255 (
            .O(N__34087),
            .I(\foc.u_Park_Transform.n16966 ));
    InMux I__4254 (
            .O(N__34084),
            .I(N__34078));
    InMux I__4253 (
            .O(N__34083),
            .I(N__34078));
    LocalMux I__4252 (
            .O(N__34078),
            .I(\foc.Look_Up_Table_out1_1_3 ));
    InMux I__4251 (
            .O(N__34075),
            .I(N__34069));
    InMux I__4250 (
            .O(N__34074),
            .I(N__34069));
    LocalMux I__4249 (
            .O(N__34069),
            .I(\foc.Look_Up_Table_out1_1_5 ));
    InMux I__4248 (
            .O(N__34066),
            .I(N__34060));
    InMux I__4247 (
            .O(N__34065),
            .I(N__34060));
    LocalMux I__4246 (
            .O(N__34060),
            .I(\foc.Look_Up_Table_out1_1_4 ));
    CascadeMux I__4245 (
            .O(N__34057),
            .I(N__34054));
    InMux I__4244 (
            .O(N__34054),
            .I(N__34051));
    LocalMux I__4243 (
            .O(N__34051),
            .I(N__34048));
    Odrv4 I__4242 (
            .O(N__34048),
            .I(\foc.u_Park_Transform.n412 ));
    InMux I__4241 (
            .O(N__34045),
            .I(bfn_12_12_0_));
    InMux I__4240 (
            .O(N__34042),
            .I(N__34039));
    LocalMux I__4239 (
            .O(N__34039),
            .I(N__34036));
    Odrv4 I__4238 (
            .O(N__34036),
            .I(\foc.u_Park_Transform.n461 ));
    InMux I__4237 (
            .O(N__34033),
            .I(\foc.u_Park_Transform.n17184 ));
    CascadeMux I__4236 (
            .O(N__34030),
            .I(N__34027));
    InMux I__4235 (
            .O(N__34027),
            .I(N__34024));
    LocalMux I__4234 (
            .O(N__34024),
            .I(N__34021));
    Odrv12 I__4233 (
            .O(N__34021),
            .I(\foc.u_Park_Transform.n510_adj_2004 ));
    InMux I__4232 (
            .O(N__34018),
            .I(\foc.u_Park_Transform.n17185 ));
    InMux I__4231 (
            .O(N__34015),
            .I(N__34012));
    LocalMux I__4230 (
            .O(N__34012),
            .I(N__34009));
    Odrv12 I__4229 (
            .O(N__34009),
            .I(\foc.u_Park_Transform.n559_adj_2001 ));
    InMux I__4228 (
            .O(N__34006),
            .I(\foc.u_Park_Transform.n17186 ));
    InMux I__4227 (
            .O(N__34003),
            .I(N__34000));
    LocalMux I__4226 (
            .O(N__34000),
            .I(N__33997));
    Odrv4 I__4225 (
            .O(N__33997),
            .I(\foc.u_Park_Transform.n608 ));
    InMux I__4224 (
            .O(N__33994),
            .I(\foc.u_Park_Transform.n17187 ));
    InMux I__4223 (
            .O(N__33991),
            .I(N__33988));
    LocalMux I__4222 (
            .O(N__33988),
            .I(N__33985));
    Odrv4 I__4221 (
            .O(N__33985),
            .I(\foc.u_Park_Transform.n657 ));
    InMux I__4220 (
            .O(N__33982),
            .I(\foc.u_Park_Transform.n17188 ));
    CascadeMux I__4219 (
            .O(N__33979),
            .I(N__33976));
    InMux I__4218 (
            .O(N__33976),
            .I(N__33973));
    LocalMux I__4217 (
            .O(N__33973),
            .I(N__33970));
    Odrv4 I__4216 (
            .O(N__33970),
            .I(\foc.u_Park_Transform.n706 ));
    InMux I__4215 (
            .O(N__33967),
            .I(\foc.u_Park_Transform.n17189 ));
    InMux I__4214 (
            .O(N__33964),
            .I(\foc.u_Park_Transform.n759_adj_2166 ));
    InMux I__4213 (
            .O(N__33961),
            .I(\foc.u_Park_Transform.n763 ));
    CascadeMux I__4212 (
            .O(N__33958),
            .I(N__33955));
    InMux I__4211 (
            .O(N__33955),
            .I(N__33952));
    LocalMux I__4210 (
            .O(N__33952),
            .I(N__33949));
    Odrv4 I__4209 (
            .O(N__33949),
            .I(\foc.u_Park_Transform.n69 ));
    InMux I__4208 (
            .O(N__33946),
            .I(\foc.u_Park_Transform.n17176 ));
    CascadeMux I__4207 (
            .O(N__33943),
            .I(N__33940));
    InMux I__4206 (
            .O(N__33940),
            .I(N__33937));
    LocalMux I__4205 (
            .O(N__33937),
            .I(N__33934));
    Odrv4 I__4204 (
            .O(N__33934),
            .I(\foc.u_Park_Transform.n118 ));
    InMux I__4203 (
            .O(N__33931),
            .I(\foc.u_Park_Transform.n17177 ));
    InMux I__4202 (
            .O(N__33928),
            .I(N__33925));
    LocalMux I__4201 (
            .O(N__33925),
            .I(N__33922));
    Odrv12 I__4200 (
            .O(N__33922),
            .I(\foc.u_Park_Transform.n167 ));
    InMux I__4199 (
            .O(N__33919),
            .I(\foc.u_Park_Transform.n17178 ));
    CascadeMux I__4198 (
            .O(N__33916),
            .I(N__33913));
    InMux I__4197 (
            .O(N__33913),
            .I(N__33910));
    LocalMux I__4196 (
            .O(N__33910),
            .I(N__33907));
    Odrv12 I__4195 (
            .O(N__33907),
            .I(\foc.u_Park_Transform.n216 ));
    InMux I__4194 (
            .O(N__33904),
            .I(\foc.u_Park_Transform.n17179 ));
    InMux I__4193 (
            .O(N__33901),
            .I(N__33898));
    LocalMux I__4192 (
            .O(N__33898),
            .I(N__33895));
    Odrv4 I__4191 (
            .O(N__33895),
            .I(\foc.u_Park_Transform.n265 ));
    InMux I__4190 (
            .O(N__33892),
            .I(\foc.u_Park_Transform.n17180 ));
    CascadeMux I__4189 (
            .O(N__33889),
            .I(N__33886));
    InMux I__4188 (
            .O(N__33886),
            .I(N__33883));
    LocalMux I__4187 (
            .O(N__33883),
            .I(N__33880));
    Odrv4 I__4186 (
            .O(N__33880),
            .I(\foc.u_Park_Transform.n314 ));
    InMux I__4185 (
            .O(N__33877),
            .I(\foc.u_Park_Transform.n17181 ));
    InMux I__4184 (
            .O(N__33874),
            .I(N__33871));
    LocalMux I__4183 (
            .O(N__33871),
            .I(N__33868));
    Odrv4 I__4182 (
            .O(N__33868),
            .I(\foc.u_Park_Transform.n363 ));
    InMux I__4181 (
            .O(N__33865),
            .I(\foc.u_Park_Transform.n17182 ));
    InMux I__4180 (
            .O(N__33862),
            .I(N__33859));
    LocalMux I__4179 (
            .O(N__33859),
            .I(N__33856));
    Odrv4 I__4178 (
            .O(N__33856),
            .I(\foc.u_Park_Transform.n366 ));
    InMux I__4177 (
            .O(N__33853),
            .I(\foc.u_Park_Transform.n17167 ));
    InMux I__4176 (
            .O(N__33850),
            .I(N__33847));
    LocalMux I__4175 (
            .O(N__33847),
            .I(N__33844));
    Span4Mux_v I__4174 (
            .O(N__33844),
            .I(N__33841));
    Odrv4 I__4173 (
            .O(N__33841),
            .I(\foc.u_Park_Transform.n415_adj_2008 ));
    InMux I__4172 (
            .O(N__33838),
            .I(bfn_12_10_0_));
    CascadeMux I__4171 (
            .O(N__33835),
            .I(N__33832));
    InMux I__4170 (
            .O(N__33832),
            .I(N__33829));
    LocalMux I__4169 (
            .O(N__33829),
            .I(N__33826));
    Odrv4 I__4168 (
            .O(N__33826),
            .I(\foc.u_Park_Transform.n464_adj_2005 ));
    InMux I__4167 (
            .O(N__33823),
            .I(\foc.u_Park_Transform.n17169 ));
    InMux I__4166 (
            .O(N__33820),
            .I(N__33817));
    LocalMux I__4165 (
            .O(N__33817),
            .I(N__33814));
    Odrv4 I__4164 (
            .O(N__33814),
            .I(\foc.u_Park_Transform.n513_adj_2002 ));
    InMux I__4163 (
            .O(N__33811),
            .I(\foc.u_Park_Transform.n17170 ));
    CascadeMux I__4162 (
            .O(N__33808),
            .I(N__33805));
    InMux I__4161 (
            .O(N__33805),
            .I(N__33802));
    LocalMux I__4160 (
            .O(N__33802),
            .I(N__33799));
    Odrv12 I__4159 (
            .O(N__33799),
            .I(\foc.u_Park_Transform.n562_adj_2000 ));
    InMux I__4158 (
            .O(N__33796),
            .I(\foc.u_Park_Transform.n17171 ));
    InMux I__4157 (
            .O(N__33793),
            .I(N__33790));
    LocalMux I__4156 (
            .O(N__33790),
            .I(N__33787));
    Odrv12 I__4155 (
            .O(N__33787),
            .I(\foc.u_Park_Transform.n611 ));
    InMux I__4154 (
            .O(N__33784),
            .I(\foc.u_Park_Transform.n17172 ));
    InMux I__4153 (
            .O(N__33781),
            .I(N__33778));
    LocalMux I__4152 (
            .O(N__33778),
            .I(N__33775));
    Odrv4 I__4151 (
            .O(N__33775),
            .I(\foc.u_Park_Transform.n660 ));
    InMux I__4150 (
            .O(N__33772),
            .I(\foc.u_Park_Transform.n17173 ));
    CascadeMux I__4149 (
            .O(N__33769),
            .I(N__33766));
    InMux I__4148 (
            .O(N__33766),
            .I(N__33763));
    LocalMux I__4147 (
            .O(N__33763),
            .I(N__33760));
    Odrv4 I__4146 (
            .O(N__33760),
            .I(\foc.u_Park_Transform.n709 ));
    InMux I__4145 (
            .O(N__33757),
            .I(\foc.u_Park_Transform.n17174 ));
    InMux I__4144 (
            .O(N__33754),
            .I(bfn_11_24_0_));
    InMux I__4143 (
            .O(N__33751),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232 ));
    CascadeMux I__4142 (
            .O(N__33748),
            .I(N__33745));
    InMux I__4141 (
            .O(N__33745),
            .I(N__33742));
    LocalMux I__4140 (
            .O(N__33742),
            .I(N__33739));
    Odrv12 I__4139 (
            .O(N__33739),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO ));
    CascadeMux I__4138 (
            .O(N__33736),
            .I(N__33733));
    InMux I__4137 (
            .O(N__33733),
            .I(N__33730));
    LocalMux I__4136 (
            .O(N__33730),
            .I(N__33727));
    Odrv4 I__4135 (
            .O(N__33727),
            .I(\foc.u_Park_Transform.n72 ));
    InMux I__4134 (
            .O(N__33724),
            .I(\foc.u_Park_Transform.n17161 ));
    CascadeMux I__4133 (
            .O(N__33721),
            .I(N__33718));
    InMux I__4132 (
            .O(N__33718),
            .I(N__33715));
    LocalMux I__4131 (
            .O(N__33715),
            .I(N__33712));
    Odrv12 I__4130 (
            .O(N__33712),
            .I(\foc.u_Park_Transform.n121 ));
    InMux I__4129 (
            .O(N__33709),
            .I(\foc.u_Park_Transform.n17162 ));
    InMux I__4128 (
            .O(N__33706),
            .I(N__33703));
    LocalMux I__4127 (
            .O(N__33703),
            .I(N__33700));
    Odrv12 I__4126 (
            .O(N__33700),
            .I(\foc.u_Park_Transform.n170 ));
    InMux I__4125 (
            .O(N__33697),
            .I(\foc.u_Park_Transform.n17163 ));
    CascadeMux I__4124 (
            .O(N__33694),
            .I(N__33691));
    InMux I__4123 (
            .O(N__33691),
            .I(N__33688));
    LocalMux I__4122 (
            .O(N__33688),
            .I(N__33685));
    Odrv12 I__4121 (
            .O(N__33685),
            .I(\foc.u_Park_Transform.n219 ));
    InMux I__4120 (
            .O(N__33682),
            .I(\foc.u_Park_Transform.n17164 ));
    InMux I__4119 (
            .O(N__33679),
            .I(N__33676));
    LocalMux I__4118 (
            .O(N__33676),
            .I(N__33673));
    Odrv12 I__4117 (
            .O(N__33673),
            .I(\foc.u_Park_Transform.n268 ));
    InMux I__4116 (
            .O(N__33670),
            .I(\foc.u_Park_Transform.n17165 ));
    CascadeMux I__4115 (
            .O(N__33667),
            .I(N__33664));
    InMux I__4114 (
            .O(N__33664),
            .I(N__33661));
    LocalMux I__4113 (
            .O(N__33661),
            .I(N__33658));
    Odrv4 I__4112 (
            .O(N__33658),
            .I(\foc.u_Park_Transform.n317 ));
    InMux I__4111 (
            .O(N__33655),
            .I(\foc.u_Park_Transform.n17166 ));
    CascadeMux I__4110 (
            .O(N__33652),
            .I(N__33649));
    InMux I__4109 (
            .O(N__33649),
            .I(N__33646));
    LocalMux I__4108 (
            .O(N__33646),
            .I(N__33643));
    Odrv4 I__4107 (
            .O(N__33643),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426 ));
    InMux I__4106 (
            .O(N__33640),
            .I(N__33637));
    LocalMux I__4105 (
            .O(N__33637),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523 ));
    InMux I__4104 (
            .O(N__33634),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403 ));
    InMux I__4103 (
            .O(N__33631),
            .I(N__33628));
    LocalMux I__4102 (
            .O(N__33628),
            .I(N__33625));
    Odrv4 I__4101 (
            .O(N__33625),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526 ));
    CascadeMux I__4100 (
            .O(N__33622),
            .I(N__33619));
    InMux I__4099 (
            .O(N__33619),
            .I(N__33616));
    LocalMux I__4098 (
            .O(N__33616),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623 ));
    InMux I__4097 (
            .O(N__33613),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404 ));
    CascadeMux I__4096 (
            .O(N__33610),
            .I(N__33607));
    InMux I__4095 (
            .O(N__33607),
            .I(N__33604));
    LocalMux I__4094 (
            .O(N__33604),
            .I(N__33601));
    Odrv12 I__4093 (
            .O(N__33601),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626 ));
    InMux I__4092 (
            .O(N__33598),
            .I(N__33595));
    LocalMux I__4091 (
            .O(N__33595),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723 ));
    InMux I__4090 (
            .O(N__33592),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405 ));
    InMux I__4089 (
            .O(N__33589),
            .I(N__33586));
    LocalMux I__4088 (
            .O(N__33586),
            .I(N__33583));
    Odrv4 I__4087 (
            .O(N__33583),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726 ));
    CascadeMux I__4086 (
            .O(N__33580),
            .I(N__33577));
    InMux I__4085 (
            .O(N__33577),
            .I(N__33574));
    LocalMux I__4084 (
            .O(N__33574),
            .I(N__33571));
    Odrv4 I__4083 (
            .O(N__33571),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823 ));
    InMux I__4082 (
            .O(N__33568),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406 ));
    InMux I__4081 (
            .O(N__33565),
            .I(N__33562));
    LocalMux I__4080 (
            .O(N__33562),
            .I(N__33559));
    Odrv4 I__4079 (
            .O(N__33559),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826 ));
    InMux I__4078 (
            .O(N__33556),
            .I(N__33553));
    LocalMux I__4077 (
            .O(N__33553),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923 ));
    InMux I__4076 (
            .O(N__33550),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407 ));
    InMux I__4075 (
            .O(N__33547),
            .I(N__33544));
    LocalMux I__4074 (
            .O(N__33544),
            .I(N__33541));
    Odrv12 I__4073 (
            .O(N__33541),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926 ));
    CascadeMux I__4072 (
            .O(N__33538),
            .I(N__33535));
    InMux I__4071 (
            .O(N__33535),
            .I(N__33532));
    LocalMux I__4070 (
            .O(N__33532),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023 ));
    InMux I__4069 (
            .O(N__33529),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408 ));
    InMux I__4068 (
            .O(N__33526),
            .I(N__33523));
    LocalMux I__4067 (
            .O(N__33523),
            .I(N__33520));
    Odrv4 I__4066 (
            .O(N__33520),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026 ));
    CascadeMux I__4065 (
            .O(N__33517),
            .I(N__33510));
    CascadeMux I__4064 (
            .O(N__33516),
            .I(N__33507));
    CascadeMux I__4063 (
            .O(N__33515),
            .I(N__33504));
    CascadeMux I__4062 (
            .O(N__33514),
            .I(N__33501));
    CascadeMux I__4061 (
            .O(N__33513),
            .I(N__33497));
    InMux I__4060 (
            .O(N__33510),
            .I(N__33490));
    InMux I__4059 (
            .O(N__33507),
            .I(N__33490));
    InMux I__4058 (
            .O(N__33504),
            .I(N__33479));
    InMux I__4057 (
            .O(N__33501),
            .I(N__33479));
    InMux I__4056 (
            .O(N__33500),
            .I(N__33479));
    InMux I__4055 (
            .O(N__33497),
            .I(N__33479));
    InMux I__4054 (
            .O(N__33496),
            .I(N__33479));
    InMux I__4053 (
            .O(N__33495),
            .I(N__33476));
    LocalMux I__4052 (
            .O(N__33490),
            .I(N__33471));
    LocalMux I__4051 (
            .O(N__33479),
            .I(N__33471));
    LocalMux I__4050 (
            .O(N__33476),
            .I(N__33468));
    Span4Mux_v I__4049 (
            .O(N__33471),
            .I(N__33465));
    Span4Mux_v I__4048 (
            .O(N__33468),
            .I(N__33462));
    Odrv4 I__4047 (
            .O(N__33465),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822 ));
    Odrv4 I__4046 (
            .O(N__33462),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822 ));
    InMux I__4045 (
            .O(N__33457),
            .I(N__33454));
    LocalMux I__4044 (
            .O(N__33454),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123 ));
    InMux I__4043 (
            .O(N__33451),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409 ));
    InMux I__4042 (
            .O(N__33448),
            .I(N__33445));
    LocalMux I__4041 (
            .O(N__33445),
            .I(N__33442));
    Odrv12 I__4040 (
            .O(N__33442),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126 ));
    InMux I__4039 (
            .O(N__33439),
            .I(N__33436));
    LocalMux I__4038 (
            .O(N__33436),
            .I(N__33433));
    Odrv12 I__4037 (
            .O(N__33433),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231 ));
    CascadeMux I__4036 (
            .O(N__33430),
            .I(N__33427));
    InMux I__4035 (
            .O(N__33427),
            .I(N__33424));
    LocalMux I__4034 (
            .O(N__33424),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629 ));
    InMux I__4033 (
            .O(N__33421),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414 ));
    InMux I__4032 (
            .O(N__33418),
            .I(N__33415));
    LocalMux I__4031 (
            .O(N__33415),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729 ));
    InMux I__4030 (
            .O(N__33412),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415 ));
    InMux I__4029 (
            .O(N__33409),
            .I(N__33406));
    LocalMux I__4028 (
            .O(N__33406),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829 ));
    InMux I__4027 (
            .O(N__33403),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416 ));
    InMux I__4026 (
            .O(N__33400),
            .I(N__33397));
    LocalMux I__4025 (
            .O(N__33397),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929 ));
    InMux I__4024 (
            .O(N__33394),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417 ));
    InMux I__4023 (
            .O(N__33391),
            .I(N__33388));
    LocalMux I__4022 (
            .O(N__33388),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029 ));
    InMux I__4021 (
            .O(N__33385),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418 ));
    InMux I__4020 (
            .O(N__33382),
            .I(N__33379));
    LocalMux I__4019 (
            .O(N__33379),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129 ));
    InMux I__4018 (
            .O(N__33376),
            .I(N__33373));
    LocalMux I__4017 (
            .O(N__33373),
            .I(N__33370));
    Odrv4 I__4016 (
            .O(N__33370),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235 ));
    InMux I__4015 (
            .O(N__33367),
            .I(bfn_11_22_0_));
    InMux I__4014 (
            .O(N__33364),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236 ));
    CascadeMux I__4013 (
            .O(N__33361),
            .I(N__33358));
    InMux I__4012 (
            .O(N__33358),
            .I(N__33355));
    LocalMux I__4011 (
            .O(N__33355),
            .I(N__33352));
    Odrv4 I__4010 (
            .O(N__33352),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO ));
    CascadeMux I__4009 (
            .O(N__33349),
            .I(N__33341));
    CascadeMux I__4008 (
            .O(N__33348),
            .I(N__33338));
    CascadeMux I__4007 (
            .O(N__33347),
            .I(N__33335));
    CascadeMux I__4006 (
            .O(N__33346),
            .I(N__33332));
    CascadeMux I__4005 (
            .O(N__33345),
            .I(N__33328));
    InMux I__4004 (
            .O(N__33344),
            .I(N__33324));
    InMux I__4003 (
            .O(N__33341),
            .I(N__33319));
    InMux I__4002 (
            .O(N__33338),
            .I(N__33319));
    InMux I__4001 (
            .O(N__33335),
            .I(N__33308));
    InMux I__4000 (
            .O(N__33332),
            .I(N__33308));
    InMux I__3999 (
            .O(N__33331),
            .I(N__33308));
    InMux I__3998 (
            .O(N__33328),
            .I(N__33308));
    InMux I__3997 (
            .O(N__33327),
            .I(N__33308));
    LocalMux I__3996 (
            .O(N__33324),
            .I(N__33301));
    LocalMux I__3995 (
            .O(N__33319),
            .I(N__33301));
    LocalMux I__3994 (
            .O(N__33308),
            .I(N__33301));
    Span4Mux_v I__3993 (
            .O(N__33301),
            .I(N__33298));
    Odrv4 I__3992 (
            .O(N__33298),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825 ));
    CascadeMux I__3991 (
            .O(N__33295),
            .I(N__33292));
    InMux I__3990 (
            .O(N__33292),
            .I(N__33289));
    LocalMux I__3989 (
            .O(N__33289),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423 ));
    InMux I__3988 (
            .O(N__33286),
            .I(N__33283));
    LocalMux I__3987 (
            .O(N__33283),
            .I(N__33280));
    Odrv12 I__3986 (
            .O(N__33280),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247 ));
    CascadeMux I__3985 (
            .O(N__33277),
            .I(N__33274));
    InMux I__3984 (
            .O(N__33274),
            .I(N__33271));
    LocalMux I__3983 (
            .O(N__33271),
            .I(N__33268));
    Span4Mux_v I__3982 (
            .O(N__33268),
            .I(N__33265));
    Odrv4 I__3981 (
            .O(N__33265),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO ));
    InMux I__3980 (
            .O(N__33262),
            .I(N__33259));
    LocalMux I__3979 (
            .O(N__33259),
            .I(N__33256));
    Odrv12 I__3978 (
            .O(N__33256),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43 ));
    InMux I__3977 (
            .O(N__33253),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500 ));
    InMux I__3976 (
            .O(N__33250),
            .I(N__33247));
    LocalMux I__3975 (
            .O(N__33247),
            .I(N__33244));
    Span4Mux_v I__3974 (
            .O(N__33244),
            .I(N__33241));
    Odrv4 I__3973 (
            .O(N__33241),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251 ));
    CascadeMux I__3972 (
            .O(N__33238),
            .I(N__33235));
    InMux I__3971 (
            .O(N__33235),
            .I(N__33232));
    LocalMux I__3970 (
            .O(N__33232),
            .I(N__33229));
    Odrv12 I__3969 (
            .O(N__33229),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO ));
    InMux I__3968 (
            .O(N__33226),
            .I(N__33223));
    LocalMux I__3967 (
            .O(N__33223),
            .I(N__33220));
    Span4Mux_v I__3966 (
            .O(N__33220),
            .I(N__33217));
    Odrv4 I__3965 (
            .O(N__33217),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44 ));
    InMux I__3964 (
            .O(N__33214),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501 ));
    InMux I__3963 (
            .O(N__33211),
            .I(N__33208));
    LocalMux I__3962 (
            .O(N__33208),
            .I(N__33205));
    Span4Mux_v I__3961 (
            .O(N__33205),
            .I(N__33202));
    Span4Mux_h I__3960 (
            .O(N__33202),
            .I(N__33199));
    Odrv4 I__3959 (
            .O(N__33199),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255 ));
    CascadeMux I__3958 (
            .O(N__33196),
            .I(N__33193));
    InMux I__3957 (
            .O(N__33193),
            .I(N__33190));
    LocalMux I__3956 (
            .O(N__33190),
            .I(N__33187));
    Span4Mux_v I__3955 (
            .O(N__33187),
            .I(N__33184));
    Odrv4 I__3954 (
            .O(N__33184),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO ));
    InMux I__3953 (
            .O(N__33181),
            .I(N__33178));
    LocalMux I__3952 (
            .O(N__33178),
            .I(N__33175));
    Span4Mux_v I__3951 (
            .O(N__33175),
            .I(N__33172));
    Odrv4 I__3950 (
            .O(N__33172),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45 ));
    InMux I__3949 (
            .O(N__33169),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502 ));
    InMux I__3948 (
            .O(N__33166),
            .I(N__33163));
    LocalMux I__3947 (
            .O(N__33163),
            .I(N__33160));
    Span4Mux_h I__3946 (
            .O(N__33160),
            .I(N__33157));
    Odrv4 I__3945 (
            .O(N__33157),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259 ));
    CascadeMux I__3944 (
            .O(N__33154),
            .I(N__33151));
    InMux I__3943 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__3942 (
            .O(N__33148),
            .I(N__33145));
    Span4Mux_v I__3941 (
            .O(N__33145),
            .I(N__33142));
    Span4Mux_v I__3940 (
            .O(N__33142),
            .I(N__33139));
    Odrv4 I__3939 (
            .O(N__33139),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO ));
    InMux I__3938 (
            .O(N__33136),
            .I(N__33133));
    LocalMux I__3937 (
            .O(N__33133),
            .I(N__33130));
    Span4Mux_v I__3936 (
            .O(N__33130),
            .I(N__33127));
    Odrv4 I__3935 (
            .O(N__33127),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46 ));
    InMux I__3934 (
            .O(N__33124),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503 ));
    InMux I__3933 (
            .O(N__33121),
            .I(N__33118));
    LocalMux I__3932 (
            .O(N__33118),
            .I(N__33115));
    Span4Mux_v I__3931 (
            .O(N__33115),
            .I(N__33112));
    Span4Mux_v I__3930 (
            .O(N__33112),
            .I(N__33109));
    Odrv4 I__3929 (
            .O(N__33109),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263 ));
    InMux I__3928 (
            .O(N__33106),
            .I(N__33103));
    LocalMux I__3927 (
            .O(N__33103),
            .I(N__33100));
    Span4Mux_h I__3926 (
            .O(N__33100),
            .I(N__33097));
    Odrv4 I__3925 (
            .O(N__33097),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO ));
    InMux I__3924 (
            .O(N__33094),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504 ));
    InMux I__3923 (
            .O(N__33091),
            .I(N__33088));
    LocalMux I__3922 (
            .O(N__33088),
            .I(N__33085));
    Span4Mux_v I__3921 (
            .O(N__33085),
            .I(N__33082));
    Odrv4 I__3920 (
            .O(N__33082),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47 ));
    InMux I__3919 (
            .O(N__33079),
            .I(N__33076));
    LocalMux I__3918 (
            .O(N__33076),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329 ));
    CascadeMux I__3917 (
            .O(N__33073),
            .I(N__33070));
    InMux I__3916 (
            .O(N__33070),
            .I(N__33067));
    LocalMux I__3915 (
            .O(N__33067),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429 ));
    InMux I__3914 (
            .O(N__33064),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412 ));
    InMux I__3913 (
            .O(N__33061),
            .I(N__33058));
    LocalMux I__3912 (
            .O(N__33058),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529 ));
    InMux I__3911 (
            .O(N__33055),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413 ));
    CascadeMux I__3910 (
            .O(N__33052),
            .I(N__33049));
    InMux I__3909 (
            .O(N__33049),
            .I(N__33046));
    LocalMux I__3908 (
            .O(N__33046),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO ));
    InMux I__3907 (
            .O(N__33043),
            .I(N__33040));
    LocalMux I__3906 (
            .O(N__33040),
            .I(N__33037));
    Odrv12 I__3905 (
            .O(N__33037),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35 ));
    InMux I__3904 (
            .O(N__33034),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492 ));
    InMux I__3903 (
            .O(N__33031),
            .I(N__33028));
    LocalMux I__3902 (
            .O(N__33028),
            .I(N__33025));
    Odrv12 I__3901 (
            .O(N__33025),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36 ));
    InMux I__3900 (
            .O(N__33022),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493 ));
    InMux I__3899 (
            .O(N__33019),
            .I(N__33016));
    LocalMux I__3898 (
            .O(N__33016),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223 ));
    InMux I__3897 (
            .O(N__33013),
            .I(N__33010));
    LocalMux I__3896 (
            .O(N__33010),
            .I(N__33007));
    Odrv12 I__3895 (
            .O(N__33007),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37 ));
    InMux I__3894 (
            .O(N__33004),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494 ));
    InMux I__3893 (
            .O(N__33001),
            .I(N__32998));
    LocalMux I__3892 (
            .O(N__32998),
            .I(N__32995));
    Span4Mux_v I__3891 (
            .O(N__32995),
            .I(N__32992));
    Odrv4 I__3890 (
            .O(N__32992),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227 ));
    CascadeMux I__3889 (
            .O(N__32989),
            .I(N__32986));
    InMux I__3888 (
            .O(N__32986),
            .I(N__32983));
    LocalMux I__3887 (
            .O(N__32983),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO ));
    InMux I__3886 (
            .O(N__32980),
            .I(N__32977));
    LocalMux I__3885 (
            .O(N__32977),
            .I(N__32974));
    Span4Mux_v I__3884 (
            .O(N__32974),
            .I(N__32971));
    Odrv4 I__3883 (
            .O(N__32971),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38 ));
    InMux I__3882 (
            .O(N__32968),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495 ));
    CascadeMux I__3881 (
            .O(N__32965),
            .I(N__32962));
    InMux I__3880 (
            .O(N__32962),
            .I(N__32959));
    LocalMux I__3879 (
            .O(N__32959),
            .I(N__32956));
    Span4Mux_v I__3878 (
            .O(N__32956),
            .I(N__32953));
    Odrv4 I__3877 (
            .O(N__32953),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO ));
    InMux I__3876 (
            .O(N__32950),
            .I(N__32947));
    LocalMux I__3875 (
            .O(N__32947),
            .I(N__32944));
    Span4Mux_v I__3874 (
            .O(N__32944),
            .I(N__32941));
    Odrv4 I__3873 (
            .O(N__32941),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39 ));
    InMux I__3872 (
            .O(N__32938),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496 ));
    InMux I__3871 (
            .O(N__32935),
            .I(N__32932));
    LocalMux I__3870 (
            .O(N__32932),
            .I(N__32929));
    Odrv12 I__3869 (
            .O(N__32929),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40 ));
    InMux I__3868 (
            .O(N__32926),
            .I(bfn_11_20_0_));
    InMux I__3867 (
            .O(N__32923),
            .I(N__32920));
    LocalMux I__3866 (
            .O(N__32920),
            .I(N__32917));
    Odrv4 I__3865 (
            .O(N__32917),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239 ));
    InMux I__3864 (
            .O(N__32914),
            .I(N__32911));
    LocalMux I__3863 (
            .O(N__32911),
            .I(N__32908));
    Odrv12 I__3862 (
            .O(N__32908),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41 ));
    InMux I__3861 (
            .O(N__32905),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498 ));
    InMux I__3860 (
            .O(N__32902),
            .I(N__32899));
    LocalMux I__3859 (
            .O(N__32899),
            .I(N__32896));
    Span4Mux_v I__3858 (
            .O(N__32896),
            .I(N__32893));
    Odrv4 I__3857 (
            .O(N__32893),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243 ));
    CascadeMux I__3856 (
            .O(N__32890),
            .I(N__32887));
    InMux I__3855 (
            .O(N__32887),
            .I(N__32884));
    LocalMux I__3854 (
            .O(N__32884),
            .I(N__32881));
    Odrv4 I__3853 (
            .O(N__32881),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO ));
    InMux I__3852 (
            .O(N__32878),
            .I(N__32875));
    LocalMux I__3851 (
            .O(N__32875),
            .I(N__32872));
    Odrv12 I__3850 (
            .O(N__32872),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42 ));
    InMux I__3849 (
            .O(N__32869),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499 ));
    InMux I__3848 (
            .O(N__32866),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363 ));
    CascadeMux I__3847 (
            .O(N__32863),
            .I(N__32857));
    CascadeMux I__3846 (
            .O(N__32862),
            .I(N__32853));
    CascadeMux I__3845 (
            .O(N__32861),
            .I(N__32849));
    InMux I__3844 (
            .O(N__32860),
            .I(N__32833));
    InMux I__3843 (
            .O(N__32857),
            .I(N__32833));
    InMux I__3842 (
            .O(N__32856),
            .I(N__32833));
    InMux I__3841 (
            .O(N__32853),
            .I(N__32833));
    InMux I__3840 (
            .O(N__32852),
            .I(N__32833));
    InMux I__3839 (
            .O(N__32849),
            .I(N__32833));
    InMux I__3838 (
            .O(N__32848),
            .I(N__32833));
    LocalMux I__3837 (
            .O(N__32833),
            .I(N__32830));
    Span4Mux_v I__3836 (
            .O(N__32830),
            .I(N__32827));
    Odrv4 I__3835 (
            .O(N__32827),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807 ));
    InMux I__3834 (
            .O(N__32824),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364 ));
    InMux I__3833 (
            .O(N__32821),
            .I(bfn_11_18_0_));
    InMux I__3832 (
            .O(N__32818),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212 ));
    InMux I__3831 (
            .O(N__32815),
            .I(N__32812));
    LocalMux I__3830 (
            .O(N__32812),
            .I(N__32809));
    Odrv4 I__3829 (
            .O(N__32809),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008 ));
    CascadeMux I__3828 (
            .O(N__32806),
            .I(N__32801));
    CascadeMux I__3827 (
            .O(N__32805),
            .I(N__32793));
    CascadeMux I__3826 (
            .O(N__32804),
            .I(N__32790));
    InMux I__3825 (
            .O(N__32801),
            .I(N__32787));
    CascadeMux I__3824 (
            .O(N__32800),
            .I(N__32784));
    CascadeMux I__3823 (
            .O(N__32799),
            .I(N__32780));
    InMux I__3822 (
            .O(N__32798),
            .I(N__32777));
    CascadeMux I__3821 (
            .O(N__32797),
            .I(N__32774));
    CascadeMux I__3820 (
            .O(N__32796),
            .I(N__32771));
    InMux I__3819 (
            .O(N__32793),
            .I(N__32767));
    InMux I__3818 (
            .O(N__32790),
            .I(N__32762));
    LocalMux I__3817 (
            .O(N__32787),
            .I(N__32759));
    InMux I__3816 (
            .O(N__32784),
            .I(N__32756));
    InMux I__3815 (
            .O(N__32783),
            .I(N__32751));
    InMux I__3814 (
            .O(N__32780),
            .I(N__32751));
    LocalMux I__3813 (
            .O(N__32777),
            .I(N__32748));
    InMux I__3812 (
            .O(N__32774),
            .I(N__32745));
    InMux I__3811 (
            .O(N__32771),
            .I(N__32742));
    CascadeMux I__3810 (
            .O(N__32770),
            .I(N__32739));
    LocalMux I__3809 (
            .O(N__32767),
            .I(N__32735));
    CascadeMux I__3808 (
            .O(N__32766),
            .I(N__32732));
    CascadeMux I__3807 (
            .O(N__32765),
            .I(N__32729));
    LocalMux I__3806 (
            .O(N__32762),
            .I(N__32725));
    Span4Mux_v I__3805 (
            .O(N__32759),
            .I(N__32714));
    LocalMux I__3804 (
            .O(N__32756),
            .I(N__32714));
    LocalMux I__3803 (
            .O(N__32751),
            .I(N__32714));
    Span4Mux_h I__3802 (
            .O(N__32748),
            .I(N__32714));
    LocalMux I__3801 (
            .O(N__32745),
            .I(N__32714));
    LocalMux I__3800 (
            .O(N__32742),
            .I(N__32711));
    InMux I__3799 (
            .O(N__32739),
            .I(N__32708));
    CascadeMux I__3798 (
            .O(N__32738),
            .I(N__32705));
    Span4Mux_v I__3797 (
            .O(N__32735),
            .I(N__32702));
    InMux I__3796 (
            .O(N__32732),
            .I(N__32697));
    InMux I__3795 (
            .O(N__32729),
            .I(N__32697));
    InMux I__3794 (
            .O(N__32728),
            .I(N__32694));
    Span4Mux_v I__3793 (
            .O(N__32725),
            .I(N__32688));
    Span4Mux_v I__3792 (
            .O(N__32714),
            .I(N__32688));
    Span4Mux_h I__3791 (
            .O(N__32711),
            .I(N__32683));
    LocalMux I__3790 (
            .O(N__32708),
            .I(N__32683));
    InMux I__3789 (
            .O(N__32705),
            .I(N__32680));
    Span4Mux_v I__3788 (
            .O(N__32702),
            .I(N__32673));
    LocalMux I__3787 (
            .O(N__32697),
            .I(N__32673));
    LocalMux I__3786 (
            .O(N__32694),
            .I(N__32673));
    InMux I__3785 (
            .O(N__32693),
            .I(N__32670));
    Odrv4 I__3784 (
            .O(N__32688),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ));
    Odrv4 I__3783 (
            .O(N__32683),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ));
    LocalMux I__3782 (
            .O(N__32680),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ));
    Odrv4 I__3781 (
            .O(N__32673),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ));
    LocalMux I__3780 (
            .O(N__32670),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ));
    InMux I__3779 (
            .O(N__32659),
            .I(N__32656));
    LocalMux I__3778 (
            .O(N__32656),
            .I(N__32653));
    Odrv4 I__3777 (
            .O(N__32653),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108 ));
    InMux I__3776 (
            .O(N__32650),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490 ));
    InMux I__3775 (
            .O(N__32647),
            .I(N__32644));
    LocalMux I__3774 (
            .O(N__32644),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211 ));
    InMux I__3773 (
            .O(N__32641),
            .I(N__32638));
    LocalMux I__3772 (
            .O(N__32638),
            .I(N__32635));
    Odrv12 I__3771 (
            .O(N__32635),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34 ));
    InMux I__3770 (
            .O(N__32632),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491 ));
    InMux I__3769 (
            .O(N__32629),
            .I(\foc.u_Park_Transform.n16959 ));
    InMux I__3768 (
            .O(N__32626),
            .I(\foc.u_Park_Transform.n16960 ));
    InMux I__3767 (
            .O(N__32623),
            .I(N__32620));
    LocalMux I__3766 (
            .O(N__32620),
            .I(N__32616));
    InMux I__3765 (
            .O(N__32619),
            .I(N__32613));
    Odrv4 I__3764 (
            .O(N__32616),
            .I(\foc.u_Park_Transform.n769 ));
    LocalMux I__3763 (
            .O(N__32613),
            .I(\foc.u_Park_Transform.n769 ));
    CascadeMux I__3762 (
            .O(N__32608),
            .I(N__32604));
    CascadeMux I__3761 (
            .O(N__32607),
            .I(N__32601));
    InMux I__3760 (
            .O(N__32604),
            .I(N__32597));
    InMux I__3759 (
            .O(N__32601),
            .I(N__32592));
    InMux I__3758 (
            .O(N__32600),
            .I(N__32592));
    LocalMux I__3757 (
            .O(N__32597),
            .I(N__32587));
    LocalMux I__3756 (
            .O(N__32592),
            .I(N__32587));
    Odrv12 I__3755 (
            .O(N__32587),
            .I(\foc.u_Park_Transform.n617 ));
    InMux I__3754 (
            .O(N__32584),
            .I(\foc.u_Park_Transform.n16961 ));
    InMux I__3753 (
            .O(N__32581),
            .I(\foc.u_Park_Transform.n771 ));
    CascadeMux I__3752 (
            .O(N__32578),
            .I(N__32575));
    InMux I__3751 (
            .O(N__32575),
            .I(N__32572));
    LocalMux I__3750 (
            .O(N__32572),
            .I(N__32569));
    Odrv12 I__3749 (
            .O(N__32569),
            .I(\foc.u_Park_Transform.n176_adj_2104 ));
    InMux I__3748 (
            .O(N__32566),
            .I(\foc.u_Park_Transform.n16950 ));
    CascadeMux I__3747 (
            .O(N__32563),
            .I(N__32560));
    InMux I__3746 (
            .O(N__32560),
            .I(N__32557));
    LocalMux I__3745 (
            .O(N__32557),
            .I(N__32554));
    Odrv12 I__3744 (
            .O(N__32554),
            .I(\foc.u_Park_Transform.n225_adj_2075 ));
    InMux I__3743 (
            .O(N__32551),
            .I(\foc.u_Park_Transform.n16951 ));
    CascadeMux I__3742 (
            .O(N__32548),
            .I(N__32545));
    InMux I__3741 (
            .O(N__32545),
            .I(N__32542));
    LocalMux I__3740 (
            .O(N__32542),
            .I(N__32539));
    Odrv4 I__3739 (
            .O(N__32539),
            .I(\foc.u_Park_Transform.n274_adj_2058 ));
    InMux I__3738 (
            .O(N__32536),
            .I(\foc.u_Park_Transform.n16952 ));
    CascadeMux I__3737 (
            .O(N__32533),
            .I(N__32530));
    InMux I__3736 (
            .O(N__32530),
            .I(N__32527));
    LocalMux I__3735 (
            .O(N__32527),
            .I(N__32524));
    Odrv12 I__3734 (
            .O(N__32524),
            .I(\foc.u_Park_Transform.n323_adj_2057 ));
    InMux I__3733 (
            .O(N__32521),
            .I(\foc.u_Park_Transform.n16953 ));
    CascadeMux I__3732 (
            .O(N__32518),
            .I(N__32515));
    InMux I__3731 (
            .O(N__32515),
            .I(N__32512));
    LocalMux I__3730 (
            .O(N__32512),
            .I(N__32509));
    Odrv4 I__3729 (
            .O(N__32509),
            .I(\foc.u_Park_Transform.n372_adj_2042 ));
    InMux I__3728 (
            .O(N__32506),
            .I(\foc.u_Park_Transform.n16954 ));
    CascadeMux I__3727 (
            .O(N__32503),
            .I(N__32500));
    InMux I__3726 (
            .O(N__32500),
            .I(N__32497));
    LocalMux I__3725 (
            .O(N__32497),
            .I(N__32494));
    Span4Mux_v I__3724 (
            .O(N__32494),
            .I(N__32491));
    Odrv4 I__3723 (
            .O(N__32491),
            .I(\foc.u_Park_Transform.n421 ));
    InMux I__3722 (
            .O(N__32488),
            .I(bfn_11_16_0_));
    InMux I__3721 (
            .O(N__32485),
            .I(N__32482));
    LocalMux I__3720 (
            .O(N__32482),
            .I(N__32479));
    Odrv4 I__3719 (
            .O(N__32479),
            .I(\foc.u_Park_Transform.n470 ));
    InMux I__3718 (
            .O(N__32476),
            .I(\foc.u_Park_Transform.n16956 ));
    CascadeMux I__3717 (
            .O(N__32473),
            .I(N__32470));
    InMux I__3716 (
            .O(N__32470),
            .I(N__32467));
    LocalMux I__3715 (
            .O(N__32467),
            .I(N__32464));
    Odrv4 I__3714 (
            .O(N__32464),
            .I(\foc.u_Park_Transform.n519 ));
    InMux I__3713 (
            .O(N__32461),
            .I(\foc.u_Park_Transform.n16957 ));
    InMux I__3712 (
            .O(N__32458),
            .I(N__32455));
    LocalMux I__3711 (
            .O(N__32455),
            .I(N__32452));
    Odrv12 I__3710 (
            .O(N__32452),
            .I(\foc.u_Park_Transform.n568 ));
    InMux I__3709 (
            .O(N__32449),
            .I(\foc.u_Park_Transform.n16958 ));
    InMux I__3708 (
            .O(N__32446),
            .I(N__32440));
    InMux I__3707 (
            .O(N__32445),
            .I(N__32440));
    LocalMux I__3706 (
            .O(N__32440),
            .I(N__32437));
    Odrv12 I__3705 (
            .O(N__32437),
            .I(\foc.Look_Up_Table_out1_1_11 ));
    InMux I__3704 (
            .O(N__32434),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952 ));
    InMux I__3703 (
            .O(N__32431),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953 ));
    InMux I__3702 (
            .O(N__32428),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954 ));
    InMux I__3701 (
            .O(N__32425),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955 ));
    InMux I__3700 (
            .O(N__32422),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956 ));
    InMux I__3699 (
            .O(N__32419),
            .I(N__32416));
    LocalMux I__3698 (
            .O(N__32416),
            .I(N__32412));
    InMux I__3697 (
            .O(N__32415),
            .I(N__32409));
    Odrv4 I__3696 (
            .O(N__32412),
            .I(\foc.Look_Up_Table_out1_1_12 ));
    LocalMux I__3695 (
            .O(N__32409),
            .I(\foc.Look_Up_Table_out1_1_12 ));
    InMux I__3694 (
            .O(N__32404),
            .I(N__32401));
    LocalMux I__3693 (
            .O(N__32401),
            .I(N__32398));
    Span4Mux_v I__3692 (
            .O(N__32398),
            .I(N__32394));
    InMux I__3691 (
            .O(N__32397),
            .I(N__32391));
    Odrv4 I__3690 (
            .O(N__32394),
            .I(\foc.u_Park_Transform.n785 ));
    LocalMux I__3689 (
            .O(N__32391),
            .I(\foc.u_Park_Transform.n785 ));
    CascadeMux I__3688 (
            .O(N__32386),
            .I(N__32377));
    CascadeMux I__3687 (
            .O(N__32385),
            .I(N__32373));
    CascadeMux I__3686 (
            .O(N__32384),
            .I(N__32360));
    InMux I__3685 (
            .O(N__32383),
            .I(N__32353));
    InMux I__3684 (
            .O(N__32382),
            .I(N__32353));
    InMux I__3683 (
            .O(N__32381),
            .I(N__32353));
    InMux I__3682 (
            .O(N__32380),
            .I(N__32343));
    InMux I__3681 (
            .O(N__32377),
            .I(N__32343));
    InMux I__3680 (
            .O(N__32376),
            .I(N__32343));
    InMux I__3679 (
            .O(N__32373),
            .I(N__32343));
    CascadeMux I__3678 (
            .O(N__32372),
            .I(N__32340));
    CascadeMux I__3677 (
            .O(N__32371),
            .I(N__32336));
    CascadeMux I__3676 (
            .O(N__32370),
            .I(N__32332));
    CascadeMux I__3675 (
            .O(N__32369),
            .I(N__32327));
    CascadeMux I__3674 (
            .O(N__32368),
            .I(N__32324));
    CascadeMux I__3673 (
            .O(N__32367),
            .I(N__32320));
    InMux I__3672 (
            .O(N__32366),
            .I(N__32307));
    InMux I__3671 (
            .O(N__32365),
            .I(N__32307));
    InMux I__3670 (
            .O(N__32364),
            .I(N__32307));
    InMux I__3669 (
            .O(N__32363),
            .I(N__32307));
    InMux I__3668 (
            .O(N__32360),
            .I(N__32307));
    LocalMux I__3667 (
            .O(N__32353),
            .I(N__32304));
    InMux I__3666 (
            .O(N__32352),
            .I(N__32301));
    LocalMux I__3665 (
            .O(N__32343),
            .I(N__32298));
    InMux I__3664 (
            .O(N__32340),
            .I(N__32285));
    InMux I__3663 (
            .O(N__32339),
            .I(N__32285));
    InMux I__3662 (
            .O(N__32336),
            .I(N__32285));
    InMux I__3661 (
            .O(N__32335),
            .I(N__32285));
    InMux I__3660 (
            .O(N__32332),
            .I(N__32285));
    InMux I__3659 (
            .O(N__32331),
            .I(N__32285));
    InMux I__3658 (
            .O(N__32330),
            .I(N__32280));
    InMux I__3657 (
            .O(N__32327),
            .I(N__32280));
    InMux I__3656 (
            .O(N__32324),
            .I(N__32271));
    InMux I__3655 (
            .O(N__32323),
            .I(N__32271));
    InMux I__3654 (
            .O(N__32320),
            .I(N__32271));
    InMux I__3653 (
            .O(N__32319),
            .I(N__32271));
    InMux I__3652 (
            .O(N__32318),
            .I(N__32268));
    LocalMux I__3651 (
            .O(N__32307),
            .I(N__32265));
    Span4Mux_h I__3650 (
            .O(N__32304),
            .I(N__32260));
    LocalMux I__3649 (
            .O(N__32301),
            .I(N__32260));
    Span4Mux_v I__3648 (
            .O(N__32298),
            .I(N__32249));
    LocalMux I__3647 (
            .O(N__32285),
            .I(N__32249));
    LocalMux I__3646 (
            .O(N__32280),
            .I(N__32249));
    LocalMux I__3645 (
            .O(N__32271),
            .I(N__32249));
    LocalMux I__3644 (
            .O(N__32268),
            .I(N__32249));
    Odrv4 I__3643 (
            .O(N__32265),
            .I(\foc.u_Park_Transform.n616 ));
    Odrv4 I__3642 (
            .O(N__32260),
            .I(\foc.u_Park_Transform.n616 ));
    Odrv4 I__3641 (
            .O(N__32249),
            .I(\foc.u_Park_Transform.n616 ));
    InMux I__3640 (
            .O(N__32242),
            .I(N__32239));
    LocalMux I__3639 (
            .O(N__32239),
            .I(N__32236));
    Odrv4 I__3638 (
            .O(N__32236),
            .I(\foc.u_Park_Transform.n78_adj_2145 ));
    InMux I__3637 (
            .O(N__32233),
            .I(\foc.u_Park_Transform.n16948 ));
    CascadeMux I__3636 (
            .O(N__32230),
            .I(N__32227));
    InMux I__3635 (
            .O(N__32227),
            .I(N__32224));
    LocalMux I__3634 (
            .O(N__32224),
            .I(N__32221));
    Odrv4 I__3633 (
            .O(N__32221),
            .I(\foc.u_Park_Transform.n127_adj_2119 ));
    InMux I__3632 (
            .O(N__32218),
            .I(\foc.u_Park_Transform.n16949 ));
    InMux I__3631 (
            .O(N__32215),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944 ));
    InMux I__3630 (
            .O(N__32212),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945 ));
    InMux I__3629 (
            .O(N__32209),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946 ));
    InMux I__3628 (
            .O(N__32206),
            .I(N__32200));
    InMux I__3627 (
            .O(N__32205),
            .I(N__32200));
    LocalMux I__3626 (
            .O(N__32200),
            .I(\foc.Look_Up_Table_out1_1_6 ));
    InMux I__3625 (
            .O(N__32197),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947 ));
    InMux I__3624 (
            .O(N__32194),
            .I(N__32188));
    InMux I__3623 (
            .O(N__32193),
            .I(N__32188));
    LocalMux I__3622 (
            .O(N__32188),
            .I(\foc.Look_Up_Table_out1_1_7 ));
    InMux I__3621 (
            .O(N__32185),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948 ));
    InMux I__3620 (
            .O(N__32182),
            .I(N__32176));
    InMux I__3619 (
            .O(N__32181),
            .I(N__32176));
    LocalMux I__3618 (
            .O(N__32176),
            .I(\foc.Look_Up_Table_out1_1_8 ));
    InMux I__3617 (
            .O(N__32173),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949 ));
    InMux I__3616 (
            .O(N__32170),
            .I(N__32164));
    InMux I__3615 (
            .O(N__32169),
            .I(N__32164));
    LocalMux I__3614 (
            .O(N__32164),
            .I(\foc.Look_Up_Table_out1_1_9 ));
    InMux I__3613 (
            .O(N__32161),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950 ));
    InMux I__3612 (
            .O(N__32158),
            .I(N__32152));
    InMux I__3611 (
            .O(N__32157),
            .I(N__32152));
    LocalMux I__3610 (
            .O(N__32152),
            .I(N__32149));
    Odrv4 I__3609 (
            .O(N__32149),
            .I(\foc.Look_Up_Table_out1_1_10 ));
    InMux I__3608 (
            .O(N__32146),
            .I(bfn_11_14_0_));
    InMux I__3607 (
            .O(N__32143),
            .I(\foc.u_Park_Transform.n787_adj_2149 ));
    CascadeMux I__3606 (
            .O(N__32140),
            .I(N__32137));
    InMux I__3605 (
            .O(N__32137),
            .I(N__32126));
    InMux I__3604 (
            .O(N__32136),
            .I(N__32126));
    InMux I__3603 (
            .O(N__32135),
            .I(N__32126));
    CascadeMux I__3602 (
            .O(N__32134),
            .I(N__32121));
    InMux I__3601 (
            .O(N__32133),
            .I(N__32118));
    LocalMux I__3600 (
            .O(N__32126),
            .I(N__32110));
    InMux I__3599 (
            .O(N__32125),
            .I(N__32103));
    InMux I__3598 (
            .O(N__32124),
            .I(N__32103));
    InMux I__3597 (
            .O(N__32121),
            .I(N__32103));
    LocalMux I__3596 (
            .O(N__32118),
            .I(N__32100));
    InMux I__3595 (
            .O(N__32117),
            .I(N__32097));
    CascadeMux I__3594 (
            .O(N__32116),
            .I(N__32094));
    CascadeMux I__3593 (
            .O(N__32115),
            .I(N__32090));
    CascadeMux I__3592 (
            .O(N__32114),
            .I(N__32086));
    CascadeMux I__3591 (
            .O(N__32113),
            .I(N__32083));
    Span4Mux_h I__3590 (
            .O(N__32110),
            .I(N__32078));
    LocalMux I__3589 (
            .O(N__32103),
            .I(N__32078));
    Span4Mux_v I__3588 (
            .O(N__32100),
            .I(N__32073));
    LocalMux I__3587 (
            .O(N__32097),
            .I(N__32073));
    InMux I__3586 (
            .O(N__32094),
            .I(N__32066));
    InMux I__3585 (
            .O(N__32093),
            .I(N__32066));
    InMux I__3584 (
            .O(N__32090),
            .I(N__32066));
    InMux I__3583 (
            .O(N__32089),
            .I(N__32059));
    InMux I__3582 (
            .O(N__32086),
            .I(N__32059));
    InMux I__3581 (
            .O(N__32083),
            .I(N__32059));
    Odrv4 I__3580 (
            .O(N__32078),
            .I(\foc.u_Park_Transform.n625 ));
    Odrv4 I__3579 (
            .O(N__32073),
            .I(\foc.u_Park_Transform.n625 ));
    LocalMux I__3578 (
            .O(N__32066),
            .I(\foc.u_Park_Transform.n625 ));
    LocalMux I__3577 (
            .O(N__32059),
            .I(\foc.u_Park_Transform.n625 ));
    CascadeMux I__3576 (
            .O(N__32050),
            .I(n21486_cascade_));
    CascadeMux I__3575 (
            .O(N__32047),
            .I(N__32044));
    InMux I__3574 (
            .O(N__32044),
            .I(N__32041));
    LocalMux I__3573 (
            .O(N__32041),
            .I(N__32037));
    InMux I__3572 (
            .O(N__32040),
            .I(N__32034));
    Odrv4 I__3571 (
            .O(N__32037),
            .I(n139));
    LocalMux I__3570 (
            .O(N__32034),
            .I(n139));
    CascadeMux I__3569 (
            .O(N__32029),
            .I(N__32026));
    InMux I__3568 (
            .O(N__32026),
            .I(N__32023));
    LocalMux I__3567 (
            .O(N__32023),
            .I(N__32019));
    InMux I__3566 (
            .O(N__32022),
            .I(N__32016));
    Odrv4 I__3565 (
            .O(N__32019),
            .I(\foc.u_Park_Transform.n90 ));
    LocalMux I__3564 (
            .O(N__32016),
            .I(\foc.u_Park_Transform.n90 ));
    InMux I__3563 (
            .O(N__32011),
            .I(N__32008));
    LocalMux I__3562 (
            .O(N__32008),
            .I(N__32005));
    Span4Mux_v I__3561 (
            .O(N__32005),
            .I(N__32001));
    InMux I__3560 (
            .O(N__32004),
            .I(N__31998));
    Odrv4 I__3559 (
            .O(N__32001),
            .I(\foc.u_Park_Transform.n781 ));
    LocalMux I__3558 (
            .O(N__31998),
            .I(\foc.u_Park_Transform.n781 ));
    CascadeMux I__3557 (
            .O(N__31993),
            .I(N__31990));
    InMux I__3556 (
            .O(N__31990),
            .I(N__31987));
    LocalMux I__3555 (
            .O(N__31987),
            .I(N__31984));
    Odrv4 I__3554 (
            .O(N__31984),
            .I(\foc.u_Park_Transform.n87_adj_2138 ));
    CascadeMux I__3553 (
            .O(N__31981),
            .I(N__31978));
    InMux I__3552 (
            .O(N__31978),
            .I(N__31975));
    LocalMux I__3551 (
            .O(N__31975),
            .I(N__31972));
    Odrv4 I__3550 (
            .O(N__31972),
            .I(\foc.u_Park_Transform.n136_adj_2127 ));
    InMux I__3549 (
            .O(N__31969),
            .I(\foc.u_Park_Transform.n17980 ));
    InMux I__3548 (
            .O(N__31966),
            .I(N__31963));
    LocalMux I__3547 (
            .O(N__31963),
            .I(N__31960));
    Odrv4 I__3546 (
            .O(N__31960),
            .I(\foc.u_Park_Transform.n185_adj_2126 ));
    InMux I__3545 (
            .O(N__31957),
            .I(\foc.u_Park_Transform.n17981 ));
    CascadeMux I__3544 (
            .O(N__31954),
            .I(N__31951));
    InMux I__3543 (
            .O(N__31951),
            .I(N__31948));
    LocalMux I__3542 (
            .O(N__31948),
            .I(N__31945));
    Odrv4 I__3541 (
            .O(N__31945),
            .I(\foc.u_Park_Transform.n234_adj_2125 ));
    InMux I__3540 (
            .O(N__31942),
            .I(\foc.u_Park_Transform.n17982 ));
    InMux I__3539 (
            .O(N__31939),
            .I(N__31936));
    LocalMux I__3538 (
            .O(N__31936),
            .I(N__31933));
    Odrv4 I__3537 (
            .O(N__31933),
            .I(\foc.u_Park_Transform.n283_adj_2122 ));
    InMux I__3536 (
            .O(N__31930),
            .I(\foc.u_Park_Transform.n17983 ));
    CascadeMux I__3535 (
            .O(N__31927),
            .I(N__31923));
    InMux I__3534 (
            .O(N__31926),
            .I(N__31917));
    InMux I__3533 (
            .O(N__31923),
            .I(N__31917));
    CascadeMux I__3532 (
            .O(N__31922),
            .I(N__31914));
    LocalMux I__3531 (
            .O(N__31917),
            .I(N__31911));
    InMux I__3530 (
            .O(N__31914),
            .I(N__31908));
    Odrv4 I__3529 (
            .O(N__31911),
            .I(\foc.u_Park_Transform.n332_adj_2110 ));
    LocalMux I__3528 (
            .O(N__31908),
            .I(\foc.u_Park_Transform.n332_adj_2110 ));
    InMux I__3527 (
            .O(N__31903),
            .I(\foc.u_Park_Transform.n17984 ));
    InMux I__3526 (
            .O(N__31900),
            .I(\foc.u_Park_Transform.n17985 ));
    InMux I__3525 (
            .O(N__31897),
            .I(N__31894));
    LocalMux I__3524 (
            .O(N__31894),
            .I(N__31891));
    Odrv4 I__3523 (
            .O(N__31891),
            .I(\foc.u_Park_Transform.n182_adj_2094 ));
    InMux I__3522 (
            .O(N__31888),
            .I(\foc.u_Park_Transform.n17099 ));
    CascadeMux I__3521 (
            .O(N__31885),
            .I(N__31882));
    InMux I__3520 (
            .O(N__31882),
            .I(N__31879));
    LocalMux I__3519 (
            .O(N__31879),
            .I(N__31876));
    Odrv4 I__3518 (
            .O(N__31876),
            .I(\foc.u_Park_Transform.n231_adj_2089 ));
    InMux I__3517 (
            .O(N__31873),
            .I(\foc.u_Park_Transform.n17100 ));
    InMux I__3516 (
            .O(N__31870),
            .I(N__31867));
    LocalMux I__3515 (
            .O(N__31867),
            .I(N__31864));
    Span4Mux_v I__3514 (
            .O(N__31864),
            .I(N__31861));
    Odrv4 I__3513 (
            .O(N__31861),
            .I(\foc.u_Park_Transform.n280_adj_2087 ));
    InMux I__3512 (
            .O(N__31858),
            .I(\foc.u_Park_Transform.n17101 ));
    CascadeMux I__3511 (
            .O(N__31855),
            .I(N__31852));
    InMux I__3510 (
            .O(N__31852),
            .I(N__31849));
    LocalMux I__3509 (
            .O(N__31849),
            .I(N__31846));
    Span4Mux_v I__3508 (
            .O(N__31846),
            .I(N__31843));
    Odrv4 I__3507 (
            .O(N__31843),
            .I(\foc.u_Park_Transform.n329_adj_2080 ));
    InMux I__3506 (
            .O(N__31840),
            .I(\foc.u_Park_Transform.n17102 ));
    InMux I__3505 (
            .O(N__31837),
            .I(N__31834));
    LocalMux I__3504 (
            .O(N__31834),
            .I(N__31831));
    Odrv12 I__3503 (
            .O(N__31831),
            .I(\foc.u_Park_Transform.n378_adj_2078 ));
    InMux I__3502 (
            .O(N__31828),
            .I(\foc.u_Park_Transform.n17103 ));
    CascadeMux I__3501 (
            .O(N__31825),
            .I(N__31821));
    CascadeMux I__3500 (
            .O(N__31824),
            .I(N__31817));
    InMux I__3499 (
            .O(N__31821),
            .I(N__31810));
    InMux I__3498 (
            .O(N__31820),
            .I(N__31810));
    InMux I__3497 (
            .O(N__31817),
            .I(N__31810));
    LocalMux I__3496 (
            .O(N__31810),
            .I(N__31807));
    Span4Mux_h I__3495 (
            .O(N__31807),
            .I(N__31804));
    Odrv4 I__3494 (
            .O(N__31804),
            .I(\foc.u_Park_Transform.n427_adj_2069 ));
    InMux I__3493 (
            .O(N__31801),
            .I(\foc.u_Park_Transform.n17104 ));
    InMux I__3492 (
            .O(N__31798),
            .I(bfn_11_10_0_));
    InMux I__3491 (
            .O(N__31795),
            .I(\foc.u_Park_Transform.n783 ));
    InMux I__3490 (
            .O(N__31792),
            .I(N__31785));
    CascadeMux I__3489 (
            .O(N__31791),
            .I(N__31782));
    CascadeMux I__3488 (
            .O(N__31790),
            .I(N__31778));
    CascadeMux I__3487 (
            .O(N__31789),
            .I(N__31774));
    CascadeMux I__3486 (
            .O(N__31788),
            .I(N__31769));
    LocalMux I__3485 (
            .O(N__31785),
            .I(N__31766));
    InMux I__3484 (
            .O(N__31782),
            .I(N__31753));
    InMux I__3483 (
            .O(N__31781),
            .I(N__31753));
    InMux I__3482 (
            .O(N__31778),
            .I(N__31753));
    InMux I__3481 (
            .O(N__31777),
            .I(N__31753));
    InMux I__3480 (
            .O(N__31774),
            .I(N__31753));
    InMux I__3479 (
            .O(N__31773),
            .I(N__31753));
    InMux I__3478 (
            .O(N__31772),
            .I(N__31748));
    InMux I__3477 (
            .O(N__31769),
            .I(N__31748));
    Span4Mux_h I__3476 (
            .O(N__31766),
            .I(N__31740));
    LocalMux I__3475 (
            .O(N__31753),
            .I(N__31740));
    LocalMux I__3474 (
            .O(N__31748),
            .I(N__31740));
    InMux I__3473 (
            .O(N__31747),
            .I(N__31737));
    Span4Mux_v I__3472 (
            .O(N__31740),
            .I(N__31730));
    LocalMux I__3471 (
            .O(N__31737),
            .I(N__31727));
    CascadeMux I__3470 (
            .O(N__31736),
            .I(N__31724));
    CascadeMux I__3469 (
            .O(N__31735),
            .I(N__31720));
    CascadeMux I__3468 (
            .O(N__31734),
            .I(N__31716));
    CascadeMux I__3467 (
            .O(N__31733),
            .I(N__31711));
    Span4Mux_h I__3466 (
            .O(N__31730),
            .I(N__31706));
    Span4Mux_h I__3465 (
            .O(N__31727),
            .I(N__31706));
    InMux I__3464 (
            .O(N__31724),
            .I(N__31693));
    InMux I__3463 (
            .O(N__31723),
            .I(N__31693));
    InMux I__3462 (
            .O(N__31720),
            .I(N__31693));
    InMux I__3461 (
            .O(N__31719),
            .I(N__31693));
    InMux I__3460 (
            .O(N__31716),
            .I(N__31693));
    InMux I__3459 (
            .O(N__31715),
            .I(N__31693));
    InMux I__3458 (
            .O(N__31714),
            .I(N__31688));
    InMux I__3457 (
            .O(N__31711),
            .I(N__31688));
    Odrv4 I__3456 (
            .O(N__31706),
            .I(\foc.u_Park_Transform.n622 ));
    LocalMux I__3455 (
            .O(N__31693),
            .I(\foc.u_Park_Transform.n622 ));
    LocalMux I__3454 (
            .O(N__31688),
            .I(\foc.u_Park_Transform.n622 ));
    CascadeMux I__3453 (
            .O(N__31681),
            .I(N__31678));
    InMux I__3452 (
            .O(N__31678),
            .I(N__31675));
    LocalMux I__3451 (
            .O(N__31675),
            .I(N__31672));
    Odrv4 I__3450 (
            .O(N__31672),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552 ));
    InMux I__3449 (
            .O(N__31669),
            .I(N__31666));
    LocalMux I__3448 (
            .O(N__31666),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470 ));
    InMux I__3447 (
            .O(N__31663),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352 ));
    InMux I__3446 (
            .O(N__31660),
            .I(N__31657));
    LocalMux I__3445 (
            .O(N__31657),
            .I(N__31654));
    Odrv4 I__3444 (
            .O(N__31654),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551 ));
    CascadeMux I__3443 (
            .O(N__31651),
            .I(N__31648));
    InMux I__3442 (
            .O(N__31648),
            .I(N__31645));
    LocalMux I__3441 (
            .O(N__31645),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469 ));
    InMux I__3440 (
            .O(N__31642),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353 ));
    InMux I__3439 (
            .O(N__31639),
            .I(N__31636));
    LocalMux I__3438 (
            .O(N__31636),
            .I(N__31633));
    Odrv4 I__3437 (
            .O(N__31633),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550 ));
    InMux I__3436 (
            .O(N__31630),
            .I(N__31627));
    LocalMux I__3435 (
            .O(N__31627),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468 ));
    InMux I__3434 (
            .O(N__31624),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354 ));
    InMux I__3433 (
            .O(N__31621),
            .I(N__31618));
    LocalMux I__3432 (
            .O(N__31618),
            .I(N__31615));
    Odrv4 I__3431 (
            .O(N__31615),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549 ));
    CascadeMux I__3430 (
            .O(N__31612),
            .I(N__31609));
    InMux I__3429 (
            .O(N__31609),
            .I(N__31606));
    LocalMux I__3428 (
            .O(N__31606),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467 ));
    InMux I__3427 (
            .O(N__31603),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355 ));
    InMux I__3426 (
            .O(N__31600),
            .I(N__31597));
    LocalMux I__3425 (
            .O(N__31597),
            .I(N__31594));
    Odrv4 I__3424 (
            .O(N__31594),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548 ));
    InMux I__3423 (
            .O(N__31591),
            .I(N__31588));
    LocalMux I__3422 (
            .O(N__31588),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466 ));
    InMux I__3421 (
            .O(N__31585),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356 ));
    InMux I__3420 (
            .O(N__31582),
            .I(N__31579));
    LocalMux I__3419 (
            .O(N__31579),
            .I(N__31576));
    Odrv4 I__3418 (
            .O(N__31576),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547 ));
    CascadeMux I__3417 (
            .O(N__31573),
            .I(N__31564));
    CascadeMux I__3416 (
            .O(N__31572),
            .I(N__31558));
    CascadeMux I__3415 (
            .O(N__31571),
            .I(N__31555));
    CascadeMux I__3414 (
            .O(N__31570),
            .I(N__31551));
    CascadeMux I__3413 (
            .O(N__31569),
            .I(N__31548));
    InMux I__3412 (
            .O(N__31568),
            .I(N__31536));
    InMux I__3411 (
            .O(N__31567),
            .I(N__31536));
    InMux I__3410 (
            .O(N__31564),
            .I(N__31536));
    InMux I__3409 (
            .O(N__31563),
            .I(N__31536));
    InMux I__3408 (
            .O(N__31562),
            .I(N__31536));
    InMux I__3407 (
            .O(N__31561),
            .I(N__31529));
    InMux I__3406 (
            .O(N__31558),
            .I(N__31529));
    InMux I__3405 (
            .O(N__31555),
            .I(N__31529));
    InMux I__3404 (
            .O(N__31554),
            .I(N__31520));
    InMux I__3403 (
            .O(N__31551),
            .I(N__31520));
    InMux I__3402 (
            .O(N__31548),
            .I(N__31520));
    InMux I__3401 (
            .O(N__31547),
            .I(N__31520));
    LocalMux I__3400 (
            .O(N__31536),
            .I(N__31511));
    LocalMux I__3399 (
            .O(N__31529),
            .I(N__31511));
    LocalMux I__3398 (
            .O(N__31520),
            .I(N__31511));
    CascadeMux I__3397 (
            .O(N__31519),
            .I(N__31506));
    CascadeMux I__3396 (
            .O(N__31518),
            .I(N__31502));
    Span4Mux_v I__3395 (
            .O(N__31511),
            .I(N__31488));
    InMux I__3394 (
            .O(N__31510),
            .I(N__31473));
    InMux I__3393 (
            .O(N__31509),
            .I(N__31473));
    InMux I__3392 (
            .O(N__31506),
            .I(N__31473));
    InMux I__3391 (
            .O(N__31505),
            .I(N__31473));
    InMux I__3390 (
            .O(N__31502),
            .I(N__31473));
    InMux I__3389 (
            .O(N__31501),
            .I(N__31473));
    InMux I__3388 (
            .O(N__31500),
            .I(N__31473));
    CascadeMux I__3387 (
            .O(N__31499),
            .I(N__31469));
    CascadeMux I__3386 (
            .O(N__31498),
            .I(N__31465));
    CascadeMux I__3385 (
            .O(N__31497),
            .I(N__31461));
    CascadeMux I__3384 (
            .O(N__31496),
            .I(N__31458));
    CascadeMux I__3383 (
            .O(N__31495),
            .I(N__31454));
    CascadeMux I__3382 (
            .O(N__31494),
            .I(N__31451));
    CascadeMux I__3381 (
            .O(N__31493),
            .I(N__31448));
    CascadeMux I__3380 (
            .O(N__31492),
            .I(N__31444));
    CascadeMux I__3379 (
            .O(N__31491),
            .I(N__31441));
    Span4Mux_h I__3378 (
            .O(N__31488),
            .I(N__31434));
    LocalMux I__3377 (
            .O(N__31473),
            .I(N__31434));
    InMux I__3376 (
            .O(N__31472),
            .I(N__31419));
    InMux I__3375 (
            .O(N__31469),
            .I(N__31419));
    InMux I__3374 (
            .O(N__31468),
            .I(N__31419));
    InMux I__3373 (
            .O(N__31465),
            .I(N__31419));
    InMux I__3372 (
            .O(N__31464),
            .I(N__31419));
    InMux I__3371 (
            .O(N__31461),
            .I(N__31419));
    InMux I__3370 (
            .O(N__31458),
            .I(N__31419));
    InMux I__3369 (
            .O(N__31457),
            .I(N__31416));
    InMux I__3368 (
            .O(N__31454),
            .I(N__31413));
    InMux I__3367 (
            .O(N__31451),
            .I(N__31406));
    InMux I__3366 (
            .O(N__31448),
            .I(N__31406));
    InMux I__3365 (
            .O(N__31447),
            .I(N__31406));
    InMux I__3364 (
            .O(N__31444),
            .I(N__31397));
    InMux I__3363 (
            .O(N__31441),
            .I(N__31397));
    InMux I__3362 (
            .O(N__31440),
            .I(N__31397));
    InMux I__3361 (
            .O(N__31439),
            .I(N__31397));
    Odrv4 I__3360 (
            .O(N__31434),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    LocalMux I__3359 (
            .O(N__31419),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    LocalMux I__3358 (
            .O(N__31416),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    LocalMux I__3357 (
            .O(N__31413),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    LocalMux I__3356 (
            .O(N__31406),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    LocalMux I__3355 (
            .O(N__31397),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ));
    InMux I__3354 (
            .O(N__31384),
            .I(bfn_10_26_0_));
    InMux I__3353 (
            .O(N__31381),
            .I(N__31378));
    LocalMux I__3352 (
            .O(N__31378),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465 ));
    CascadeMux I__3351 (
            .O(N__31375),
            .I(N__31372));
    InMux I__3350 (
            .O(N__31372),
            .I(N__31369));
    LocalMux I__3349 (
            .O(N__31369),
            .I(N__31366));
    Odrv4 I__3348 (
            .O(N__31366),
            .I(\foc.u_Park_Transform.n84 ));
    CascadeMux I__3347 (
            .O(N__31363),
            .I(N__31360));
    InMux I__3346 (
            .O(N__31360),
            .I(N__31357));
    LocalMux I__3345 (
            .O(N__31357),
            .I(N__31354));
    Odrv4 I__3344 (
            .O(N__31354),
            .I(\foc.u_Park_Transform.n133_adj_2101 ));
    InMux I__3343 (
            .O(N__31351),
            .I(\foc.u_Park_Transform.n17098 ));
    InMux I__3342 (
            .O(N__31348),
            .I(N__31345));
    LocalMux I__3341 (
            .O(N__31345),
            .I(N__31342));
    Odrv12 I__3340 (
            .O(N__31342),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920 ));
    InMux I__3339 (
            .O(N__31339),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398 ));
    CascadeMux I__3338 (
            .O(N__31336),
            .I(N__31333));
    InMux I__3337 (
            .O(N__31333),
            .I(N__31330));
    LocalMux I__3336 (
            .O(N__31330),
            .I(N__31327));
    Odrv12 I__3335 (
            .O(N__31327),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020 ));
    InMux I__3334 (
            .O(N__31324),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399 ));
    CascadeMux I__3333 (
            .O(N__31321),
            .I(N__31315));
    CascadeMux I__3332 (
            .O(N__31320),
            .I(N__31311));
    CascadeMux I__3331 (
            .O(N__31319),
            .I(N__31307));
    InMux I__3330 (
            .O(N__31318),
            .I(N__31291));
    InMux I__3329 (
            .O(N__31315),
            .I(N__31291));
    InMux I__3328 (
            .O(N__31314),
            .I(N__31291));
    InMux I__3327 (
            .O(N__31311),
            .I(N__31291));
    InMux I__3326 (
            .O(N__31310),
            .I(N__31291));
    InMux I__3325 (
            .O(N__31307),
            .I(N__31291));
    InMux I__3324 (
            .O(N__31306),
            .I(N__31291));
    LocalMux I__3323 (
            .O(N__31291),
            .I(N__31288));
    Span4Mux_v I__3322 (
            .O(N__31288),
            .I(N__31284));
    InMux I__3321 (
            .O(N__31287),
            .I(N__31281));
    Odrv4 I__3320 (
            .O(N__31284),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819 ));
    LocalMux I__3319 (
            .O(N__31281),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819 ));
    InMux I__3318 (
            .O(N__31276),
            .I(N__31273));
    LocalMux I__3317 (
            .O(N__31273),
            .I(N__31270));
    Odrv12 I__3316 (
            .O(N__31270),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120 ));
    InMux I__3315 (
            .O(N__31267),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400 ));
    InMux I__3314 (
            .O(N__31264),
            .I(bfn_10_24_0_));
    InMux I__3313 (
            .O(N__31261),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228 ));
    InMux I__3312 (
            .O(N__31258),
            .I(N__31255));
    LocalMux I__3311 (
            .O(N__31255),
            .I(N__31252));
    Span4Mux_v I__3310 (
            .O(N__31252),
            .I(N__31249));
    Span4Mux_h I__3309 (
            .O(N__31249),
            .I(N__31246));
    Odrv4 I__3308 (
            .O(N__31246),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554 ));
    InMux I__3307 (
            .O(N__31243),
            .I(N__31240));
    LocalMux I__3306 (
            .O(N__31240),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472 ));
    InMux I__3305 (
            .O(N__31237),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350 ));
    CascadeMux I__3304 (
            .O(N__31234),
            .I(N__31231));
    InMux I__3303 (
            .O(N__31231),
            .I(N__31228));
    LocalMux I__3302 (
            .O(N__31228),
            .I(N__31225));
    Odrv4 I__3301 (
            .O(N__31225),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553 ));
    CascadeMux I__3300 (
            .O(N__31222),
            .I(N__31219));
    InMux I__3299 (
            .O(N__31219),
            .I(N__31216));
    LocalMux I__3298 (
            .O(N__31216),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471 ));
    InMux I__3297 (
            .O(N__31213),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351 ));
    InMux I__3296 (
            .O(N__31210),
            .I(N__31207));
    LocalMux I__3295 (
            .O(N__31207),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932 ));
    InMux I__3294 (
            .O(N__31204),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427 ));
    InMux I__3293 (
            .O(N__31201),
            .I(N__31198));
    LocalMux I__3292 (
            .O(N__31198),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032 ));
    CascadeMux I__3291 (
            .O(N__31195),
            .I(N__31188));
    CascadeMux I__3290 (
            .O(N__31194),
            .I(N__31185));
    CascadeMux I__3289 (
            .O(N__31193),
            .I(N__31182));
    CascadeMux I__3288 (
            .O(N__31192),
            .I(N__31179));
    CascadeMux I__3287 (
            .O(N__31191),
            .I(N__31175));
    InMux I__3286 (
            .O(N__31188),
            .I(N__31170));
    InMux I__3285 (
            .O(N__31185),
            .I(N__31167));
    InMux I__3284 (
            .O(N__31182),
            .I(N__31154));
    InMux I__3283 (
            .O(N__31179),
            .I(N__31154));
    InMux I__3282 (
            .O(N__31178),
            .I(N__31154));
    InMux I__3281 (
            .O(N__31175),
            .I(N__31154));
    InMux I__3280 (
            .O(N__31174),
            .I(N__31154));
    InMux I__3279 (
            .O(N__31173),
            .I(N__31154));
    LocalMux I__3278 (
            .O(N__31170),
            .I(N__31147));
    LocalMux I__3277 (
            .O(N__31167),
            .I(N__31147));
    LocalMux I__3276 (
            .O(N__31154),
            .I(N__31147));
    Odrv4 I__3275 (
            .O(N__31147),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828 ));
    InMux I__3274 (
            .O(N__31144),
            .I(bfn_10_22_0_));
    InMux I__3273 (
            .O(N__31141),
            .I(N__31138));
    LocalMux I__3272 (
            .O(N__31138),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132 ));
    InMux I__3271 (
            .O(N__31135),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429 ));
    InMux I__3270 (
            .O(N__31132),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240 ));
    CascadeMux I__3269 (
            .O(N__31129),
            .I(N__31126));
    InMux I__3268 (
            .O(N__31126),
            .I(N__31123));
    LocalMux I__3267 (
            .O(N__31123),
            .I(N__31120));
    Span12Mux_h I__3266 (
            .O(N__31120),
            .I(N__31117));
    Odrv12 I__3265 (
            .O(N__31117),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420 ));
    InMux I__3264 (
            .O(N__31114),
            .I(N__31111));
    LocalMux I__3263 (
            .O(N__31111),
            .I(N__31108));
    Span4Mux_v I__3262 (
            .O(N__31108),
            .I(N__31105));
    Odrv4 I__3261 (
            .O(N__31105),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520 ));
    InMux I__3260 (
            .O(N__31102),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394 ));
    CascadeMux I__3259 (
            .O(N__31099),
            .I(N__31096));
    InMux I__3258 (
            .O(N__31096),
            .I(N__31093));
    LocalMux I__3257 (
            .O(N__31093),
            .I(N__31090));
    Span4Mux_v I__3256 (
            .O(N__31090),
            .I(N__31087));
    Odrv4 I__3255 (
            .O(N__31087),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620 ));
    InMux I__3254 (
            .O(N__31084),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395 ));
    InMux I__3253 (
            .O(N__31081),
            .I(N__31078));
    LocalMux I__3252 (
            .O(N__31078),
            .I(N__31075));
    Odrv12 I__3251 (
            .O(N__31075),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720 ));
    InMux I__3250 (
            .O(N__31072),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396 ));
    CascadeMux I__3249 (
            .O(N__31069),
            .I(N__31066));
    InMux I__3248 (
            .O(N__31066),
            .I(N__31063));
    LocalMux I__3247 (
            .O(N__31063),
            .I(N__31060));
    Odrv12 I__3246 (
            .O(N__31060),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820 ));
    InMux I__3245 (
            .O(N__31057),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397 ));
    InMux I__3244 (
            .O(N__31054),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224 ));
    InMux I__3243 (
            .O(N__31051),
            .I(N__31048));
    LocalMux I__3242 (
            .O(N__31048),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332 ));
    InMux I__3241 (
            .O(N__31045),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421 ));
    CascadeMux I__3240 (
            .O(N__31042),
            .I(N__31039));
    InMux I__3239 (
            .O(N__31039),
            .I(N__31036));
    LocalMux I__3238 (
            .O(N__31036),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432 ));
    InMux I__3237 (
            .O(N__31033),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422 ));
    InMux I__3236 (
            .O(N__31030),
            .I(N__31027));
    LocalMux I__3235 (
            .O(N__31027),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532 ));
    InMux I__3234 (
            .O(N__31024),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423 ));
    CascadeMux I__3233 (
            .O(N__31021),
            .I(N__31018));
    InMux I__3232 (
            .O(N__31018),
            .I(N__31015));
    LocalMux I__3231 (
            .O(N__31015),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632 ));
    InMux I__3230 (
            .O(N__31012),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424 ));
    InMux I__3229 (
            .O(N__31009),
            .I(N__31006));
    LocalMux I__3228 (
            .O(N__31006),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732 ));
    InMux I__3227 (
            .O(N__31003),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425 ));
    InMux I__3226 (
            .O(N__31000),
            .I(N__30997));
    LocalMux I__3225 (
            .O(N__30997),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832 ));
    InMux I__3224 (
            .O(N__30994),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426 ));
    InMux I__3223 (
            .O(N__30991),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385 ));
    InMux I__3222 (
            .O(N__30988),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386 ));
    InMux I__3221 (
            .O(N__30985),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387 ));
    InMux I__3220 (
            .O(N__30982),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388 ));
    InMux I__3219 (
            .O(N__30979),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389 ));
    InMux I__3218 (
            .O(N__30976),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390 ));
    InMux I__3217 (
            .O(N__30973),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391 ));
    InMux I__3216 (
            .O(N__30970),
            .I(bfn_10_20_0_));
    CascadeMux I__3215 (
            .O(N__30967),
            .I(N__30964));
    InMux I__3214 (
            .O(N__30964),
            .I(N__30961));
    LocalMux I__3213 (
            .O(N__30961),
            .I(N__30958));
    Odrv12 I__3212 (
            .O(N__30958),
            .I(\foc.u_Park_Transform.n231 ));
    CascadeMux I__3211 (
            .O(N__30955),
            .I(N__30952));
    InMux I__3210 (
            .O(N__30952),
            .I(N__30949));
    LocalMux I__3209 (
            .O(N__30949),
            .I(N__30946));
    Span4Mux_v I__3208 (
            .O(N__30946),
            .I(N__30943));
    Odrv4 I__3207 (
            .O(N__30943),
            .I(\foc.u_Park_Transform.n277 ));
    InMux I__3206 (
            .O(N__30940),
            .I(\foc.u_Park_Transform.n16927 ));
    InMux I__3205 (
            .O(N__30937),
            .I(N__30934));
    LocalMux I__3204 (
            .O(N__30934),
            .I(N__30931));
    Odrv4 I__3203 (
            .O(N__30931),
            .I(\foc.u_Park_Transform.n280 ));
    CascadeMux I__3202 (
            .O(N__30928),
            .I(N__30925));
    InMux I__3201 (
            .O(N__30925),
            .I(N__30922));
    LocalMux I__3200 (
            .O(N__30922),
            .I(N__30919));
    Odrv4 I__3199 (
            .O(N__30919),
            .I(\foc.u_Park_Transform.n326 ));
    InMux I__3198 (
            .O(N__30916),
            .I(\foc.u_Park_Transform.n16928 ));
    CascadeMux I__3197 (
            .O(N__30913),
            .I(N__30910));
    InMux I__3196 (
            .O(N__30910),
            .I(N__30907));
    LocalMux I__3195 (
            .O(N__30907),
            .I(N__30904));
    Odrv4 I__3194 (
            .O(N__30904),
            .I(\foc.u_Park_Transform.n329 ));
    CascadeMux I__3193 (
            .O(N__30901),
            .I(N__30898));
    InMux I__3192 (
            .O(N__30898),
            .I(N__30895));
    LocalMux I__3191 (
            .O(N__30895),
            .I(N__30892));
    Span4Mux_v I__3190 (
            .O(N__30892),
            .I(N__30889));
    Odrv4 I__3189 (
            .O(N__30889),
            .I(\foc.u_Park_Transform.n375 ));
    InMux I__3188 (
            .O(N__30886),
            .I(\foc.u_Park_Transform.n16929 ));
    InMux I__3187 (
            .O(N__30883),
            .I(N__30880));
    LocalMux I__3186 (
            .O(N__30880),
            .I(N__30877));
    Odrv4 I__3185 (
            .O(N__30877),
            .I(\foc.u_Park_Transform.n378 ));
    InMux I__3184 (
            .O(N__30874),
            .I(N__30871));
    LocalMux I__3183 (
            .O(N__30871),
            .I(\foc.u_Park_Transform.n424 ));
    InMux I__3182 (
            .O(N__30868),
            .I(\foc.u_Park_Transform.n16930 ));
    CascadeMux I__3181 (
            .O(N__30865),
            .I(N__30862));
    InMux I__3180 (
            .O(N__30862),
            .I(N__30859));
    LocalMux I__3179 (
            .O(N__30859),
            .I(N__30856));
    Odrv4 I__3178 (
            .O(N__30856),
            .I(\foc.u_Park_Transform.n473 ));
    InMux I__3177 (
            .O(N__30853),
            .I(bfn_10_18_0_));
    CascadeMux I__3176 (
            .O(N__30850),
            .I(N__30841));
    CascadeMux I__3175 (
            .O(N__30849),
            .I(N__30834));
    CascadeMux I__3174 (
            .O(N__30848),
            .I(N__30830));
    CascadeMux I__3173 (
            .O(N__30847),
            .I(N__30826));
    CascadeMux I__3172 (
            .O(N__30846),
            .I(N__30822));
    CascadeMux I__3171 (
            .O(N__30845),
            .I(N__30817));
    InMux I__3170 (
            .O(N__30844),
            .I(N__30812));
    InMux I__3169 (
            .O(N__30841),
            .I(N__30812));
    CascadeMux I__3168 (
            .O(N__30840),
            .I(N__30809));
    CascadeMux I__3167 (
            .O(N__30839),
            .I(N__30805));
    CascadeMux I__3166 (
            .O(N__30838),
            .I(N__30801));
    CascadeMux I__3165 (
            .O(N__30837),
            .I(N__30797));
    InMux I__3164 (
            .O(N__30834),
            .I(N__30791));
    InMux I__3163 (
            .O(N__30833),
            .I(N__30791));
    InMux I__3162 (
            .O(N__30830),
            .I(N__30778));
    InMux I__3161 (
            .O(N__30829),
            .I(N__30778));
    InMux I__3160 (
            .O(N__30826),
            .I(N__30778));
    InMux I__3159 (
            .O(N__30825),
            .I(N__30778));
    InMux I__3158 (
            .O(N__30822),
            .I(N__30778));
    InMux I__3157 (
            .O(N__30821),
            .I(N__30778));
    InMux I__3156 (
            .O(N__30820),
            .I(N__30773));
    InMux I__3155 (
            .O(N__30817),
            .I(N__30773));
    LocalMux I__3154 (
            .O(N__30812),
            .I(N__30770));
    InMux I__3153 (
            .O(N__30809),
            .I(N__30765));
    InMux I__3152 (
            .O(N__30808),
            .I(N__30765));
    InMux I__3151 (
            .O(N__30805),
            .I(N__30751));
    InMux I__3150 (
            .O(N__30804),
            .I(N__30751));
    InMux I__3149 (
            .O(N__30801),
            .I(N__30751));
    InMux I__3148 (
            .O(N__30800),
            .I(N__30751));
    InMux I__3147 (
            .O(N__30797),
            .I(N__30751));
    InMux I__3146 (
            .O(N__30796),
            .I(N__30751));
    LocalMux I__3145 (
            .O(N__30791),
            .I(N__30748));
    LocalMux I__3144 (
            .O(N__30778),
            .I(N__30743));
    LocalMux I__3143 (
            .O(N__30773),
            .I(N__30743));
    Span4Mux_v I__3142 (
            .O(N__30770),
            .I(N__30738));
    LocalMux I__3141 (
            .O(N__30765),
            .I(N__30738));
    InMux I__3140 (
            .O(N__30764),
            .I(N__30735));
    LocalMux I__3139 (
            .O(N__30751),
            .I(N__30731));
    Span4Mux_v I__3138 (
            .O(N__30748),
            .I(N__30722));
    Span4Mux_v I__3137 (
            .O(N__30743),
            .I(N__30722));
    Span4Mux_h I__3136 (
            .O(N__30738),
            .I(N__30722));
    LocalMux I__3135 (
            .O(N__30735),
            .I(N__30722));
    InMux I__3134 (
            .O(N__30734),
            .I(N__30719));
    Odrv12 I__3133 (
            .O(N__30731),
            .I(\foc.u_Park_Transform.n619 ));
    Odrv4 I__3132 (
            .O(N__30722),
            .I(\foc.u_Park_Transform.n619 ));
    LocalMux I__3131 (
            .O(N__30719),
            .I(\foc.u_Park_Transform.n619 ));
    CascadeMux I__3130 (
            .O(N__30712),
            .I(N__30708));
    InMux I__3129 (
            .O(N__30711),
            .I(N__30700));
    InMux I__3128 (
            .O(N__30708),
            .I(N__30700));
    InMux I__3127 (
            .O(N__30707),
            .I(N__30700));
    LocalMux I__3126 (
            .O(N__30700),
            .I(N__30697));
    Odrv4 I__3125 (
            .O(N__30697),
            .I(\foc.u_Park_Transform.n522 ));
    InMux I__3124 (
            .O(N__30694),
            .I(\foc.u_Park_Transform.n16932 ));
    InMux I__3123 (
            .O(N__30691),
            .I(N__30688));
    LocalMux I__3122 (
            .O(N__30688),
            .I(N__30684));
    InMux I__3121 (
            .O(N__30687),
            .I(N__30681));
    Span12Mux_h I__3120 (
            .O(N__30684),
            .I(N__30676));
    LocalMux I__3119 (
            .O(N__30681),
            .I(N__30676));
    Odrv12 I__3118 (
            .O(N__30676),
            .I(\foc.u_Park_Transform.n777 ));
    CascadeMux I__3117 (
            .O(N__30673),
            .I(N__30669));
    CascadeMux I__3116 (
            .O(N__30672),
            .I(N__30665));
    InMux I__3115 (
            .O(N__30669),
            .I(N__30658));
    InMux I__3114 (
            .O(N__30668),
            .I(N__30658));
    InMux I__3113 (
            .O(N__30665),
            .I(N__30658));
    LocalMux I__3112 (
            .O(N__30658),
            .I(N__30655));
    Odrv12 I__3111 (
            .O(N__30655),
            .I(\foc.u_Park_Transform.n427 ));
    InMux I__3110 (
            .O(N__30652),
            .I(\foc.u_Park_Transform.n16933 ));
    InMux I__3109 (
            .O(N__30649),
            .I(\foc.u_Park_Transform.n779 ));
    InMux I__3108 (
            .O(N__30646),
            .I(N__30643));
    LocalMux I__3107 (
            .O(N__30643),
            .I(\foc.u_Park_Transform.n283 ));
    InMux I__3106 (
            .O(N__30640),
            .I(\foc.u_Park_Transform.n16919 ));
    InMux I__3105 (
            .O(N__30637),
            .I(\foc.u_Park_Transform.n16920 ));
    InMux I__3104 (
            .O(N__30634),
            .I(\foc.u_Park_Transform.n16921 ));
    CascadeMux I__3103 (
            .O(N__30631),
            .I(N__30628));
    InMux I__3102 (
            .O(N__30628),
            .I(N__30624));
    CascadeMux I__3101 (
            .O(N__30627),
            .I(N__30620));
    LocalMux I__3100 (
            .O(N__30624),
            .I(N__30617));
    InMux I__3099 (
            .O(N__30623),
            .I(N__30612));
    InMux I__3098 (
            .O(N__30620),
            .I(N__30612));
    Odrv4 I__3097 (
            .O(N__30617),
            .I(\foc.u_Park_Transform.n332 ));
    LocalMux I__3096 (
            .O(N__30612),
            .I(\foc.u_Park_Transform.n332 ));
    InMux I__3095 (
            .O(N__30607),
            .I(bfn_10_16_0_));
    InMux I__3094 (
            .O(N__30604),
            .I(\foc.u_Park_Transform.n783_adj_2167 ));
    CascadeMux I__3093 (
            .O(N__30601),
            .I(N__30598));
    InMux I__3092 (
            .O(N__30598),
            .I(N__30595));
    LocalMux I__3091 (
            .O(N__30595),
            .I(N__30592));
    Odrv4 I__3090 (
            .O(N__30592),
            .I(\foc.u_Park_Transform.n81_adj_2120 ));
    CascadeMux I__3089 (
            .O(N__30589),
            .I(N__30586));
    InMux I__3088 (
            .O(N__30586),
            .I(N__30583));
    LocalMux I__3087 (
            .O(N__30583),
            .I(N__30580));
    Odrv4 I__3086 (
            .O(N__30580),
            .I(\foc.u_Park_Transform.n84_adj_2118 ));
    CascadeMux I__3085 (
            .O(N__30577),
            .I(N__30574));
    InMux I__3084 (
            .O(N__30574),
            .I(N__30571));
    LocalMux I__3083 (
            .O(N__30571),
            .I(N__30568));
    Span4Mux_h I__3082 (
            .O(N__30568),
            .I(N__30565));
    Odrv4 I__3081 (
            .O(N__30565),
            .I(\foc.u_Park_Transform.n130_adj_2105 ));
    InMux I__3080 (
            .O(N__30562),
            .I(\foc.u_Park_Transform.n16924 ));
    CascadeMux I__3079 (
            .O(N__30559),
            .I(N__30556));
    InMux I__3078 (
            .O(N__30556),
            .I(N__30553));
    LocalMux I__3077 (
            .O(N__30553),
            .I(N__30550));
    Odrv12 I__3076 (
            .O(N__30550),
            .I(\foc.u_Park_Transform.n133 ));
    CascadeMux I__3075 (
            .O(N__30547),
            .I(N__30544));
    InMux I__3074 (
            .O(N__30544),
            .I(N__30541));
    LocalMux I__3073 (
            .O(N__30541),
            .I(N__30538));
    Odrv4 I__3072 (
            .O(N__30538),
            .I(\foc.u_Park_Transform.n179_adj_2076 ));
    InMux I__3071 (
            .O(N__30535),
            .I(\foc.u_Park_Transform.n16925 ));
    InMux I__3070 (
            .O(N__30532),
            .I(N__30529));
    LocalMux I__3069 (
            .O(N__30529),
            .I(N__30526));
    Odrv4 I__3068 (
            .O(N__30526),
            .I(\foc.u_Park_Transform.n182 ));
    CascadeMux I__3067 (
            .O(N__30523),
            .I(N__30520));
    InMux I__3066 (
            .O(N__30520),
            .I(N__30517));
    LocalMux I__3065 (
            .O(N__30517),
            .I(N__30514));
    Odrv4 I__3064 (
            .O(N__30514),
            .I(\foc.u_Park_Transform.n228 ));
    InMux I__3063 (
            .O(N__30511),
            .I(\foc.u_Park_Transform.n16926 ));
    InMux I__3062 (
            .O(N__30508),
            .I(\foc.u_Park_Transform.n18164 ));
    InMux I__3061 (
            .O(N__30505),
            .I(\foc.u_Park_Transform.n18165 ));
    InMux I__3060 (
            .O(N__30502),
            .I(\foc.u_Park_Transform.n787 ));
    CascadeMux I__3059 (
            .O(N__30499),
            .I(N__30496));
    InMux I__3058 (
            .O(N__30496),
            .I(N__30493));
    LocalMux I__3057 (
            .O(N__30493),
            .I(\foc.u_Park_Transform.n87 ));
    InMux I__3056 (
            .O(N__30490),
            .I(\foc.u_Park_Transform.n16915 ));
    CascadeMux I__3055 (
            .O(N__30487),
            .I(N__30484));
    InMux I__3054 (
            .O(N__30484),
            .I(N__30481));
    LocalMux I__3053 (
            .O(N__30481),
            .I(\foc.u_Park_Transform.n136 ));
    InMux I__3052 (
            .O(N__30478),
            .I(\foc.u_Park_Transform.n16916 ));
    InMux I__3051 (
            .O(N__30475),
            .I(N__30472));
    LocalMux I__3050 (
            .O(N__30472),
            .I(\foc.u_Park_Transform.n185 ));
    InMux I__3049 (
            .O(N__30469),
            .I(\foc.u_Park_Transform.n16917 ));
    CascadeMux I__3048 (
            .O(N__30466),
            .I(N__30463));
    InMux I__3047 (
            .O(N__30463),
            .I(N__30460));
    LocalMux I__3046 (
            .O(N__30460),
            .I(\foc.u_Park_Transform.n234 ));
    InMux I__3045 (
            .O(N__30457),
            .I(\foc.u_Park_Transform.n16918 ));
    InMux I__3044 (
            .O(N__30454),
            .I(\foc.u_Park_Transform.n771_adj_2032 ));
    CascadeMux I__3043 (
            .O(N__30451),
            .I(N__30448));
    InMux I__3042 (
            .O(N__30448),
            .I(N__30444));
    CascadeMux I__3041 (
            .O(N__30447),
            .I(N__30441));
    LocalMux I__3040 (
            .O(N__30444),
            .I(N__30438));
    InMux I__3039 (
            .O(N__30441),
            .I(N__30435));
    Odrv4 I__3038 (
            .O(N__30438),
            .I(\foc.u_Park_Transform.n773 ));
    LocalMux I__3037 (
            .O(N__30435),
            .I(\foc.u_Park_Transform.n773 ));
    InMux I__3036 (
            .O(N__30430),
            .I(\foc.u_Park_Transform.n18160 ));
    InMux I__3035 (
            .O(N__30427),
            .I(\foc.u_Park_Transform.n18161 ));
    InMux I__3034 (
            .O(N__30424),
            .I(\foc.u_Park_Transform.n18162 ));
    InMux I__3033 (
            .O(N__30421),
            .I(\foc.u_Park_Transform.n18163 ));
    InMux I__3032 (
            .O(N__30418),
            .I(N__30415));
    LocalMux I__3031 (
            .O(N__30415),
            .I(\foc.u_Park_Transform.n372 ));
    InMux I__3030 (
            .O(N__30412),
            .I(N__30409));
    LocalMux I__3029 (
            .O(N__30409),
            .I(\foc.u_Park_Transform.n418_adj_2024 ));
    InMux I__3028 (
            .O(N__30406),
            .I(\foc.u_Park_Transform.n17137 ));
    InMux I__3027 (
            .O(N__30403),
            .I(N__30400));
    LocalMux I__3026 (
            .O(N__30400),
            .I(\foc.u_Park_Transform.n421_adj_2039 ));
    CascadeMux I__3025 (
            .O(N__30397),
            .I(N__30394));
    InMux I__3024 (
            .O(N__30394),
            .I(N__30391));
    LocalMux I__3023 (
            .O(N__30391),
            .I(N__30388));
    Odrv4 I__3022 (
            .O(N__30388),
            .I(\foc.u_Park_Transform.n467_adj_2019 ));
    InMux I__3021 (
            .O(N__30385),
            .I(bfn_10_12_0_));
    CascadeMux I__3020 (
            .O(N__30382),
            .I(N__30379));
    InMux I__3019 (
            .O(N__30379),
            .I(N__30376));
    LocalMux I__3018 (
            .O(N__30376),
            .I(\foc.u_Park_Transform.n470_adj_2038 ));
    InMux I__3017 (
            .O(N__30373),
            .I(N__30370));
    LocalMux I__3016 (
            .O(N__30370),
            .I(N__30367));
    Odrv4 I__3015 (
            .O(N__30367),
            .I(\foc.u_Park_Transform.n516_adj_2018 ));
    InMux I__3014 (
            .O(N__30364),
            .I(\foc.u_Park_Transform.n17139 ));
    InMux I__3013 (
            .O(N__30361),
            .I(N__30358));
    LocalMux I__3012 (
            .O(N__30358),
            .I(\foc.u_Park_Transform.n519_adj_2035 ));
    CascadeMux I__3011 (
            .O(N__30355),
            .I(N__30352));
    InMux I__3010 (
            .O(N__30352),
            .I(N__30349));
    LocalMux I__3009 (
            .O(N__30349),
            .I(N__30346));
    Odrv4 I__3008 (
            .O(N__30346),
            .I(\foc.u_Park_Transform.n565 ));
    InMux I__3007 (
            .O(N__30343),
            .I(\foc.u_Park_Transform.n17140 ));
    CascadeMux I__3006 (
            .O(N__30340),
            .I(N__30337));
    InMux I__3005 (
            .O(N__30337),
            .I(N__30334));
    LocalMux I__3004 (
            .O(N__30334),
            .I(\foc.u_Park_Transform.n568_adj_2034 ));
    InMux I__3003 (
            .O(N__30331),
            .I(N__30328));
    LocalMux I__3002 (
            .O(N__30328),
            .I(N__30325));
    Odrv4 I__3001 (
            .O(N__30325),
            .I(\foc.u_Park_Transform.n614_adj_2017 ));
    InMux I__3000 (
            .O(N__30322),
            .I(\foc.u_Park_Transform.n17141 ));
    CascadeMux I__2999 (
            .O(N__30319),
            .I(N__30316));
    InMux I__2998 (
            .O(N__30316),
            .I(N__30313));
    LocalMux I__2997 (
            .O(N__30313),
            .I(N__30310));
    Odrv4 I__2996 (
            .O(N__30310),
            .I(\foc.u_Park_Transform.n663_adj_2016 ));
    InMux I__2995 (
            .O(N__30307),
            .I(\foc.u_Park_Transform.n17142 ));
    CascadeMux I__2994 (
            .O(N__30304),
            .I(N__30301));
    InMux I__2993 (
            .O(N__30301),
            .I(N__30298));
    LocalMux I__2992 (
            .O(N__30298),
            .I(N__30295));
    Odrv4 I__2991 (
            .O(N__30295),
            .I(\foc.u_Park_Transform.n712_adj_2015 ));
    InMux I__2990 (
            .O(N__30292),
            .I(\foc.u_Park_Transform.n17143 ));
    CascadeMux I__2989 (
            .O(N__30289),
            .I(N__30285));
    CascadeMux I__2988 (
            .O(N__30288),
            .I(N__30282));
    InMux I__2987 (
            .O(N__30285),
            .I(N__30278));
    InMux I__2986 (
            .O(N__30282),
            .I(N__30273));
    InMux I__2985 (
            .O(N__30281),
            .I(N__30273));
    LocalMux I__2984 (
            .O(N__30278),
            .I(\foc.u_Park_Transform.n617_adj_2031 ));
    LocalMux I__2983 (
            .O(N__30273),
            .I(\foc.u_Park_Transform.n617_adj_2031 ));
    InMux I__2982 (
            .O(N__30268),
            .I(\foc.u_Park_Transform.n17144 ));
    InMux I__2981 (
            .O(N__30265),
            .I(\foc.u_Park_Transform.n767 ));
    CascadeMux I__2980 (
            .O(N__30262),
            .I(N__30259));
    InMux I__2979 (
            .O(N__30259),
            .I(N__30256));
    LocalMux I__2978 (
            .O(N__30256),
            .I(N__30253));
    Odrv4 I__2977 (
            .O(N__30253),
            .I(\foc.u_Park_Transform.n75 ));
    CascadeMux I__2976 (
            .O(N__30250),
            .I(N__30247));
    InMux I__2975 (
            .O(N__30247),
            .I(N__30244));
    LocalMux I__2974 (
            .O(N__30244),
            .I(\foc.u_Park_Transform.n78 ));
    CascadeMux I__2973 (
            .O(N__30241),
            .I(N__30238));
    InMux I__2972 (
            .O(N__30238),
            .I(N__30235));
    LocalMux I__2971 (
            .O(N__30235),
            .I(N__30232));
    Odrv4 I__2970 (
            .O(N__30232),
            .I(\foc.u_Park_Transform.n124 ));
    InMux I__2969 (
            .O(N__30229),
            .I(\foc.u_Park_Transform.n17131 ));
    CascadeMux I__2968 (
            .O(N__30226),
            .I(N__30223));
    InMux I__2967 (
            .O(N__30223),
            .I(N__30220));
    LocalMux I__2966 (
            .O(N__30220),
            .I(\foc.u_Park_Transform.n127 ));
    InMux I__2965 (
            .O(N__30217),
            .I(N__30214));
    LocalMux I__2964 (
            .O(N__30214),
            .I(N__30211));
    Odrv4 I__2963 (
            .O(N__30211),
            .I(\foc.u_Park_Transform.n173 ));
    InMux I__2962 (
            .O(N__30208),
            .I(\foc.u_Park_Transform.n17132 ));
    InMux I__2961 (
            .O(N__30205),
            .I(N__30202));
    LocalMux I__2960 (
            .O(N__30202),
            .I(\foc.u_Park_Transform.n176 ));
    CascadeMux I__2959 (
            .O(N__30199),
            .I(N__30196));
    InMux I__2958 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__2957 (
            .O(N__30193),
            .I(N__30190));
    Odrv4 I__2956 (
            .O(N__30190),
            .I(\foc.u_Park_Transform.n222 ));
    InMux I__2955 (
            .O(N__30187),
            .I(\foc.u_Park_Transform.n17133 ));
    CascadeMux I__2954 (
            .O(N__30184),
            .I(N__30181));
    InMux I__2953 (
            .O(N__30181),
            .I(N__30178));
    LocalMux I__2952 (
            .O(N__30178),
            .I(\foc.u_Park_Transform.n225 ));
    InMux I__2951 (
            .O(N__30175),
            .I(N__30172));
    LocalMux I__2950 (
            .O(N__30172),
            .I(N__30169));
    Odrv4 I__2949 (
            .O(N__30169),
            .I(\foc.u_Park_Transform.n271 ));
    InMux I__2948 (
            .O(N__30166),
            .I(\foc.u_Park_Transform.n17134 ));
    InMux I__2947 (
            .O(N__30163),
            .I(N__30160));
    LocalMux I__2946 (
            .O(N__30160),
            .I(\foc.u_Park_Transform.n274 ));
    CascadeMux I__2945 (
            .O(N__30157),
            .I(N__30154));
    InMux I__2944 (
            .O(N__30154),
            .I(N__30151));
    LocalMux I__2943 (
            .O(N__30151),
            .I(N__30148));
    Odrv4 I__2942 (
            .O(N__30148),
            .I(\foc.u_Park_Transform.n320 ));
    InMux I__2941 (
            .O(N__30145),
            .I(\foc.u_Park_Transform.n17135 ));
    CascadeMux I__2940 (
            .O(N__30142),
            .I(N__30139));
    InMux I__2939 (
            .O(N__30139),
            .I(N__30136));
    LocalMux I__2938 (
            .O(N__30136),
            .I(\foc.u_Park_Transform.n323 ));
    InMux I__2937 (
            .O(N__30133),
            .I(N__30130));
    LocalMux I__2936 (
            .O(N__30130),
            .I(N__30127));
    Odrv12 I__2935 (
            .O(N__30127),
            .I(\foc.u_Park_Transform.n369 ));
    InMux I__2934 (
            .O(N__30124),
            .I(\foc.u_Park_Transform.n17136 ));
    InMux I__2933 (
            .O(N__30121),
            .I(\foc.u_Park_Transform.n17151 ));
    InMux I__2932 (
            .O(N__30118),
            .I(\foc.u_Park_Transform.n17152 ));
    InMux I__2931 (
            .O(N__30115),
            .I(bfn_10_10_0_));
    InMux I__2930 (
            .O(N__30112),
            .I(\foc.u_Park_Transform.n17154 ));
    InMux I__2929 (
            .O(N__30109),
            .I(\foc.u_Park_Transform.n17155 ));
    InMux I__2928 (
            .O(N__30106),
            .I(\foc.u_Park_Transform.n17156 ));
    InMux I__2927 (
            .O(N__30103),
            .I(\foc.u_Park_Transform.n17157 ));
    InMux I__2926 (
            .O(N__30100),
            .I(\foc.u_Park_Transform.n17158 ));
    InMux I__2925 (
            .O(N__30097),
            .I(\foc.u_Park_Transform.n17159 ));
    InMux I__2924 (
            .O(N__30094),
            .I(N__30091));
    LocalMux I__2923 (
            .O(N__30091),
            .I(N__30088));
    Odrv4 I__2922 (
            .O(N__30088),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047 ));
    InMux I__2921 (
            .O(N__30085),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487 ));
    InMux I__2920 (
            .O(N__30082),
            .I(N__30079));
    LocalMux I__2919 (
            .O(N__30079),
            .I(N__30076));
    Span4Mux_v I__2918 (
            .O(N__30076),
            .I(N__30073));
    Odrv4 I__2917 (
            .O(N__30073),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147 ));
    InMux I__2916 (
            .O(N__30070),
            .I(bfn_9_25_0_));
    InMux I__2915 (
            .O(N__30067),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489 ));
    InMux I__2914 (
            .O(N__30064),
            .I(\foc.u_Park_Transform.n17146 ));
    InMux I__2913 (
            .O(N__30061),
            .I(\foc.u_Park_Transform.n17147 ));
    InMux I__2912 (
            .O(N__30058),
            .I(\foc.u_Park_Transform.n17148 ));
    InMux I__2911 (
            .O(N__30055),
            .I(\foc.u_Park_Transform.n17149 ));
    InMux I__2910 (
            .O(N__30052),
            .I(\foc.u_Park_Transform.n17150 ));
    InMux I__2909 (
            .O(N__30049),
            .I(N__30046));
    LocalMux I__2908 (
            .O(N__30046),
            .I(N__30043));
    Span4Mux_h I__2907 (
            .O(N__30043),
            .I(N__30040));
    Odrv4 I__2906 (
            .O(N__30040),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891 ));
    InMux I__2905 (
            .O(N__30037),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343 ));
    InMux I__2904 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__2903 (
            .O(N__30031),
            .I(N__30028));
    Span4Mux_v I__2902 (
            .O(N__30028),
            .I(N__30025));
    Odrv4 I__2901 (
            .O(N__30025),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347 ));
    InMux I__2900 (
            .O(N__30022),
            .I(N__30019));
    LocalMux I__2899 (
            .O(N__30019),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473 ));
    CascadeMux I__2898 (
            .O(N__30016),
            .I(N__30013));
    InMux I__2897 (
            .O(N__30013),
            .I(N__30010));
    LocalMux I__2896 (
            .O(N__30010),
            .I(N__30007));
    Span4Mux_v I__2895 (
            .O(N__30007),
            .I(N__30004));
    Odrv4 I__2894 (
            .O(N__30004),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447 ));
    InMux I__2893 (
            .O(N__30001),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481 ));
    InMux I__2892 (
            .O(N__29998),
            .I(N__29995));
    LocalMux I__2891 (
            .O(N__29995),
            .I(N__29992));
    Span4Mux_h I__2890 (
            .O(N__29992),
            .I(N__29989));
    Odrv4 I__2889 (
            .O(N__29989),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547 ));
    InMux I__2888 (
            .O(N__29986),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482 ));
    CascadeMux I__2887 (
            .O(N__29983),
            .I(N__29980));
    InMux I__2886 (
            .O(N__29980),
            .I(N__29977));
    LocalMux I__2885 (
            .O(N__29977),
            .I(N__29974));
    Span4Mux_v I__2884 (
            .O(N__29974),
            .I(N__29971));
    Odrv4 I__2883 (
            .O(N__29971),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647 ));
    InMux I__2882 (
            .O(N__29968),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483 ));
    InMux I__2881 (
            .O(N__29965),
            .I(N__29962));
    LocalMux I__2880 (
            .O(N__29962),
            .I(N__29959));
    Span4Mux_h I__2879 (
            .O(N__29959),
            .I(N__29956));
    Odrv4 I__2878 (
            .O(N__29956),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747 ));
    InMux I__2877 (
            .O(N__29953),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484 ));
    InMux I__2876 (
            .O(N__29950),
            .I(N__29947));
    LocalMux I__2875 (
            .O(N__29947),
            .I(N__29944));
    Span4Mux_h I__2874 (
            .O(N__29944),
            .I(N__29941));
    Odrv4 I__2873 (
            .O(N__29941),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847 ));
    InMux I__2872 (
            .O(N__29938),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485 ));
    InMux I__2871 (
            .O(N__29935),
            .I(N__29932));
    LocalMux I__2870 (
            .O(N__29932),
            .I(N__29929));
    Span4Mux_v I__2869 (
            .O(N__29929),
            .I(N__29926));
    Odrv4 I__2868 (
            .O(N__29926),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947 ));
    InMux I__2867 (
            .O(N__29923),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486 ));
    InMux I__2866 (
            .O(N__29920),
            .I(N__29917));
    LocalMux I__2865 (
            .O(N__29917),
            .I(N__29914));
    Span4Mux_v I__2864 (
            .O(N__29914),
            .I(N__29911));
    Odrv4 I__2863 (
            .O(N__29911),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135 ));
    InMux I__2862 (
            .O(N__29908),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439 ));
    InMux I__2861 (
            .O(N__29905),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244 ));
    InMux I__2860 (
            .O(N__29902),
            .I(N__29899));
    LocalMux I__2859 (
            .O(N__29899),
            .I(N__29896));
    Span4Mux_v I__2858 (
            .O(N__29896),
            .I(N__29893));
    Odrv4 I__2857 (
            .O(N__29893),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897 ));
    InMux I__2856 (
            .O(N__29890),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337 ));
    CascadeMux I__2855 (
            .O(N__29887),
            .I(N__29884));
    InMux I__2854 (
            .O(N__29884),
            .I(N__29881));
    LocalMux I__2853 (
            .O(N__29881),
            .I(N__29878));
    Span4Mux_h I__2852 (
            .O(N__29878),
            .I(N__29875));
    Odrv4 I__2851 (
            .O(N__29875),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896 ));
    InMux I__2850 (
            .O(N__29872),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338 ));
    InMux I__2849 (
            .O(N__29869),
            .I(N__29866));
    LocalMux I__2848 (
            .O(N__29866),
            .I(N__29863));
    Span4Mux_v I__2847 (
            .O(N__29863),
            .I(N__29860));
    Odrv4 I__2846 (
            .O(N__29860),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895 ));
    InMux I__2845 (
            .O(N__29857),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339 ));
    CascadeMux I__2844 (
            .O(N__29854),
            .I(N__29851));
    InMux I__2843 (
            .O(N__29851),
            .I(N__29848));
    LocalMux I__2842 (
            .O(N__29848),
            .I(N__29845));
    Span4Mux_v I__2841 (
            .O(N__29845),
            .I(N__29842));
    Odrv4 I__2840 (
            .O(N__29842),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894 ));
    InMux I__2839 (
            .O(N__29839),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340 ));
    InMux I__2838 (
            .O(N__29836),
            .I(N__29833));
    LocalMux I__2837 (
            .O(N__29833),
            .I(N__29830));
    Span4Mux_h I__2836 (
            .O(N__29830),
            .I(N__29827));
    Odrv4 I__2835 (
            .O(N__29827),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893 ));
    InMux I__2834 (
            .O(N__29824),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341 ));
    CascadeMux I__2833 (
            .O(N__29821),
            .I(N__29818));
    InMux I__2832 (
            .O(N__29818),
            .I(N__29815));
    LocalMux I__2831 (
            .O(N__29815),
            .I(N__29812));
    Span12Mux_s11_v I__2830 (
            .O(N__29812),
            .I(N__29809));
    Odrv12 I__2829 (
            .O(N__29809),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892 ));
    InMux I__2828 (
            .O(N__29806),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342 ));
    InMux I__2827 (
            .O(N__29803),
            .I(N__29800));
    LocalMux I__2826 (
            .O(N__29800),
            .I(N__29797));
    Span4Mux_h I__2825 (
            .O(N__29797),
            .I(N__29794));
    Odrv4 I__2824 (
            .O(N__29794),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335 ));
    InMux I__2823 (
            .O(N__29791),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431 ));
    InMux I__2822 (
            .O(N__29788),
            .I(N__29785));
    LocalMux I__2821 (
            .O(N__29785),
            .I(N__29782));
    Span4Mux_v I__2820 (
            .O(N__29782),
            .I(N__29779));
    Odrv4 I__2819 (
            .O(N__29779),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435 ));
    InMux I__2818 (
            .O(N__29776),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432 ));
    CascadeMux I__2817 (
            .O(N__29773),
            .I(N__29770));
    InMux I__2816 (
            .O(N__29770),
            .I(N__29767));
    LocalMux I__2815 (
            .O(N__29767),
            .I(N__29764));
    Span4Mux_v I__2814 (
            .O(N__29764),
            .I(N__29761));
    Odrv4 I__2813 (
            .O(N__29761),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535 ));
    InMux I__2812 (
            .O(N__29758),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433 ));
    InMux I__2811 (
            .O(N__29755),
            .I(N__29752));
    LocalMux I__2810 (
            .O(N__29752),
            .I(N__29749));
    Span4Mux_v I__2809 (
            .O(N__29749),
            .I(N__29746));
    Odrv4 I__2808 (
            .O(N__29746),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635 ));
    InMux I__2807 (
            .O(N__29743),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434 ));
    CascadeMux I__2806 (
            .O(N__29740),
            .I(N__29737));
    InMux I__2805 (
            .O(N__29737),
            .I(N__29734));
    LocalMux I__2804 (
            .O(N__29734),
            .I(N__29731));
    Span4Mux_v I__2803 (
            .O(N__29731),
            .I(N__29728));
    Odrv4 I__2802 (
            .O(N__29728),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735 ));
    InMux I__2801 (
            .O(N__29725),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435 ));
    InMux I__2800 (
            .O(N__29722),
            .I(N__29719));
    LocalMux I__2799 (
            .O(N__29719),
            .I(N__29716));
    Span4Mux_v I__2798 (
            .O(N__29716),
            .I(N__29713));
    Odrv4 I__2797 (
            .O(N__29713),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835 ));
    InMux I__2796 (
            .O(N__29710),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436 ));
    InMux I__2795 (
            .O(N__29707),
            .I(N__29704));
    LocalMux I__2794 (
            .O(N__29704),
            .I(N__29701));
    Span4Mux_v I__2793 (
            .O(N__29701),
            .I(N__29698));
    Odrv4 I__2792 (
            .O(N__29698),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935 ));
    InMux I__2791 (
            .O(N__29695),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437 ));
    InMux I__2790 (
            .O(N__29692),
            .I(N__29689));
    LocalMux I__2789 (
            .O(N__29689),
            .I(N__29686));
    Span4Mux_h I__2788 (
            .O(N__29686),
            .I(N__29683));
    Odrv4 I__2787 (
            .O(N__29683),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035 ));
    CascadeMux I__2786 (
            .O(N__29680),
            .I(N__29677));
    InMux I__2785 (
            .O(N__29677),
            .I(N__29669));
    CascadeMux I__2784 (
            .O(N__29676),
            .I(N__29666));
    CascadeMux I__2783 (
            .O(N__29675),
            .I(N__29663));
    CascadeMux I__2782 (
            .O(N__29674),
            .I(N__29659));
    CascadeMux I__2781 (
            .O(N__29673),
            .I(N__29655));
    CascadeMux I__2780 (
            .O(N__29672),
            .I(N__29652));
    LocalMux I__2779 (
            .O(N__29669),
            .I(N__29649));
    InMux I__2778 (
            .O(N__29666),
            .I(N__29646));
    InMux I__2777 (
            .O(N__29663),
            .I(N__29633));
    InMux I__2776 (
            .O(N__29662),
            .I(N__29633));
    InMux I__2775 (
            .O(N__29659),
            .I(N__29633));
    InMux I__2774 (
            .O(N__29658),
            .I(N__29633));
    InMux I__2773 (
            .O(N__29655),
            .I(N__29633));
    InMux I__2772 (
            .O(N__29652),
            .I(N__29633));
    Odrv12 I__2771 (
            .O(N__29649),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831 ));
    LocalMux I__2770 (
            .O(N__29646),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831 ));
    LocalMux I__2769 (
            .O(N__29633),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831 ));
    InMux I__2768 (
            .O(N__29626),
            .I(bfn_9_22_0_));
    InMux I__2767 (
            .O(N__29623),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464 ));
    InMux I__2766 (
            .O(N__29620),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465 ));
    InMux I__2765 (
            .O(N__29617),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466 ));
    InMux I__2764 (
            .O(N__29614),
            .I(bfn_9_20_0_));
    CascadeMux I__2763 (
            .O(N__29611),
            .I(N__29606));
    CascadeMux I__2762 (
            .O(N__29610),
            .I(N__29602));
    CascadeMux I__2761 (
            .O(N__29609),
            .I(N__29598));
    InMux I__2760 (
            .O(N__29606),
            .I(N__29580));
    InMux I__2759 (
            .O(N__29605),
            .I(N__29580));
    InMux I__2758 (
            .O(N__29602),
            .I(N__29580));
    InMux I__2757 (
            .O(N__29601),
            .I(N__29580));
    InMux I__2756 (
            .O(N__29598),
            .I(N__29580));
    InMux I__2755 (
            .O(N__29597),
            .I(N__29580));
    InMux I__2754 (
            .O(N__29596),
            .I(N__29580));
    CascadeMux I__2753 (
            .O(N__29595),
            .I(N__29577));
    LocalMux I__2752 (
            .O(N__29580),
            .I(N__29574));
    InMux I__2751 (
            .O(N__29577),
            .I(N__29571));
    Span4Mux_v I__2750 (
            .O(N__29574),
            .I(N__29566));
    LocalMux I__2749 (
            .O(N__29571),
            .I(N__29566));
    Odrv4 I__2748 (
            .O(N__29566),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834 ));
    InMux I__2747 (
            .O(N__29563),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468 ));
    CascadeMux I__2746 (
            .O(N__29560),
            .I(N__29557));
    InMux I__2745 (
            .O(N__29557),
            .I(N__29554));
    LocalMux I__2744 (
            .O(N__29554),
            .I(N__29548));
    CascadeMux I__2743 (
            .O(N__29553),
            .I(N__29544));
    CascadeMux I__2742 (
            .O(N__29552),
            .I(N__29540));
    CascadeMux I__2741 (
            .O(N__29551),
            .I(N__29536));
    Span4Mux_h I__2740 (
            .O(N__29548),
            .I(N__29528));
    CascadeMux I__2739 (
            .O(N__29547),
            .I(N__29525));
    InMux I__2738 (
            .O(N__29544),
            .I(N__29510));
    InMux I__2737 (
            .O(N__29543),
            .I(N__29510));
    InMux I__2736 (
            .O(N__29540),
            .I(N__29510));
    InMux I__2735 (
            .O(N__29539),
            .I(N__29510));
    InMux I__2734 (
            .O(N__29536),
            .I(N__29510));
    InMux I__2733 (
            .O(N__29535),
            .I(N__29510));
    InMux I__2732 (
            .O(N__29534),
            .I(N__29510));
    CascadeMux I__2731 (
            .O(N__29533),
            .I(N__29507));
    CascadeMux I__2730 (
            .O(N__29532),
            .I(N__29503));
    CascadeMux I__2729 (
            .O(N__29531),
            .I(N__29499));
    Span4Mux_v I__2728 (
            .O(N__29528),
            .I(N__29494));
    InMux I__2727 (
            .O(N__29525),
            .I(N__29491));
    LocalMux I__2726 (
            .O(N__29510),
            .I(N__29488));
    InMux I__2725 (
            .O(N__29507),
            .I(N__29473));
    InMux I__2724 (
            .O(N__29506),
            .I(N__29473));
    InMux I__2723 (
            .O(N__29503),
            .I(N__29473));
    InMux I__2722 (
            .O(N__29502),
            .I(N__29473));
    InMux I__2721 (
            .O(N__29499),
            .I(N__29473));
    InMux I__2720 (
            .O(N__29498),
            .I(N__29473));
    InMux I__2719 (
            .O(N__29497),
            .I(N__29473));
    Sp12to4 I__2718 (
            .O(N__29494),
            .I(N__29468));
    LocalMux I__2717 (
            .O(N__29491),
            .I(N__29468));
    Span4Mux_h I__2716 (
            .O(N__29488),
            .I(N__29465));
    LocalMux I__2715 (
            .O(N__29473),
            .I(N__29462));
    Span12Mux_s8_h I__2714 (
            .O(N__29468),
            .I(N__29459));
    Span4Mux_v I__2713 (
            .O(N__29465),
            .I(N__29454));
    Span4Mux_h I__2712 (
            .O(N__29462),
            .I(N__29454));
    Odrv12 I__2711 (
            .O(N__29459),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840 ));
    Odrv4 I__2710 (
            .O(N__29454),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840 ));
    InMux I__2709 (
            .O(N__29449),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469 ));
    CascadeMux I__2708 (
            .O(N__29446),
            .I(N__29443));
    InMux I__2707 (
            .O(N__29443),
            .I(N__29436));
    CascadeMux I__2706 (
            .O(N__29442),
            .I(N__29433));
    CascadeMux I__2705 (
            .O(N__29441),
            .I(N__29430));
    CascadeMux I__2704 (
            .O(N__29440),
            .I(N__29427));
    CascadeMux I__2703 (
            .O(N__29439),
            .I(N__29423));
    LocalMux I__2702 (
            .O(N__29436),
            .I(N__29418));
    InMux I__2701 (
            .O(N__29433),
            .I(N__29415));
    InMux I__2700 (
            .O(N__29430),
            .I(N__29402));
    InMux I__2699 (
            .O(N__29427),
            .I(N__29402));
    InMux I__2698 (
            .O(N__29426),
            .I(N__29402));
    InMux I__2697 (
            .O(N__29423),
            .I(N__29402));
    InMux I__2696 (
            .O(N__29422),
            .I(N__29402));
    InMux I__2695 (
            .O(N__29421),
            .I(N__29402));
    Span4Mux_v I__2694 (
            .O(N__29418),
            .I(N__29399));
    LocalMux I__2693 (
            .O(N__29415),
            .I(N__29394));
    LocalMux I__2692 (
            .O(N__29402),
            .I(N__29394));
    Span4Mux_v I__2691 (
            .O(N__29399),
            .I(N__29391));
    Span4Mux_h I__2690 (
            .O(N__29394),
            .I(N__29388));
    Odrv4 I__2689 (
            .O(N__29391),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843 ));
    Odrv4 I__2688 (
            .O(N__29388),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843 ));
    InMux I__2687 (
            .O(N__29383),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470 ));
    InMux I__2686 (
            .O(N__29380),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471 ));
    InMux I__2685 (
            .O(N__29377),
            .I(\foc.u_Park_Transform.n16944 ));
    InMux I__2684 (
            .O(N__29374),
            .I(\foc.u_Park_Transform.n16945 ));
    InMux I__2683 (
            .O(N__29371),
            .I(\foc.u_Park_Transform.n16946 ));
    InMux I__2682 (
            .O(N__29368),
            .I(\foc.u_Park_Transform.n775 ));
    InMux I__2681 (
            .O(N__29365),
            .I(bfn_9_19_0_));
    InMux I__2680 (
            .O(N__29362),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460 ));
    InMux I__2679 (
            .O(N__29359),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461 ));
    InMux I__2678 (
            .O(N__29356),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462 ));
    InMux I__2677 (
            .O(N__29353),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463 ));
    InMux I__2676 (
            .O(N__29350),
            .I(\foc.u_Park_Transform.n16935 ));
    InMux I__2675 (
            .O(N__29347),
            .I(\foc.u_Park_Transform.n16936 ));
    InMux I__2674 (
            .O(N__29344),
            .I(\foc.u_Park_Transform.n16937 ));
    InMux I__2673 (
            .O(N__29341),
            .I(\foc.u_Park_Transform.n16938 ));
    InMux I__2672 (
            .O(N__29338),
            .I(\foc.u_Park_Transform.n16939 ));
    InMux I__2671 (
            .O(N__29335),
            .I(\foc.u_Park_Transform.n16940 ));
    InMux I__2670 (
            .O(N__29332),
            .I(\foc.u_Park_Transform.n16941 ));
    InMux I__2669 (
            .O(N__29329),
            .I(bfn_9_16_0_));
    InMux I__2668 (
            .O(N__29326),
            .I(\foc.u_Park_Transform.n16943 ));
    CascadeMux I__2667 (
            .O(N__29323),
            .I(N__29320));
    InMux I__2666 (
            .O(N__29320),
            .I(N__29317));
    LocalMux I__2665 (
            .O(N__29317),
            .I(N__29314));
    Odrv12 I__2664 (
            .O(N__29314),
            .I(\foc.u_Park_Transform.n424_adj_2052 ));
    InMux I__2663 (
            .O(N__29311),
            .I(bfn_9_12_0_));
    InMux I__2662 (
            .O(N__29308),
            .I(N__29305));
    LocalMux I__2661 (
            .O(N__29305),
            .I(N__29302));
    Odrv4 I__2660 (
            .O(N__29302),
            .I(\foc.u_Park_Transform.n473_adj_2050 ));
    InMux I__2659 (
            .O(N__29299),
            .I(\foc.u_Park_Transform.n17126 ));
    InMux I__2658 (
            .O(N__29296),
            .I(\foc.u_Park_Transform.n17127 ));
    InMux I__2657 (
            .O(N__29293),
            .I(\foc.u_Park_Transform.n17128 ));
    CascadeMux I__2656 (
            .O(N__29290),
            .I(N__29285));
    InMux I__2655 (
            .O(N__29289),
            .I(N__29282));
    InMux I__2654 (
            .O(N__29288),
            .I(N__29277));
    InMux I__2653 (
            .O(N__29285),
            .I(N__29277));
    LocalMux I__2652 (
            .O(N__29282),
            .I(N__29272));
    LocalMux I__2651 (
            .O(N__29277),
            .I(N__29272));
    Odrv4 I__2650 (
            .O(N__29272),
            .I(\foc.u_Park_Transform.n522_adj_2046 ));
    InMux I__2649 (
            .O(N__29269),
            .I(\foc.u_Park_Transform.n17129 ));
    InMux I__2648 (
            .O(N__29266),
            .I(\foc.u_Park_Transform.n775_adj_2047 ));
    InMux I__2647 (
            .O(N__29263),
            .I(\foc.u_Park_Transform.n779_adj_2070 ));
    CascadeMux I__2646 (
            .O(N__29260),
            .I(N__29257));
    InMux I__2645 (
            .O(N__29257),
            .I(N__29254));
    LocalMux I__2644 (
            .O(N__29254),
            .I(N__29251));
    Odrv4 I__2643 (
            .O(N__29251),
            .I(\foc.u_Park_Transform.n81 ));
    InMux I__2642 (
            .O(N__29248),
            .I(\foc.u_Park_Transform.n17118 ));
    CascadeMux I__2641 (
            .O(N__29245),
            .I(N__29242));
    InMux I__2640 (
            .O(N__29242),
            .I(N__29239));
    LocalMux I__2639 (
            .O(N__29239),
            .I(N__29236));
    Odrv12 I__2638 (
            .O(N__29236),
            .I(\foc.u_Park_Transform.n130 ));
    InMux I__2637 (
            .O(N__29233),
            .I(\foc.u_Park_Transform.n17119 ));
    InMux I__2636 (
            .O(N__29230),
            .I(N__29227));
    LocalMux I__2635 (
            .O(N__29227),
            .I(N__29224));
    Odrv12 I__2634 (
            .O(N__29224),
            .I(\foc.u_Park_Transform.n179 ));
    InMux I__2633 (
            .O(N__29221),
            .I(\foc.u_Park_Transform.n17120 ));
    CascadeMux I__2632 (
            .O(N__29218),
            .I(N__29215));
    InMux I__2631 (
            .O(N__29215),
            .I(N__29212));
    LocalMux I__2630 (
            .O(N__29212),
            .I(N__29209));
    Odrv12 I__2629 (
            .O(N__29209),
            .I(\foc.u_Park_Transform.n228_adj_2063 ));
    InMux I__2628 (
            .O(N__29206),
            .I(\foc.u_Park_Transform.n17121 ));
    InMux I__2627 (
            .O(N__29203),
            .I(N__29200));
    LocalMux I__2626 (
            .O(N__29200),
            .I(N__29197));
    Odrv4 I__2625 (
            .O(N__29197),
            .I(\foc.u_Park_Transform.n277_adj_2060 ));
    InMux I__2624 (
            .O(N__29194),
            .I(\foc.u_Park_Transform.n17122 ));
    CascadeMux I__2623 (
            .O(N__29191),
            .I(N__29188));
    InMux I__2622 (
            .O(N__29188),
            .I(N__29185));
    LocalMux I__2621 (
            .O(N__29185),
            .I(N__29182));
    Odrv4 I__2620 (
            .O(N__29182),
            .I(\foc.u_Park_Transform.n326_adj_2056 ));
    InMux I__2619 (
            .O(N__29179),
            .I(\foc.u_Park_Transform.n17123 ));
    InMux I__2618 (
            .O(N__29176),
            .I(N__29173));
    LocalMux I__2617 (
            .O(N__29173),
            .I(N__29170));
    Odrv4 I__2616 (
            .O(N__29170),
            .I(\foc.u_Park_Transform.n375_adj_2055 ));
    InMux I__2615 (
            .O(N__29167),
            .I(\foc.u_Park_Transform.n17124 ));
    InMux I__2614 (
            .O(N__29164),
            .I(\foc.u_Park_Transform.n17108 ));
    InMux I__2613 (
            .O(N__29161),
            .I(\foc.u_Park_Transform.n17109 ));
    InMux I__2612 (
            .O(N__29158),
            .I(\foc.u_Park_Transform.n17110 ));
    InMux I__2611 (
            .O(N__29155),
            .I(\foc.u_Park_Transform.n17111 ));
    InMux I__2610 (
            .O(N__29152),
            .I(\foc.u_Park_Transform.n17112 ));
    InMux I__2609 (
            .O(N__29149),
            .I(\foc.u_Park_Transform.n17113 ));
    InMux I__2608 (
            .O(N__29146),
            .I(bfn_9_10_0_));
    InMux I__2607 (
            .O(N__29143),
            .I(\foc.u_Park_Transform.n17115 ));
    InMux I__2606 (
            .O(N__29140),
            .I(\foc.u_Park_Transform.n17116 ));
    InMux I__2605 (
            .O(N__29137),
            .I(N__29134));
    LocalMux I__2604 (
            .O(N__29134),
            .I(N__29131));
    Odrv4 I__2603 (
            .O(N__29131),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744 ));
    CascadeMux I__2602 (
            .O(N__29128),
            .I(N__29125));
    InMux I__2601 (
            .O(N__29125),
            .I(N__29122));
    LocalMux I__2600 (
            .O(N__29122),
            .I(N__29119));
    Odrv12 I__2599 (
            .O(N__29119),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841 ));
    InMux I__2598 (
            .O(N__29116),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465 ));
    CascadeMux I__2597 (
            .O(N__29113),
            .I(N__29110));
    InMux I__2596 (
            .O(N__29110),
            .I(N__29107));
    LocalMux I__2595 (
            .O(N__29107),
            .I(N__29104));
    Odrv4 I__2594 (
            .O(N__29104),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844 ));
    InMux I__2593 (
            .O(N__29101),
            .I(N__29098));
    LocalMux I__2592 (
            .O(N__29098),
            .I(N__29095));
    Odrv12 I__2591 (
            .O(N__29095),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941 ));
    InMux I__2590 (
            .O(N__29092),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466 ));
    InMux I__2589 (
            .O(N__29089),
            .I(N__29086));
    LocalMux I__2588 (
            .O(N__29086),
            .I(N__29083));
    Odrv4 I__2587 (
            .O(N__29083),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944 ));
    InMux I__2586 (
            .O(N__29080),
            .I(N__29077));
    LocalMux I__2585 (
            .O(N__29077),
            .I(N__29074));
    Odrv12 I__2584 (
            .O(N__29074),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041 ));
    InMux I__2583 (
            .O(N__29071),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467 ));
    InMux I__2582 (
            .O(N__29068),
            .I(N__29065));
    LocalMux I__2581 (
            .O(N__29065),
            .I(N__29062));
    Odrv4 I__2580 (
            .O(N__29062),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044 ));
    InMux I__2579 (
            .O(N__29059),
            .I(N__29056));
    LocalMux I__2578 (
            .O(N__29056),
            .I(N__29053));
    Odrv12 I__2577 (
            .O(N__29053),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141 ));
    InMux I__2576 (
            .O(N__29050),
            .I(bfn_7_26_0_));
    InMux I__2575 (
            .O(N__29047),
            .I(N__29044));
    LocalMux I__2574 (
            .O(N__29044),
            .I(N__29041));
    Odrv4 I__2573 (
            .O(N__29041),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144 ));
    InMux I__2572 (
            .O(N__29038),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469 ));
    InMux I__2571 (
            .O(N__29035),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256 ));
    InMux I__2570 (
            .O(N__29032),
            .I(\foc.u_Park_Transform.n17107 ));
    InMux I__2569 (
            .O(N__29029),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477 ));
    InMux I__2568 (
            .O(N__29026),
            .I(bfn_7_24_0_));
    InMux I__2567 (
            .O(N__29023),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479 ));
    InMux I__2566 (
            .O(N__29020),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260 ));
    InMux I__2565 (
            .O(N__29017),
            .I(N__29014));
    LocalMux I__2564 (
            .O(N__29014),
            .I(N__29011));
    Span4Mux_v I__2563 (
            .O(N__29011),
            .I(N__29008));
    Odrv4 I__2562 (
            .O(N__29008),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341 ));
    InMux I__2561 (
            .O(N__29005),
            .I(N__29002));
    LocalMux I__2560 (
            .O(N__29002),
            .I(N__28999));
    Odrv4 I__2559 (
            .O(N__28999),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344 ));
    CascadeMux I__2558 (
            .O(N__28996),
            .I(N__28993));
    InMux I__2557 (
            .O(N__28993),
            .I(N__28990));
    LocalMux I__2556 (
            .O(N__28990),
            .I(N__28987));
    Span4Mux_v I__2555 (
            .O(N__28987),
            .I(N__28984));
    Odrv4 I__2554 (
            .O(N__28984),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441 ));
    InMux I__2553 (
            .O(N__28981),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461 ));
    CascadeMux I__2552 (
            .O(N__28978),
            .I(N__28975));
    InMux I__2551 (
            .O(N__28975),
            .I(N__28972));
    LocalMux I__2550 (
            .O(N__28972),
            .I(N__28969));
    Odrv4 I__2549 (
            .O(N__28969),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444 ));
    InMux I__2548 (
            .O(N__28966),
            .I(N__28963));
    LocalMux I__2547 (
            .O(N__28963),
            .I(N__28960));
    Sp12to4 I__2546 (
            .O(N__28960),
            .I(N__28957));
    Odrv12 I__2545 (
            .O(N__28957),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541 ));
    InMux I__2544 (
            .O(N__28954),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462 ));
    InMux I__2543 (
            .O(N__28951),
            .I(N__28948));
    LocalMux I__2542 (
            .O(N__28948),
            .I(N__28945));
    Odrv12 I__2541 (
            .O(N__28945),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544 ));
    CascadeMux I__2540 (
            .O(N__28942),
            .I(N__28939));
    InMux I__2539 (
            .O(N__28939),
            .I(N__28936));
    LocalMux I__2538 (
            .O(N__28936),
            .I(N__28933));
    Odrv12 I__2537 (
            .O(N__28933),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641 ));
    InMux I__2536 (
            .O(N__28930),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463 ));
    CascadeMux I__2535 (
            .O(N__28927),
            .I(N__28924));
    InMux I__2534 (
            .O(N__28924),
            .I(N__28921));
    LocalMux I__2533 (
            .O(N__28921),
            .I(N__28918));
    Odrv12 I__2532 (
            .O(N__28918),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644 ));
    InMux I__2531 (
            .O(N__28915),
            .I(N__28912));
    LocalMux I__2530 (
            .O(N__28912),
            .I(N__28909));
    Odrv12 I__2529 (
            .O(N__28909),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741 ));
    InMux I__2528 (
            .O(N__28906),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464 ));
    InMux I__2527 (
            .O(N__28903),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459 ));
    InMux I__2526 (
            .O(N__28900),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252 ));
    InMux I__2525 (
            .O(N__28897),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471 ));
    InMux I__2524 (
            .O(N__28894),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472 ));
    InMux I__2523 (
            .O(N__28891),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473 ));
    InMux I__2522 (
            .O(N__28888),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474 ));
    InMux I__2521 (
            .O(N__28885),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475 ));
    InMux I__2520 (
            .O(N__28882),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476 ));
    CascadeMux I__2519 (
            .O(N__28879),
            .I(N__28876));
    InMux I__2518 (
            .O(N__28876),
            .I(N__28873));
    LocalMux I__2517 (
            .O(N__28873),
            .I(N__28870));
    Odrv4 I__2516 (
            .O(N__28870),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438 ));
    InMux I__2515 (
            .O(N__28867),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451 ));
    InMux I__2514 (
            .O(N__28864),
            .I(N__28861));
    LocalMux I__2513 (
            .O(N__28861),
            .I(N__28858));
    Odrv4 I__2512 (
            .O(N__28858),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538 ));
    InMux I__2511 (
            .O(N__28855),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452 ));
    CascadeMux I__2510 (
            .O(N__28852),
            .I(N__28849));
    InMux I__2509 (
            .O(N__28849),
            .I(N__28846));
    LocalMux I__2508 (
            .O(N__28846),
            .I(N__28843));
    Odrv4 I__2507 (
            .O(N__28843),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638 ));
    InMux I__2506 (
            .O(N__28840),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453 ));
    InMux I__2505 (
            .O(N__28837),
            .I(N__28834));
    LocalMux I__2504 (
            .O(N__28834),
            .I(N__28831));
    Odrv4 I__2503 (
            .O(N__28831),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738 ));
    InMux I__2502 (
            .O(N__28828),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454 ));
    CascadeMux I__2501 (
            .O(N__28825),
            .I(N__28822));
    InMux I__2500 (
            .O(N__28822),
            .I(N__28819));
    LocalMux I__2499 (
            .O(N__28819),
            .I(N__28816));
    Odrv4 I__2498 (
            .O(N__28816),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838 ));
    InMux I__2497 (
            .O(N__28813),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455 ));
    InMux I__2496 (
            .O(N__28810),
            .I(N__28807));
    LocalMux I__2495 (
            .O(N__28807),
            .I(N__28804));
    Odrv4 I__2494 (
            .O(N__28804),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938 ));
    InMux I__2493 (
            .O(N__28801),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456 ));
    InMux I__2492 (
            .O(N__28798),
            .I(N__28795));
    LocalMux I__2491 (
            .O(N__28795),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038 ));
    InMux I__2490 (
            .O(N__28792),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457 ));
    InMux I__2489 (
            .O(N__28789),
            .I(N__28786));
    LocalMux I__2488 (
            .O(N__28786),
            .I(N__28783));
    Odrv4 I__2487 (
            .O(N__28783),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138 ));
    InMux I__2486 (
            .O(N__28780),
            .I(bfn_7_22_0_));
    InMux I__2485 (
            .O(N__28777),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444 ));
    InMux I__2484 (
            .O(N__28774),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445 ));
    InMux I__2483 (
            .O(N__28771),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446 ));
    InMux I__2482 (
            .O(N__28768),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447 ));
    InMux I__2481 (
            .O(N__28765),
            .I(bfn_7_20_0_));
    InMux I__2480 (
            .O(N__28762),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449 ));
    InMux I__2479 (
            .O(N__28759),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248 ));
    CascadeMux I__2478 (
            .O(N__28756),
            .I(N__28752));
    InMux I__2477 (
            .O(N__28755),
            .I(N__28741));
    InMux I__2476 (
            .O(N__28752),
            .I(N__28741));
    InMux I__2475 (
            .O(N__28751),
            .I(N__28741));
    InMux I__2474 (
            .O(N__28750),
            .I(N__28741));
    LocalMux I__2473 (
            .O(N__28741),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490 ));
    InMux I__2472 (
            .O(N__28738),
            .I(N__28735));
    LocalMux I__2471 (
            .O(N__28735),
            .I(N__28732));
    Odrv4 I__2470 (
            .O(N__28732),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338 ));
    InMux I__2469 (
            .O(N__28729),
            .I(N__28726));
    LocalMux I__2468 (
            .O(N__28726),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175 ));
    InMux I__2467 (
            .O(N__28723),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346 ));
    InMux I__2466 (
            .O(N__28720),
            .I(N__28717));
    LocalMux I__2465 (
            .O(N__28717),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174 ));
    InMux I__2464 (
            .O(N__28714),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347 ));
    InMux I__2463 (
            .O(N__28711),
            .I(N__28708));
    LocalMux I__2462 (
            .O(N__28708),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173 ));
    InMux I__2461 (
            .O(N__28705),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348 ));
    InMux I__2460 (
            .O(N__28702),
            .I(N__28699));
    LocalMux I__2459 (
            .O(N__28699),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172 ));
    InMux I__2458 (
            .O(N__28696),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349 ));
    InMux I__2457 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__2456 (
            .O(N__28690),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177 ));
    InMux I__2455 (
            .O(N__28687),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441 ));
    InMux I__2454 (
            .O(N__28684),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442 ));
    InMux I__2453 (
            .O(N__28681),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443 ));
    InMux I__2452 (
            .O(N__28678),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332 ));
    InMux I__2451 (
            .O(N__28675),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333 ));
    InMux I__2450 (
            .O(N__28672),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334 ));
    InMux I__2449 (
            .O(N__28669),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335 ));
    InMux I__2448 (
            .O(N__28666),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336 ));
    InMux I__2447 (
            .O(N__28663),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344 ));
    InMux I__2446 (
            .O(N__28660),
            .I(N__28657));
    LocalMux I__2445 (
            .O(N__28657),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176 ));
    InMux I__2444 (
            .O(N__28654),
            .I(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345 ));
    IoInMux I__2443 (
            .O(N__28651),
            .I(N__28648));
    LocalMux I__2442 (
            .O(N__28648),
            .I(N__28645));
    Span12Mux_s8_h I__2441 (
            .O(N__28645),
            .I(N__28642));
    Span12Mux_v I__2440 (
            .O(N__28642),
            .I(N__28639));
    Odrv12 I__2439 (
            .O(N__28639),
            .I(pin3_clk_16mhz_pad_gb_input));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17090 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\foc.u_Park_Transform.n16907 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_19_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_21_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18151 ),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18159 ),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17964 ),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17972 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15727 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15735 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15743 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_18_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_26_0_));
    defparam IN_MUX_bfv_18_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_27_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18361 ),
            .carryinitout(bfn_18_27_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_19_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_18_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17718 ),
            .carryinitout(bfn_19_18_0_));
    defparam IN_MUX_bfv_19_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_19_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17726 ),
            .carryinitout(bfn_19_19_0_));
    defparam IN_MUX_bfv_20_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_14_0_));
    defparam IN_MUX_bfv_20_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_15_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17512 ),
            .carryinitout(bfn_20_15_0_));
    defparam IN_MUX_bfv_20_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_16_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17520 ),
            .carryinitout(bfn_20_16_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15782 ),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15790 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15798 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_19_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_9_0_));
    defparam IN_MUX_bfv_19_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_10_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17934 ),
            .carryinitout(bfn_19_10_0_));
    defparam IN_MUX_bfv_6_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357 ),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478 ),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468 ),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\foc.u_Park_Transform.n15755 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\foc.u_Park_Transform.n15763 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\foc.u_Park_Transform.n15771 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\foc.u_Park_Transform.n17284 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\foc.u_Park_Transform.n17292 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17300 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n16922 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\foc.u_Park_Transform.n16931 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n16942 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n16955 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n16970 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n16985 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\foc.u_Park_Transform.n17000 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\foc.u_Park_Transform.n17015 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\foc.u_Park_Transform.n17030 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\foc.u_Park_Transform.n17045 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n17060 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\foc.u_Park_Transform.n17075 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17105 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17114 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17125 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17138 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17153 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17168 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17183 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17198 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17213 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17228 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\foc.u_Park_Transform.n17243 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\foc.u_Park_Transform.n17258 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17734 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17863 ),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17663 ),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18114 ),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18099 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18084 ),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18069 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18054 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18039 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_16_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18024 ),
            .carryinitout(bfn_16_26_0_));
    defparam IN_MUX_bfv_16_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_27_0_));
    defparam IN_MUX_bfv_16_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_28_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18009 ),
            .carryinitout(bfn_16_28_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17994 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_21_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_23_0_));
    defparam IN_MUX_bfv_21_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15920 ),
            .carryinitout(bfn_21_24_0_));
    defparam IN_MUX_bfv_21_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_25_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15928 ),
            .carryinitout(bfn_21_25_0_));
    defparam IN_MUX_bfv_21_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15936 ),
            .carryinitout(bfn_21_26_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15890 ),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15898 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_18_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_25_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15906 ),
            .carryinitout(bfn_18_25_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18376 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_19_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_26_0_));
    defparam IN_MUX_bfv_19_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_27_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18346 ),
            .carryinitout(bfn_19_27_0_));
    defparam IN_MUX_bfv_19_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_28_0_));
    defparam IN_MUX_bfv_19_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_29_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18331 ),
            .carryinitout(bfn_19_29_0_));
    defparam IN_MUX_bfv_20_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_28_0_));
    defparam IN_MUX_bfv_20_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_29_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18316 ),
            .carryinitout(bfn_20_29_0_));
    defparam IN_MUX_bfv_21_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_28_0_));
    defparam IN_MUX_bfv_21_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_29_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18301 ),
            .carryinitout(bfn_21_29_0_));
    defparam IN_MUX_bfv_22_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_28_0_));
    defparam IN_MUX_bfv_22_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_29_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18286 ),
            .carryinitout(bfn_22_29_0_));
    defparam IN_MUX_bfv_23_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_27_0_));
    defparam IN_MUX_bfv_23_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_28_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18271 ),
            .carryinitout(bfn_23_28_0_));
    defparam IN_MUX_bfv_23_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_25_0_));
    defparam IN_MUX_bfv_23_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18256 ),
            .carryinitout(bfn_23_26_0_));
    defparam IN_MUX_bfv_22_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_25_0_));
    defparam IN_MUX_bfv_22_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18241 ),
            .carryinitout(bfn_22_26_0_));
    defparam IN_MUX_bfv_20_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_25_0_));
    defparam IN_MUX_bfv_20_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_26_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18226 ),
            .carryinitout(bfn_20_26_0_));
    defparam IN_MUX_bfv_20_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_23_0_));
    defparam IN_MUX_bfv_20_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_24_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18211 ),
            .carryinitout(bfn_20_24_0_));
    defparam IN_MUX_bfv_19_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_24_0_));
    defparam IN_MUX_bfv_19_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_25_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18196 ),
            .carryinitout(bfn_19_25_0_));
    defparam IN_MUX_bfv_21_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_21_0_));
    defparam IN_MUX_bfv_21_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_22_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18181 ),
            .carryinitout(bfn_21_22_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18142 ),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_18_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_5_0_));
    defparam IN_MUX_bfv_18_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_6_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17273 ),
            .carryinitout(bfn_18_6_0_));
    defparam IN_MUX_bfv_20_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_5_0_));
    defparam IN_MUX_bfv_20_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_6_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18129 ),
            .carryinitout(bfn_20_6_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17648 ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17633 ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_20_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_7_0_));
    defparam IN_MUX_bfv_20_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_8_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17618 ),
            .carryinitout(bfn_20_8_0_));
    defparam IN_MUX_bfv_21_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_7_0_));
    defparam IN_MUX_bfv_21_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_8_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17603 ),
            .carryinitout(bfn_21_8_0_));
    defparam IN_MUX_bfv_20_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_9_0_));
    defparam IN_MUX_bfv_20_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_10_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17588 ),
            .carryinitout(bfn_20_10_0_));
    defparam IN_MUX_bfv_21_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_9_0_));
    defparam IN_MUX_bfv_21_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_10_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17573 ),
            .carryinitout(bfn_21_10_0_));
    defparam IN_MUX_bfv_21_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_11_0_));
    defparam IN_MUX_bfv_21_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_12_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17558 ),
            .carryinitout(bfn_21_12_0_));
    defparam IN_MUX_bfv_22_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_11_0_));
    defparam IN_MUX_bfv_22_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_12_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17543 ),
            .carryinitout(bfn_22_12_0_));
    defparam IN_MUX_bfv_23_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_11_0_));
    defparam IN_MUX_bfv_23_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_12_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17528 ),
            .carryinitout(bfn_23_12_0_));
    defparam IN_MUX_bfv_22_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_19_0_));
    defparam IN_MUX_bfv_22_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_20_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15980 ),
            .carryinitout(bfn_22_20_0_));
    defparam IN_MUX_bfv_22_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_21_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15988 ),
            .carryinitout(bfn_22_21_0_));
    defparam IN_MUX_bfv_22_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_22_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15996 ),
            .carryinitout(bfn_22_22_0_));
    defparam IN_MUX_bfv_24_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_16_0_));
    defparam IN_MUX_bfv_24_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_17_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_24_17_0_));
    defparam IN_MUX_bfv_24_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_18_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_24_18_0_));
    defparam IN_MUX_bfv_24_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_19_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15588 ),
            .carryinitout(bfn_24_19_0_));
    defparam IN_MUX_bfv_24_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_20_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15596 ),
            .carryinitout(bfn_24_20_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17949 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_19_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_11_0_));
    defparam IN_MUX_bfv_19_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_12_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17919 ),
            .carryinitout(bfn_19_12_0_));
    defparam IN_MUX_bfv_20_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_11_0_));
    defparam IN_MUX_bfv_20_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_12_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17904 ),
            .carryinitout(bfn_20_12_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17889 ),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17874 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17848 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17833 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_19_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_13_0_));
    defparam IN_MUX_bfv_19_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_14_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17818 ),
            .carryinitout(bfn_19_14_0_));
    defparam IN_MUX_bfv_19_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_15_0_));
    defparam IN_MUX_bfv_19_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_16_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17803 ),
            .carryinitout(bfn_19_16_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17788 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17773 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17758 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_21_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_17_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17743 ),
            .carryinitout(bfn_21_18_0_));
    ICE_GB pin3_clk_16mhz_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__28651),
            .GLOBALBUFFEROUTPUT(pin3_clk_16mhz_N));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_2_lut_LC_6_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_2_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_2_lut_LC_6_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_2_lut_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(N__31562),
            .in2(N__32765),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7897 ),
            .ltout(),
            .carryin(bfn_6_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_3_lut_LC_6_20_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_3_lut_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_3_lut_LC_6_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_3_lut_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(N__28750),
            .in2(_gnd_net_),
            .in3(N__28678),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8176 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17332 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_4_lut_LC_6_20_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_4_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_4_lut_LC_6_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_4_lut_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(N__31563),
            .in2(N__32766),
            .in3(N__28675),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8175 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17333 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_5_lut_LC_6_20_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_5_lut_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_5_lut_LC_6_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_5_lut_LC_6_20_3  (
            .in0(_gnd_net_),
            .in1(N__28751),
            .in2(N__31573),
            .in3(N__28672),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8174 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17334 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_6_lut_LC_6_20_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_6_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_6_lut_LC_6_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_6_lut_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__31567),
            .in2(N__28756),
            .in3(N__28669),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8173 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17335 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17336 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_7_lut_LC_6_20_5 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_7_lut_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_7_lut_LC_6_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_7_lut_LC_6_20_5  (
            .in0(N__31568),
            .in1(N__28755),
            .in2(_gnd_net_),
            .in3(N__28666),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_2_lut_LC_6_21_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_2_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_2_lut_LC_6_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_2_lut_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(N__31547),
            .in2(N__32799),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7554 ),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_3_lut_LC_6_21_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_3_lut_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_3_lut_LC_6_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_3_lut_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(N__28693),
            .in2(_gnd_net_),
            .in3(N__28663),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7896 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17344 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_4_lut_LC_6_21_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_4_lut_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_4_lut_LC_6_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_4_lut_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(N__28660),
            .in2(N__31571),
            .in3(N__28654),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7895 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17345 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_5_lut_LC_6_21_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_5_lut_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_5_lut_LC_6_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_5_lut_LC_6_21_3  (
            .in0(_gnd_net_),
            .in1(N__28729),
            .in2(N__31569),
            .in3(N__28723),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7894 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17346 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_6_lut_LC_6_21_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_6_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_6_lut_LC_6_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_6_lut_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__28720),
            .in2(N__31572),
            .in3(N__28714),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7893 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17347 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_7_lut_LC_6_21_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_7_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_7_lut_LC_6_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_7_lut_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(N__28711),
            .in2(N__31570),
            .in3(N__28705),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7892 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17348 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17349 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_8_lut_LC_6_21_6 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_8_lut_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_8_lut_LC_6_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6236_8_lut_LC_6_21_6  (
            .in0(N__28702),
            .in1(N__31554),
            .in2(_gnd_net_),
            .in3(N__28696),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_2_lut_LC_6_21_7 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_2_lut_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_2_lut_LC_6_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_6484_2_lut_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(N__31561),
            .in2(_gnd_net_),
            .in3(N__32783),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_2_lut_LC_7_19_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_2_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_2_lut_LC_7_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_2_lut_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__29596),
            .in2(N__32796),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2335 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_3_lut_LC_7_19_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_3_lut_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_3_lut_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_3_lut_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__28738),
            .in2(_gnd_net_),
            .in3(N__28687),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2435 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17441 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_4_lut_LC_7_19_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_4_lut_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_4_lut_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_4_lut_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__29597),
            .in2(N__28879),
            .in3(N__28684),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2535 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17442 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_5_lut_LC_7_19_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_5_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_5_lut_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_5_lut_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__28864),
            .in2(N__29609),
            .in3(N__28681),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2635 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17443 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_6_lut_LC_7_19_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_6_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_6_lut_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_6_lut_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__29601),
            .in2(N__28852),
            .in3(N__28777),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2735 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17444 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_7_lut_LC_7_19_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_7_lut_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_7_lut_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_7_lut_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__28837),
            .in2(N__29610),
            .in3(N__28774),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2835 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17445 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_8_lut_LC_7_19_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_8_lut_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_8_lut_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_8_lut_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__29605),
            .in2(N__28825),
            .in3(N__28771),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2935 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17446 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_9_lut_LC_7_19_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_9_lut_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_9_lut_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_9_lut_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__28810),
            .in2(N__29611),
            .in3(N__28768),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3035 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17447 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17448 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_10_lut_LC_7_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_10_lut_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_10_lut_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_10_lut_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__28798),
            .in2(N__29595),
            .in3(N__28765),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3135 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_11_lut_LC_7_20_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_11_lut_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_11_lut_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2272_11_lut_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__28789),
            .in2(_gnd_net_),
            .in3(N__28762),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3247 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17449 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_LUT4_0_LC_7_20_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_LUT4_0_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_LUT4_0_LC_7_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_LUT4_0_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28759),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3248_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.i13555_2_lut_LC_7_20_4 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.i13555_2_lut_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.i13555_2_lut_LC_7_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.i13555_2_lut_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__32728),
            .in2(_gnd_net_),
            .in3(N__44911),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n8490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_2_lut_LC_7_21_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_2_lut_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_2_lut_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_2_lut_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__29497),
            .in2(N__32797),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2338 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_3_lut_LC_7_21_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_3_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_3_lut_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_3_lut_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__29017),
            .in2(_gnd_net_),
            .in3(N__28867),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2438 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17451 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_4_lut_LC_7_21_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_4_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_4_lut_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_4_lut_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__29498),
            .in2(N__28996),
            .in3(N__28855),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2538 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17452 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_5_lut_LC_7_21_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_5_lut_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_5_lut_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_5_lut_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__28966),
            .in2(N__29531),
            .in3(N__28840),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2638 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17453 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_6_lut_LC_7_21_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_6_lut_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_6_lut_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_6_lut_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__29502),
            .in2(N__28942),
            .in3(N__28828),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2738 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17454 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_7_lut_LC_7_21_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_7_lut_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_7_lut_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_7_lut_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__28915),
            .in2(N__29532),
            .in3(N__28813),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2838 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17455 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_8_lut_LC_7_21_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_8_lut_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_8_lut_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_8_lut_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__29506),
            .in2(N__29128),
            .in3(N__28801),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2938 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17456 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_9_lut_LC_7_21_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_9_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_9_lut_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_9_lut_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__29101),
            .in2(N__29533),
            .in3(N__28792),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3038 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17457 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17458 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_10_lut_LC_7_22_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_10_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_10_lut_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_10_lut_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__29080),
            .in2(N__29547),
            .in3(N__28780),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3138 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_11_lut_LC_7_22_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_11_lut_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_11_lut_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2273_11_lut_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__29059),
            .in2(_gnd_net_),
            .in3(N__28903),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3251 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17459 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_LUT4_0_LC_7_22_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_LUT4_0_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_LUT4_0_LC_7_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_LUT4_0_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28900),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3252_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_2_lut_LC_7_23_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_2_lut_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_2_lut_LC_7_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_2_lut_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__29421),
            .in2(N__32800),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2344 ),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_3_lut_LC_7_23_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_3_lut_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_3_lut_LC_7_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_3_lut_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__30034),
            .in2(_gnd_net_),
            .in3(N__28897),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2444 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17471 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_4_lut_LC_7_23_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_4_lut_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_4_lut_LC_7_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_4_lut_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__29422),
            .in2(N__30016),
            .in3(N__28894),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2544 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17472 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_5_lut_LC_7_23_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_5_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_5_lut_LC_7_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_5_lut_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__29998),
            .in2(N__29439),
            .in3(N__28891),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2644 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17473 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_6_lut_LC_7_23_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_6_lut_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_6_lut_LC_7_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_6_lut_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__29426),
            .in2(N__29983),
            .in3(N__28888),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2744 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17474 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_7_lut_LC_7_23_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_7_lut_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_7_lut_LC_7_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_7_lut_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__29965),
            .in2(N__29440),
            .in3(N__28885),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2844 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17475 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_8_lut_LC_7_23_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_8_lut_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_8_lut_LC_7_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_8_lut_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(N__29950),
            .in2(N__29442),
            .in3(N__28882),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2944 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17476 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_9_lut_LC_7_23_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_9_lut_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_9_lut_LC_7_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_9_lut_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(N__29935),
            .in2(N__29441),
            .in3(N__29029),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3044 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17477 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17478 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_10_lut_LC_7_24_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_10_lut_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_10_lut_LC_7_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_10_lut_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__30094),
            .in2(N__29446),
            .in3(N__29026),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3144 ),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_11_lut_LC_7_24_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_11_lut_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_11_lut_LC_7_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2275_11_lut_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(N__30082),
            .in2(_gnd_net_),
            .in3(N__29023),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3259 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17479 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_LUT4_0_LC_7_24_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_LUT4_0_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_LUT4_0_LC_7_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_LUT4_0_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29020),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3260_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_2_lut_LC_7_25_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_2_lut_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_2_lut_LC_7_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_2_lut_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__29534),
            .in2(N__32806),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2341 ),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_3_lut_LC_7_25_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_3_lut_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_3_lut_LC_7_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_3_lut_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__29005),
            .in2(_gnd_net_),
            .in3(N__28981),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2441 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17461 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_4_lut_LC_7_25_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_4_lut_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_4_lut_LC_7_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_4_lut_LC_7_25_2  (
            .in0(_gnd_net_),
            .in1(N__29535),
            .in2(N__28978),
            .in3(N__28954),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2541 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17462 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_5_lut_LC_7_25_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_5_lut_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_5_lut_LC_7_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_5_lut_LC_7_25_3  (
            .in0(_gnd_net_),
            .in1(N__28951),
            .in2(N__29551),
            .in3(N__28930),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2641 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17463 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_6_lut_LC_7_25_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_6_lut_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_6_lut_LC_7_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_6_lut_LC_7_25_4  (
            .in0(_gnd_net_),
            .in1(N__29539),
            .in2(N__28927),
            .in3(N__28906),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2741 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17464 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_7_lut_LC_7_25_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_7_lut_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_7_lut_LC_7_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_7_lut_LC_7_25_5  (
            .in0(_gnd_net_),
            .in1(N__29137),
            .in2(N__29552),
            .in3(N__29116),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2841 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17465 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_8_lut_LC_7_25_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_8_lut_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_8_lut_LC_7_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_8_lut_LC_7_25_6  (
            .in0(_gnd_net_),
            .in1(N__29543),
            .in2(N__29113),
            .in3(N__29092),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2941 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17466 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_9_lut_LC_7_25_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_9_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_9_lut_LC_7_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_9_lut_LC_7_25_7  (
            .in0(_gnd_net_),
            .in1(N__29089),
            .in2(N__29553),
            .in3(N__29071),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3041 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17467 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17468 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_10_lut_LC_7_26_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_10_lut_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_10_lut_LC_7_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_10_lut_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(N__29068),
            .in2(N__29560),
            .in3(N__29050),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3141 ),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_11_lut_LC_7_26_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_11_lut_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_11_lut_LC_7_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2274_11_lut_LC_7_26_1  (
            .in0(_gnd_net_),
            .in1(N__29047),
            .in2(_gnd_net_),
            .in3(N__29038),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3255 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17469 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_LUT4_0_LC_7_26_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_LUT4_0_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_LUT4_0_LC_7_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_LUT4_0_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29035),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3256_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_2_lut_LC_9_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_2_lut_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_2_lut_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_2_lut_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__31747),
            .in2(N__30850),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n81 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\foc.u_Park_Transform.n17107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_3_lut_LC_9_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_3_lut_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_3_lut_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_3_lut_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__30844),
            .in2(N__31375),
            .in3(N__29032),
            .lcout(\foc.u_Park_Transform.n130 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17107 ),
            .carryout(\foc.u_Park_Transform.n17108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_4_lut_LC_9_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_4_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_4_lut_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_4_lut_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__30796),
            .in2(N__31363),
            .in3(N__29164),
            .lcout(\foc.u_Park_Transform.n179 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17108 ),
            .carryout(\foc.u_Park_Transform.n17109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_5_lut_LC_9_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_5_lut_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_5_lut_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_5_lut_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__31897),
            .in2(N__30837),
            .in3(N__29161),
            .lcout(\foc.u_Park_Transform.n228_adj_2063 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17109 ),
            .carryout(\foc.u_Park_Transform.n17110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_6_lut_LC_9_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_6_lut_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_6_lut_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_6_lut_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__30800),
            .in2(N__31885),
            .in3(N__29158),
            .lcout(\foc.u_Park_Transform.n277_adj_2060 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17110 ),
            .carryout(\foc.u_Park_Transform.n17111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_7_lut_LC_9_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_7_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_7_lut_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_7_lut_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__31870),
            .in2(N__30838),
            .in3(N__29155),
            .lcout(\foc.u_Park_Transform.n326_adj_2056 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17111 ),
            .carryout(\foc.u_Park_Transform.n17112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_8_lut_LC_9_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_8_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_8_lut_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_8_lut_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__30804),
            .in2(N__31855),
            .in3(N__29152),
            .lcout(\foc.u_Park_Transform.n375_adj_2055 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17112 ),
            .carryout(\foc.u_Park_Transform.n17113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_9_lut_LC_9_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_9_lut_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_9_lut_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_9_lut_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__31837),
            .in2(N__30839),
            .in3(N__29149),
            .lcout(\foc.u_Park_Transform.n424_adj_2052 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17113 ),
            .carryout(\foc.u_Park_Transform.n17114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_10_lut_LC_9_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_10_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_10_lut_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_10_lut_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__30808),
            .in2(N__31824),
            .in3(N__29146),
            .lcout(\foc.u_Park_Transform.n473_adj_2050 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\foc.u_Park_Transform.n17115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_11_lut_LC_9_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_11_lut_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_11_lut_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_11_lut_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__31820),
            .in2(N__30840),
            .in3(N__29143),
            .lcout(\foc.u_Park_Transform.n522_adj_2046 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17115 ),
            .carryout(\foc.u_Park_Transform.n17116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_12_lut_LC_9_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_12_lut_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_12_lut_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_571_12_lut_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__30687),
            .in2(N__31825),
            .in3(N__29140),
            .lcout(\foc.u_Park_Transform.n778_adj_2068 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17116 ),
            .carryout(\foc.u_Park_Transform.n779_adj_2070 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n779_adj_2070_THRU_LUT4_0_LC_9_10_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n779_adj_2070_THRU_LUT4_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n779_adj_2070_THRU_LUT4_0_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n779_adj_2070_THRU_LUT4_0_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29263),
            .lcout(\foc.u_Park_Transform.n779_adj_2070_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_2_lut_LC_9_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_2_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_2_lut_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_2_lut_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__30764),
            .in2(N__32369),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n78 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\foc.u_Park_Transform.n17118 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_3_lut_LC_9_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_3_lut_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_3_lut_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_3_lut_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__32330),
            .in2(N__29260),
            .in3(N__29248),
            .lcout(\foc.u_Park_Transform.n127 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17118 ),
            .carryout(\foc.u_Park_Transform.n17119 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_4_lut_LC_9_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_4_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_4_lut_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_4_lut_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__32331),
            .in2(N__29245),
            .in3(N__29233),
            .lcout(\foc.u_Park_Transform.n176 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17119 ),
            .carryout(\foc.u_Park_Transform.n17120 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_5_lut_LC_9_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_5_lut_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_5_lut_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_5_lut_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__29230),
            .in2(N__32370),
            .in3(N__29221),
            .lcout(\foc.u_Park_Transform.n225 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17120 ),
            .carryout(\foc.u_Park_Transform.n17121 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_6_lut_LC_9_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_6_lut_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_6_lut_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_6_lut_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__32335),
            .in2(N__29218),
            .in3(N__29206),
            .lcout(\foc.u_Park_Transform.n274 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17121 ),
            .carryout(\foc.u_Park_Transform.n17122 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_7_lut_LC_9_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_7_lut_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_7_lut_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_7_lut_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__29203),
            .in2(N__32371),
            .in3(N__29194),
            .lcout(\foc.u_Park_Transform.n323 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17122 ),
            .carryout(\foc.u_Park_Transform.n17123 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_8_lut_LC_9_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_8_lut_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_8_lut_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_8_lut_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__32339),
            .in2(N__29191),
            .in3(N__29179),
            .lcout(\foc.u_Park_Transform.n372 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17123 ),
            .carryout(\foc.u_Park_Transform.n17124 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_9_lut_LC_9_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_9_lut_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_9_lut_LC_9_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_9_lut_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__29176),
            .in2(N__32372),
            .in3(N__29167),
            .lcout(\foc.u_Park_Transform.n421_adj_2039 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17124 ),
            .carryout(\foc.u_Park_Transform.n17125 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_10_lut_LC_9_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_10_lut_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_10_lut_LC_9_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_10_lut_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__32319),
            .in2(N__29323),
            .in3(N__29311),
            .lcout(\foc.u_Park_Transform.n470_adj_2038 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\foc.u_Park_Transform.n17126 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_11_lut_LC_9_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_11_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_11_lut_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_11_lut_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__29308),
            .in2(N__32367),
            .in3(N__29299),
            .lcout(\foc.u_Park_Transform.n519_adj_2035 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17126 ),
            .carryout(\foc.u_Park_Transform.n17127 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_12_lut_LC_9_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_12_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_12_lut_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_12_lut_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__32323),
            .in2(N__29290),
            .in3(N__29296),
            .lcout(\foc.u_Park_Transform.n568_adj_2034 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17127 ),
            .carryout(\foc.u_Park_Transform.n17128 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_13_lut_LC_9_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_13_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_13_lut_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_13_lut_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__29288),
            .in2(N__32368),
            .in3(N__29293),
            .lcout(\foc.u_Park_Transform.n617_adj_2031 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17128 ),
            .carryout(\foc.u_Park_Transform.n17129 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_14_lut_LC_9_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_14_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_14_lut_LC_9_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_570_14_lut_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__29289),
            .in2(N__30447),
            .in3(N__29269),
            .lcout(\foc.u_Park_Transform.n774_adj_2045 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17129 ),
            .carryout(\foc.u_Park_Transform.n775_adj_2047 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n775_adj_2047_THRU_LUT4_0_LC_9_12_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n775_adj_2047_THRU_LUT4_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n775_adj_2047_THRU_LUT4_0_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n775_adj_2047_THRU_LUT4_0_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29266),
            .lcout(\foc.u_Park_Transform.n775_adj_2047_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i22_2_lut_LC_9_14_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i22_2_lut_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i22_2_lut_LC_9_14_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i22_2_lut_LC_9_14_3  (
            .in0(N__32157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i528_2_lut_LC_9_14_4 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i528_2_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i528_2_lut_LC_9_14_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i528_2_lut_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32158),
            .lcout(\foc.u_Park_Transform.n777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_2_lut_LC_9_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_2_lut_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_2_lut_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_2_lut_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__30734),
            .in2(N__32384),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n78_adj_2145 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\foc.u_Park_Transform.n16935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_3_lut_LC_9_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_3_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_3_lut_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_3_lut_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__32363),
            .in2(N__30601),
            .in3(N__29350),
            .lcout(\foc.u_Park_Transform.n127_adj_2119 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16935 ),
            .carryout(\foc.u_Park_Transform.n16936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_4_lut_LC_9_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_4_lut_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_4_lut_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_4_lut_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__32381),
            .in2(N__30577),
            .in3(N__29347),
            .lcout(\foc.u_Park_Transform.n176_adj_2104 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16936 ),
            .carryout(\foc.u_Park_Transform.n16937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_5_lut_LC_9_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_5_lut_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_5_lut_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_5_lut_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__32364),
            .in2(N__30547),
            .in3(N__29344),
            .lcout(\foc.u_Park_Transform.n225_adj_2075 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16937 ),
            .carryout(\foc.u_Park_Transform.n16938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_6_lut_LC_9_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_6_lut_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_6_lut_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_6_lut_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__32382),
            .in2(N__30523),
            .in3(N__29341),
            .lcout(\foc.u_Park_Transform.n274_adj_2058 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16938 ),
            .carryout(\foc.u_Park_Transform.n16939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_7_lut_LC_9_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_7_lut_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_7_lut_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_7_lut_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__32365),
            .in2(N__30955),
            .in3(N__29338),
            .lcout(\foc.u_Park_Transform.n323_adj_2057 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16939 ),
            .carryout(\foc.u_Park_Transform.n16940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_8_lut_LC_9_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_8_lut_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_8_lut_LC_9_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_8_lut_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__32383),
            .in2(N__30928),
            .in3(N__29335),
            .lcout(\foc.u_Park_Transform.n372_adj_2042 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16940 ),
            .carryout(\foc.u_Park_Transform.n16941 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_9_lut_LC_9_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_9_lut_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_9_lut_LC_9_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_9_lut_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__32366),
            .in2(N__30901),
            .in3(N__29332),
            .lcout(\foc.u_Park_Transform.n421 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16941 ),
            .carryout(\foc.u_Park_Transform.n16942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_10_lut_LC_9_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_10_lut_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_10_lut_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_10_lut_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__30874),
            .in2(N__32385),
            .in3(N__29329),
            .lcout(\foc.u_Park_Transform.n470 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\foc.u_Park_Transform.n16943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_11_lut_LC_9_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_11_lut_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_11_lut_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_11_lut_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__32376),
            .in2(N__30865),
            .in3(N__29326),
            .lcout(\foc.u_Park_Transform.n519 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16943 ),
            .carryout(\foc.u_Park_Transform.n16944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_12_lut_LC_9_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_12_lut_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_12_lut_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_12_lut_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__30707),
            .in2(N__32386),
            .in3(N__29377),
            .lcout(\foc.u_Park_Transform.n568 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16944 ),
            .carryout(\foc.u_Park_Transform.n16945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_13_lut_LC_9_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_13_lut_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_13_lut_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_13_lut_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__32380),
            .in2(N__30712),
            .in3(N__29374),
            .lcout(\foc.u_Park_Transform.n617 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16945 ),
            .carryout(\foc.u_Park_Transform.n16946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_14_lut_LC_9_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_14_lut_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_570_14_lut_LC_9_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_570_14_lut_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__30711),
            .in2(N__30451),
            .in3(N__29371),
            .lcout(\foc.u_Park_Transform.n774 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16946 ),
            .carryout(\foc.u_Park_Transform.n775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n775_THRU_LUT4_0_LC_9_16_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n775_THRU_LUT4_0_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n775_THRU_LUT4_0_LC_9_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n775_THRU_LUT4_0_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29368),
            .lcout(\foc.u_Park_Transform.n775_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut_LC_9_19_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut_LC_9_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__44946),
            .in2(_gnd_net_),
            .in3(N__29365),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2807 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut_LC_9_19_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut_LC_9_19_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__44949),
            .in2(_gnd_net_),
            .in3(N__29362),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2810 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15460 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut_LC_9_19_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut_LC_9_19_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__68428),
            .in2(_gnd_net_),
            .in3(N__29359),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2813 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15461 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut_LC_9_19_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut_LC_9_19_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__44950),
            .in2(_gnd_net_),
            .in3(N__29356),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2816 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15462 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut_LC_9_19_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut_LC_9_19_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__44947),
            .in2(_gnd_net_),
            .in3(N__29353),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2819 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15463 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut_LC_9_19_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut_LC_9_19_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__44951),
            .in2(_gnd_net_),
            .in3(N__29623),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2822 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15464 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut_LC_9_19_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut_LC_9_19_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__44948),
            .in2(_gnd_net_),
            .in3(N__29620),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2825 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15465 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut_LC_9_19_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut_LC_9_19_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__44952),
            .in2(_gnd_net_),
            .in3(N__29617),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2828 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15466 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15467 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut_LC_9_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut_LC_9_20_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__44954),
            .in2(_gnd_net_),
            .in3(N__29614),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2831 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut_LC_9_20_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut_LC_9_20_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__44953),
            .in2(_gnd_net_),
            .in3(N__29563),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2834 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15468 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut_LC_9_20_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut_LC_9_20_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__44955),
            .in2(_gnd_net_),
            .in3(N__29449),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2840 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15469 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut_LC_9_20_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut_LC_9_20_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__68436),
            .in2(_gnd_net_),
            .in3(N__29383),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2843 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15470 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15471 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut_LC_9_20_4 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut_LC_9_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut_LC_9_20_4  (
            .in0(N__68437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29380),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_sub_temp1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_2_lut_LC_9_21_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_2_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_2_lut_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_2_lut_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__32693),
            .in2(N__29672),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2332 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_3_lut_LC_9_21_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_3_lut_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_3_lut_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_3_lut_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__29803),
            .in2(_gnd_net_),
            .in3(N__29791),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2432 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17431 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_4_lut_LC_9_21_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_4_lut_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_4_lut_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_4_lut_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__29788),
            .in2(N__29673),
            .in3(N__29776),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2532 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17432 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_5_lut_LC_9_21_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_5_lut_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_5_lut_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_5_lut_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__29658),
            .in2(N__29773),
            .in3(N__29758),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2632 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17433 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_6_lut_LC_9_21_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_6_lut_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_6_lut_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_6_lut_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__29755),
            .in2(N__29674),
            .in3(N__29743),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2732 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17434 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_7_lut_LC_9_21_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_7_lut_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_7_lut_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_7_lut_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__29662),
            .in2(N__29740),
            .in3(N__29725),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2832 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17435 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_8_lut_LC_9_21_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_8_lut_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_8_lut_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_8_lut_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__29722),
            .in2(N__29675),
            .in3(N__29710),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2932 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17436 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_9_lut_LC_9_21_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_9_lut_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_9_lut_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_9_lut_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__29707),
            .in2(N__29676),
            .in3(N__29695),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3032 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17437 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17438 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_10_lut_LC_9_22_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_10_lut_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_10_lut_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_10_lut_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__29692),
            .in2(N__29680),
            .in3(N__29626),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3132 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_11_lut_LC_9_22_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_11_lut_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_11_lut_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2271_11_lut_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__29920),
            .in2(_gnd_net_),
            .in3(N__29908),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3243 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17439 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_LUT4_0_LC_9_22_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_LUT4_0_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_LUT4_0_LC_9_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_LUT4_0_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29905),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3244_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_2_lut_LC_9_23_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_2_lut_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_2_lut_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_2_lut_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__31500),
            .in2(N__32770),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7473 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_3_lut_LC_9_23_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_3_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_3_lut_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_3_lut_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__29902),
            .in2(_gnd_net_),
            .in3(N__29890),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7553 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17337 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_4_lut_LC_9_23_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_4_lut_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_4_lut_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_4_lut_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__31501),
            .in2(N__29887),
            .in3(N__29872),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7552 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17338 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_5_lut_LC_9_23_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_5_lut_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_5_lut_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_5_lut_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__29869),
            .in2(N__31518),
            .in3(N__29857),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7551 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17339 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_6_lut_LC_9_23_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_6_lut_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_6_lut_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_6_lut_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__31505),
            .in2(N__29854),
            .in3(N__29839),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7550 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17340 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_7_lut_LC_9_23_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_7_lut_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_7_lut_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_7_lut_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__29836),
            .in2(N__31519),
            .in3(N__29824),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7549 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17341 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_8_lut_LC_9_23_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_8_lut_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_8_lut_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_8_lut_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__31509),
            .in2(N__29821),
            .in3(N__29806),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7548 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17342 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17343 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_9_lut_LC_9_23_7 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_9_lut_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_9_lut_LC_9_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5953_9_lut_LC_9_23_7  (
            .in0(N__31510),
            .in1(N__30049),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_2_lut_LC_9_24_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_2_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_2_lut_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_2_lut_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__32798),
            .in2(N__31496),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2347 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_3_lut_LC_9_24_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_3_lut_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_3_lut_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_3_lut_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__30022),
            .in2(_gnd_net_),
            .in3(N__30001),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2447 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17481 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_4_lut_LC_9_24_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_4_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_4_lut_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_4_lut_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__31243),
            .in2(N__31497),
            .in3(N__29986),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2547 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17482 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_5_lut_LC_9_24_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_5_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_5_lut_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_5_lut_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__31464),
            .in2(N__31222),
            .in3(N__29968),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2647 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17483 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_6_lut_LC_9_24_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_6_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_6_lut_LC_9_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_6_lut_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__31669),
            .in2(N__31498),
            .in3(N__29953),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2747 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17484 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_7_lut_LC_9_24_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_7_lut_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_7_lut_LC_9_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_7_lut_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__31468),
            .in2(N__31651),
            .in3(N__29938),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2847 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17485 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_8_lut_LC_9_24_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_8_lut_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_8_lut_LC_9_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_8_lut_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__31630),
            .in2(N__31499),
            .in3(N__29923),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2947 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17486 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_9_lut_LC_9_24_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_9_lut_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_9_lut_LC_9_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_9_lut_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__31472),
            .in2(N__31612),
            .in3(N__30085),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3047 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17487 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17488 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_10_lut_LC_9_25_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_10_lut_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_10_lut_LC_9_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_10_lut_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__31591),
            .in2(N__31495),
            .in3(N__30070),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3147 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17489 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_11_lut_LC_9_25_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_11_lut_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_11_lut_LC_9_25_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2276_11_lut_LC_9_25_1  (
            .in0(N__31381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30067),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_2_lut_LC_10_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_2_lut_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_2_lut_LC_10_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_2_lut_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__34278),
            .in2(N__35893),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n72 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\foc.u_Park_Transform.n17146 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_3_lut_LC_10_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_3_lut_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_3_lut_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_3_lut_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__35870),
            .in2(N__30262),
            .in3(N__30064),
            .lcout(\foc.u_Park_Transform.n121 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17146 ),
            .carryout(\foc.u_Park_Transform.n17147 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_4_lut_LC_10_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_4_lut_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_4_lut_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_4_lut_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__35871),
            .in2(N__30241),
            .in3(N__30061),
            .lcout(\foc.u_Park_Transform.n170 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17147 ),
            .carryout(\foc.u_Park_Transform.n17148 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_5_lut_LC_10_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_5_lut_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_5_lut_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_5_lut_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__30217),
            .in2(N__35894),
            .in3(N__30058),
            .lcout(\foc.u_Park_Transform.n219 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17148 ),
            .carryout(\foc.u_Park_Transform.n17149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_6_lut_LC_10_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_6_lut_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_6_lut_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_6_lut_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__35875),
            .in2(N__30199),
            .in3(N__30055),
            .lcout(\foc.u_Park_Transform.n268 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17149 ),
            .carryout(\foc.u_Park_Transform.n17150 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_7_lut_LC_10_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_7_lut_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_7_lut_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_7_lut_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__30175),
            .in2(N__35895),
            .in3(N__30052),
            .lcout(\foc.u_Park_Transform.n317 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17150 ),
            .carryout(\foc.u_Park_Transform.n17151 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_8_lut_LC_10_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_8_lut_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_8_lut_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_8_lut_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__35879),
            .in2(N__30157),
            .in3(N__30121),
            .lcout(\foc.u_Park_Transform.n366 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17151 ),
            .carryout(\foc.u_Park_Transform.n17152 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_9_lut_LC_10_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_9_lut_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_9_lut_LC_10_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_9_lut_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__30133),
            .in2(N__35896),
            .in3(N__30118),
            .lcout(\foc.u_Park_Transform.n415_adj_2008 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17152 ),
            .carryout(\foc.u_Park_Transform.n17153 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_10_lut_LC_10_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_10_lut_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_10_lut_LC_10_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_10_lut_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__30412),
            .in2(N__35810),
            .in3(N__30115),
            .lcout(\foc.u_Park_Transform.n464_adj_2005 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\foc.u_Park_Transform.n17154 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_11_lut_LC_10_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_11_lut_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_11_lut_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_11_lut_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__35758),
            .in2(N__30397),
            .in3(N__30112),
            .lcout(\foc.u_Park_Transform.n513_adj_2002 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17154 ),
            .carryout(\foc.u_Park_Transform.n17155 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_12_lut_LC_10_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_12_lut_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_12_lut_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_12_lut_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__30373),
            .in2(N__35811),
            .in3(N__30109),
            .lcout(\foc.u_Park_Transform.n562_adj_2000 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17155 ),
            .carryout(\foc.u_Park_Transform.n17156 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_13_lut_LC_10_10_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_13_lut_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_13_lut_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_13_lut_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__35762),
            .in2(N__30355),
            .in3(N__30106),
            .lcout(\foc.u_Park_Transform.n611 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17156 ),
            .carryout(\foc.u_Park_Transform.n17157 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_14_lut_LC_10_10_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_14_lut_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_14_lut_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_14_lut_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__30331),
            .in2(N__35812),
            .in3(N__30103),
            .lcout(\foc.u_Park_Transform.n660 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17157 ),
            .carryout(\foc.u_Park_Transform.n17158 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_15_lut_LC_10_10_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_15_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_15_lut_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_15_lut_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__35766),
            .in2(N__30319),
            .in3(N__30100),
            .lcout(\foc.u_Park_Transform.n709 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17158 ),
            .carryout(\foc.u_Park_Transform.n17159 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_16_lut_LC_10_10_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_16_lut_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_16_lut_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_568_16_lut_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__34500),
            .in2(N__30304),
            .in3(N__30097),
            .lcout(\foc.u_Park_Transform.n766 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17159 ),
            .carryout(\foc.u_Park_Transform.n767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n767_THRU_LUT4_0_LC_10_10_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n767_THRU_LUT4_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n767_THRU_LUT4_0_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n767_THRU_LUT4_0_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30265),
            .lcout(\foc.u_Park_Transform.n767_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_2_lut_LC_10_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_2_lut_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_2_lut_LC_10_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_2_lut_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__32318),
            .in2(N__34272),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n75 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\foc.u_Park_Transform.n17131 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_3_lut_LC_10_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_3_lut_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_3_lut_LC_10_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_3_lut_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__34227),
            .in2(N__30250),
            .in3(N__30229),
            .lcout(\foc.u_Park_Transform.n124 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17131 ),
            .carryout(\foc.u_Park_Transform.n17132 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_4_lut_LC_10_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_4_lut_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_4_lut_LC_10_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_4_lut_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__34228),
            .in2(N__30226),
            .in3(N__30208),
            .lcout(\foc.u_Park_Transform.n173 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17132 ),
            .carryout(\foc.u_Park_Transform.n17133 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_5_lut_LC_10_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_5_lut_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_5_lut_LC_10_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_5_lut_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__30205),
            .in2(N__34273),
            .in3(N__30187),
            .lcout(\foc.u_Park_Transform.n222 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17133 ),
            .carryout(\foc.u_Park_Transform.n17134 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_6_lut_LC_10_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_6_lut_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_6_lut_LC_10_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_6_lut_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__34232),
            .in2(N__30184),
            .in3(N__30166),
            .lcout(\foc.u_Park_Transform.n271 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17134 ),
            .carryout(\foc.u_Park_Transform.n17135 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_7_lut_LC_10_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_7_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_7_lut_LC_10_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_7_lut_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__30163),
            .in2(N__34274),
            .in3(N__30145),
            .lcout(\foc.u_Park_Transform.n320 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17135 ),
            .carryout(\foc.u_Park_Transform.n17136 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_8_lut_LC_10_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_8_lut_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_8_lut_LC_10_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_8_lut_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__34236),
            .in2(N__30142),
            .in3(N__30124),
            .lcout(\foc.u_Park_Transform.n369 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17136 ),
            .carryout(\foc.u_Park_Transform.n17137 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_9_lut_LC_10_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_9_lut_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_9_lut_LC_10_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_9_lut_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__30418),
            .in2(N__34275),
            .in3(N__30406),
            .lcout(\foc.u_Park_Transform.n418_adj_2024 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17137 ),
            .carryout(\foc.u_Park_Transform.n17138 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_10_lut_LC_10_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_10_lut_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_10_lut_LC_10_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_10_lut_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__30403),
            .in2(N__34221),
            .in3(N__30385),
            .lcout(\foc.u_Park_Transform.n467_adj_2019 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\foc.u_Park_Transform.n17139 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_11_lut_LC_10_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_11_lut_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_11_lut_LC_10_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_11_lut_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__34165),
            .in2(N__30382),
            .in3(N__30364),
            .lcout(\foc.u_Park_Transform.n516_adj_2018 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17139 ),
            .carryout(\foc.u_Park_Transform.n17140 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_12_lut_LC_10_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_12_lut_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_12_lut_LC_10_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_12_lut_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__30361),
            .in2(N__34222),
            .in3(N__30343),
            .lcout(\foc.u_Park_Transform.n565 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17140 ),
            .carryout(\foc.u_Park_Transform.n17141 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_13_lut_LC_10_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_13_lut_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_13_lut_LC_10_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_13_lut_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__34169),
            .in2(N__30340),
            .in3(N__30322),
            .lcout(\foc.u_Park_Transform.n614_adj_2017 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17141 ),
            .carryout(\foc.u_Park_Transform.n17142 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_14_lut_LC_10_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_14_lut_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_14_lut_LC_10_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_14_lut_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__30281),
            .in2(N__34223),
            .in3(N__30307),
            .lcout(\foc.u_Park_Transform.n663_adj_2016 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17142 ),
            .carryout(\foc.u_Park_Transform.n17143 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_15_lut_LC_10_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_15_lut_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_15_lut_LC_10_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_15_lut_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__34173),
            .in2(N__30288),
            .in3(N__30292),
            .lcout(\foc.u_Park_Transform.n712_adj_2015 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17143 ),
            .carryout(\foc.u_Park_Transform.n17144 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_16_lut_LC_10_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_16_lut_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_16_lut_LC_10_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_569_16_lut_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__32619),
            .in2(N__30289),
            .in3(N__30268),
            .lcout(\foc.u_Park_Transform.n770_adj_2030 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17144 ),
            .carryout(\foc.u_Park_Transform.n771_adj_2032 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n771_adj_2032_THRU_LUT4_0_LC_10_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n771_adj_2032_THRU_LUT4_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n771_adj_2032_THRU_LUT4_0_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n771_adj_2032_THRU_LUT4_0_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30454),
            .lcout(\foc.u_Park_Transform.n771_adj_2032_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i20_2_lut_LC_10_13_0 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i20_2_lut_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i20_2_lut_LC_10_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i20_2_lut_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32169),
            .lcout(\foc.u_Park_Transform.n616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i18_2_lut_LC_10_13_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i18_2_lut_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i18_2_lut_LC_10_13_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i18_2_lut_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32181),
            .lcout(\foc.u_Park_Transform.n613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i525_2_lut_LC_10_13_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i525_2_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i525_2_lut_LC_10_13_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i525_2_lut_LC_10_13_3  (
            .in0(N__32170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i522_2_lut_LC_10_13_6 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i522_2_lut_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i522_2_lut_LC_10_13_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i522_2_lut_LC_10_13_6  (
            .in0(N__32182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_2_lut_LC_10_14_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_2_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_2_lut_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_2_lut_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__44241),
            .in2(N__32134),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n87 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\foc.u_Park_Transform.n18160 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_3_lut_LC_10_14_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_3_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_3_lut_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_3_lut_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__32124),
            .in2(N__32029),
            .in3(N__30430),
            .lcout(\foc.u_Park_Transform.n136 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18160 ),
            .carryout(\foc.u_Park_Transform.n18161 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_4_lut_LC_10_14_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_4_lut_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_4_lut_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_4_lut_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__32135),
            .in2(N__32047),
            .in3(N__30427),
            .lcout(\foc.u_Park_Transform.n185 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18161 ),
            .carryout(\foc.u_Park_Transform.n18162 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_5_lut_LC_10_14_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_5_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_5_lut_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_5_lut_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__32125),
            .in2(N__34317),
            .in3(N__30424),
            .lcout(\foc.u_Park_Transform.n234 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18162 ),
            .carryout(\foc.u_Park_Transform.n18163 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_6_lut_LC_10_14_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_6_lut_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_6_lut_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_6_lut_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__32136),
            .in2(N__34360),
            .in3(N__30421),
            .lcout(\foc.u_Park_Transform.n283 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18163 ),
            .carryout(\foc.u_Park_Transform.n18164 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_7_lut_LC_10_14_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_7_lut_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_7_lut_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_7_lut_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__34349),
            .in2(N__32140),
            .in3(N__30508),
            .lcout(\foc.u_Park_Transform.n332 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18164 ),
            .carryout(\foc.u_Park_Transform.n18165 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_8_lut_LC_10_14_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_8_lut_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_573_8_lut_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_573_8_lut_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__32397),
            .in2(N__34361),
            .in3(N__30505),
            .lcout(\foc.u_Park_Transform.n786 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n18165 ),
            .carryout(\foc.u_Park_Transform.n787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n787_THRU_LUT4_0_LC_10_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n787_THRU_LUT4_0_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n787_THRU_LUT4_0_LC_10_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n787_THRU_LUT4_0_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30502),
            .lcout(\foc.u_Park_Transform.n787_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_2_lut_LC_10_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_2_lut_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_2_lut_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_2_lut_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__32133),
            .in2(N__31788),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n84_adj_2118 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\foc.u_Park_Transform.n16915 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_3_lut_LC_10_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_3_lut_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_3_lut_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_3_lut_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__31772),
            .in2(N__30499),
            .in3(N__30490),
            .lcout(\foc.u_Park_Transform.n133 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16915 ),
            .carryout(\foc.u_Park_Transform.n16916 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_4_lut_LC_10_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_4_lut_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_4_lut_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_4_lut_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__31773),
            .in2(N__30487),
            .in3(N__30478),
            .lcout(\foc.u_Park_Transform.n182 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16916 ),
            .carryout(\foc.u_Park_Transform.n16917 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_5_lut_LC_10_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_5_lut_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_5_lut_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_5_lut_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__30475),
            .in2(N__31789),
            .in3(N__30469),
            .lcout(\foc.u_Park_Transform.n231 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16917 ),
            .carryout(\foc.u_Park_Transform.n16918 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_6_lut_LC_10_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_6_lut_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_6_lut_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_6_lut_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__31777),
            .in2(N__30466),
            .in3(N__30457),
            .lcout(\foc.u_Park_Transform.n280 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16918 ),
            .carryout(\foc.u_Park_Transform.n16919 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_7_lut_LC_10_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_7_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_7_lut_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_7_lut_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__30646),
            .in2(N__31790),
            .in3(N__30640),
            .lcout(\foc.u_Park_Transform.n329 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16919 ),
            .carryout(\foc.u_Park_Transform.n16920 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_8_lut_LC_10_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_8_lut_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_8_lut_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_8_lut_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__31781),
            .in2(N__30627),
            .in3(N__30637),
            .lcout(\foc.u_Park_Transform.n378 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16920 ),
            .carryout(\foc.u_Park_Transform.n16921 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_9_lut_LC_10_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_9_lut_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_9_lut_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_9_lut_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__30623),
            .in2(N__31791),
            .in3(N__30634),
            .lcout(\foc.u_Park_Transform.n427 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16921 ),
            .carryout(\foc.u_Park_Transform.n16922 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_10_lut_LC_10_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_10_lut_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_572_10_lut_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_572_10_lut_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__32011),
            .in2(N__30631),
            .in3(N__30607),
            .lcout(\foc.u_Park_Transform.n782 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\foc.u_Park_Transform.n783_adj_2167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n783_adj_2167_THRU_LUT4_0_LC_10_16_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n783_adj_2167_THRU_LUT4_0_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n783_adj_2167_THRU_LUT4_0_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n783_adj_2167_THRU_LUT4_0_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30604),
            .lcout(\foc.u_Park_Transform.n783_adj_2167_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_2_lut_LC_10_17_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_2_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_2_lut_LC_10_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_2_lut_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__31792),
            .in2(N__30845),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n81_adj_2120 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\foc.u_Park_Transform.n16924 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_3_lut_LC_10_17_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_3_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_3_lut_LC_10_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_3_lut_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__30820),
            .in2(N__30589),
            .in3(N__30562),
            .lcout(\foc.u_Park_Transform.n130_adj_2105 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16924 ),
            .carryout(\foc.u_Park_Transform.n16925 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_4_lut_LC_10_17_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_4_lut_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_4_lut_LC_10_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_4_lut_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__30821),
            .in2(N__30559),
            .in3(N__30535),
            .lcout(\foc.u_Park_Transform.n179_adj_2076 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16925 ),
            .carryout(\foc.u_Park_Transform.n16926 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_5_lut_LC_10_17_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_5_lut_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_5_lut_LC_10_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_5_lut_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__30532),
            .in2(N__30846),
            .in3(N__30511),
            .lcout(\foc.u_Park_Transform.n228 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16926 ),
            .carryout(\foc.u_Park_Transform.n16927 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_6_lut_LC_10_17_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_6_lut_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_6_lut_LC_10_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_6_lut_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__30825),
            .in2(N__30967),
            .in3(N__30940),
            .lcout(\foc.u_Park_Transform.n277 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16927 ),
            .carryout(\foc.u_Park_Transform.n16928 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_7_lut_LC_10_17_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_7_lut_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_7_lut_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_7_lut_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__30937),
            .in2(N__30847),
            .in3(N__30916),
            .lcout(\foc.u_Park_Transform.n326 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16928 ),
            .carryout(\foc.u_Park_Transform.n16929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_8_lut_LC_10_17_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_8_lut_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_8_lut_LC_10_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_8_lut_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__30829),
            .in2(N__30913),
            .in3(N__30886),
            .lcout(\foc.u_Park_Transform.n375 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16929 ),
            .carryout(\foc.u_Park_Transform.n16930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_9_lut_LC_10_17_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_9_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_9_lut_LC_10_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_9_lut_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__30883),
            .in2(N__30848),
            .in3(N__30868),
            .lcout(\foc.u_Park_Transform.n424 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16930 ),
            .carryout(\foc.u_Park_Transform.n16931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_10_lut_LC_10_18_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_10_lut_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_10_lut_LC_10_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_10_lut_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__30833),
            .in2(N__30672),
            .in3(N__30853),
            .lcout(\foc.u_Park_Transform.n473 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\foc.u_Park_Transform.n16932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_11_lut_LC_10_18_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_11_lut_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_11_lut_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_11_lut_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__30668),
            .in2(N__30849),
            .in3(N__30694),
            .lcout(\foc.u_Park_Transform.n522 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16932 ),
            .carryout(\foc.u_Park_Transform.n16933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_12_lut_LC_10_18_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_12_lut_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_571_12_lut_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_571_12_lut_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__30691),
            .in2(N__30673),
            .in3(N__30652),
            .lcout(\foc.u_Park_Transform.n778 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16933 ),
            .carryout(\foc.u_Park_Transform.n779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n779_THRU_LUT4_0_LC_10_18_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n779_THRU_LUT4_0_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n779_THRU_LUT4_0_LC_10_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n779_THRU_LUT4_0_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30649),
            .lcout(\foc.u_Park_Transform.n779_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_2_lut_LC_10_19_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_2_lut_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_2_lut_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_2_lut_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__31287),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2417 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_3_lut_LC_10_19_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_3_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_3_lut_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_3_lut_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__34779),
            .in2(N__31129),
            .in3(N__30991),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2517 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17385 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_4_lut_LC_10_19_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_4_lut_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_4_lut_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_4_lut_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__31114),
            .in2(N__34795),
            .in3(N__30988),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2617 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17386 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_5_lut_LC_10_19_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_5_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_5_lut_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_5_lut_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__34783),
            .in2(N__31099),
            .in3(N__30985),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2717 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17387 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_6_lut_LC_10_19_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_6_lut_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_6_lut_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_6_lut_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__31081),
            .in2(N__34796),
            .in3(N__30982),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2817 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17388 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_7_lut_LC_10_19_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_7_lut_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_7_lut_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_7_lut_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__34787),
            .in2(N__31069),
            .in3(N__30979),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2917 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17389 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_8_lut_LC_10_19_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_8_lut_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_8_lut_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_8_lut_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__31348),
            .in2(N__34797),
            .in3(N__30976),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3017 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17390 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_9_lut_LC_10_19_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_9_lut_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_9_lut_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_9_lut_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__34791),
            .in2(N__31336),
            .in3(N__30973),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3117 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17391 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17392 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_10_lut_LC_10_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_10_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_10_lut_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5958_10_lut_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__31276),
            .in2(_gnd_net_),
            .in3(N__30970),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3223 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_LUT4_0_LC_10_20_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_LUT4_0_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_LUT4_0_LC_10_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_LUT4_0_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31054),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3224_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_2_lut_LC_10_21_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_2_lut_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_2_lut_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_2_lut_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__31173),
            .in2(N__32738),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2329 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_3_lut_LC_10_21_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_3_lut_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_3_lut_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_3_lut_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__31051),
            .in2(_gnd_net_),
            .in3(N__31045),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2429 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17421 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_4_lut_LC_10_21_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_4_lut_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_4_lut_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_4_lut_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__31174),
            .in2(N__31042),
            .in3(N__31033),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2529 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17422 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_5_lut_LC_10_21_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_5_lut_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_5_lut_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_5_lut_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__31030),
            .in2(N__31191),
            .in3(N__31024),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2629 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17423 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_6_lut_LC_10_21_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_6_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_6_lut_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_6_lut_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__31178),
            .in2(N__31021),
            .in3(N__31012),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2729 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17424 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_7_lut_LC_10_21_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_7_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_7_lut_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_7_lut_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__31009),
            .in2(N__31192),
            .in3(N__31003),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2829 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17425 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_8_lut_LC_10_21_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_8_lut_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_8_lut_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_8_lut_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__31000),
            .in2(N__31194),
            .in3(N__30994),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2929 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17426 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_9_lut_LC_10_21_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_9_lut_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_9_lut_LC_10_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_9_lut_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__31210),
            .in2(N__31193),
            .in3(N__31204),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3029 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17427 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17428 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_10_lut_LC_10_22_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_10_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_10_lut_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_10_lut_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__31201),
            .in2(N__31195),
            .in3(N__31144),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3129 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_11_lut_LC_10_22_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_11_lut_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_11_lut_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_add_2270_11_lut_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__31141),
            .in2(_gnd_net_),
            .in3(N__31135),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3239 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17429 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_LUT4_0_LC_10_22_2 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_LUT4_0_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_LUT4_0_LC_10_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_LUT4_0_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31132),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3240_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_2_lut_LC_10_23_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_2_lut_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_2_lut_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_2_lut_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__33495),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2420 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_3_lut_LC_10_23_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_3_lut_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_3_lut_LC_10_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_3_lut_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__31306),
            .in2(N__33295),
            .in3(N__31102),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2520 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17394 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_4_lut_LC_10_23_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_4_lut_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_4_lut_LC_10_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_4_lut_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__33640),
            .in2(N__31319),
            .in3(N__31084),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2620 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17395 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_5_lut_LC_10_23_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_5_lut_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_5_lut_LC_10_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_5_lut_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__31310),
            .in2(N__33622),
            .in3(N__31072),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2720 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17396 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_6_lut_LC_10_23_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_6_lut_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_6_lut_LC_10_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_6_lut_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__33598),
            .in2(N__31320),
            .in3(N__31057),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2820 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17397 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_7_lut_LC_10_23_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_7_lut_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_7_lut_LC_10_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_7_lut_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__31314),
            .in2(N__33580),
            .in3(N__31339),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2920 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17398 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_8_lut_LC_10_23_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_8_lut_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_8_lut_LC_10_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_8_lut_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__33556),
            .in2(N__31321),
            .in3(N__31324),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3020 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17399 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_9_lut_LC_10_23_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_9_lut_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_9_lut_LC_10_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_9_lut_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__31318),
            .in2(N__33538),
            .in3(N__31267),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3120 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17400 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17401 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_10_lut_LC_10_24_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_10_lut_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_10_lut_LC_10_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5959_10_lut_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__33457),
            .in2(_gnd_net_),
            .in3(N__31264),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3227 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_LUT4_0_LC_10_24_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_LUT4_0_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_LUT4_0_LC_10_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_LUT4_0_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31261),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3228_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_i1719_2_lut_LC_10_25_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_i1719_2_lut_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_i1719_2_lut_LC_10_25_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_f1_31__I_0_i1719_2_lut_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__31439),
            .in2(N__32805),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2652 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_3_lut_LC_10_25_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_3_lut_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_3_lut_LC_10_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_3_lut_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__31258),
            .in2(_gnd_net_),
            .in3(N__31237),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7472 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17350 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_4_lut_LC_10_25_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_4_lut_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_4_lut_LC_10_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_4_lut_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(N__31440),
            .in2(N__31234),
            .in3(N__31213),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7471 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17351 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_5_lut_LC_10_25_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_5_lut_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_5_lut_LC_10_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_5_lut_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__31447),
            .in2(N__31681),
            .in3(N__31663),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7470 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17352 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_6_lut_LC_10_25_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_6_lut_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_6_lut_LC_10_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_6_lut_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__31660),
            .in2(N__31493),
            .in3(N__31642),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7469 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17353 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_7_lut_LC_10_25_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_7_lut_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_7_lut_LC_10_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_7_lut_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(N__31639),
            .in2(N__31491),
            .in3(N__31624),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7468 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17354 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_8_lut_LC_10_25_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_8_lut_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_8_lut_LC_10_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_8_lut_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(N__31621),
            .in2(N__31494),
            .in3(N__31603),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7467 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17355 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_9_lut_LC_10_25_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_9_lut_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_9_lut_LC_10_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_9_lut_LC_10_25_7  (
            .in0(_gnd_net_),
            .in1(N__31600),
            .in2(N__31492),
            .in3(N__31585),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7466 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17356 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17357 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_10_lut_LC_10_26_0 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_10_lut_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_10_lut_LC_10_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5928_10_lut_LC_10_26_0  (
            .in0(N__31582),
            .in1(N__31457),
            .in2(_gnd_net_),
            .in3(N__31384),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n7465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_2_lut_LC_11_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_2_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_2_lut_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_2_lut_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__32117),
            .in2(N__31733),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n84 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\foc.u_Park_Transform.n17098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_3_lut_LC_11_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_3_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_3_lut_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_3_lut_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__31714),
            .in2(N__31993),
            .in3(N__31351),
            .lcout(\foc.u_Park_Transform.n133_adj_2101 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17098 ),
            .carryout(\foc.u_Park_Transform.n17099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_4_lut_LC_11_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_4_lut_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_4_lut_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__31715),
            .in2(N__31981),
            .in3(N__31888),
            .lcout(\foc.u_Park_Transform.n182_adj_2094 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17099 ),
            .carryout(\foc.u_Park_Transform.n17100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_5_lut_LC_11_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_5_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_5_lut_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_5_lut_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__31966),
            .in2(N__31734),
            .in3(N__31873),
            .lcout(\foc.u_Park_Transform.n231_adj_2089 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17100 ),
            .carryout(\foc.u_Park_Transform.n17101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_6_lut_LC_11_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_6_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_6_lut_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_6_lut_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__31719),
            .in2(N__31954),
            .in3(N__31858),
            .lcout(\foc.u_Park_Transform.n280_adj_2087 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17101 ),
            .carryout(\foc.u_Park_Transform.n17102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_7_lut_LC_11_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_7_lut_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_7_lut_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_7_lut_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__31939),
            .in2(N__31735),
            .in3(N__31840),
            .lcout(\foc.u_Park_Transform.n329_adj_2080 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17102 ),
            .carryout(\foc.u_Park_Transform.n17103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_8_lut_LC_11_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_8_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_8_lut_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_8_lut_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__31723),
            .in2(N__31927),
            .in3(N__31828),
            .lcout(\foc.u_Park_Transform.n378_adj_2078 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17103 ),
            .carryout(\foc.u_Park_Transform.n17104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_9_lut_LC_11_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_9_lut_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_9_lut_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_9_lut_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__31926),
            .in2(N__31736),
            .in3(N__31801),
            .lcout(\foc.u_Park_Transform.n427_adj_2069 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17104 ),
            .carryout(\foc.u_Park_Transform.n17105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_10_lut_LC_11_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_10_lut_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_10_lut_LC_11_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_572_10_lut_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__32004),
            .in2(N__31922),
            .in3(N__31798),
            .lcout(\foc.u_Park_Transform.n782_adj_2109 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\foc.u_Park_Transform.n783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n783_THRU_LUT4_0_LC_11_10_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n783_THRU_LUT4_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n783_THRU_LUT4_0_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n783_THRU_LUT4_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31795),
            .lcout(\foc.u_Park_Transform.n783_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i24_2_lut_LC_11_10_2 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i24_2_lut_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i24_2_lut_LC_11_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i24_2_lut_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32445),
            .lcout(\foc.u_Park_Transform.n622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i531_2_lut_LC_11_10_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i531_2_lut_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i531_2_lut_LC_11_10_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i531_2_lut_LC_11_10_5  (
            .in0(N__32446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_2_lut_LC_11_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_2_lut_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_2_lut_LC_11_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_2_lut_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__44254),
            .in2(N__32113),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n87_adj_2138 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\foc.u_Park_Transform.n17980 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_3_lut_LC_11_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_3_lut_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_3_lut_LC_11_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_3_lut_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__32022),
            .in2(N__32115),
            .in3(N__31969),
            .lcout(\foc.u_Park_Transform.n136_adj_2127 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17980 ),
            .carryout(\foc.u_Park_Transform.n17981 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_4_lut_LC_11_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_4_lut_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_4_lut_LC_11_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_4_lut_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__32040),
            .in2(N__32114),
            .in3(N__31957),
            .lcout(\foc.u_Park_Transform.n185_adj_2126 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17981 ),
            .carryout(\foc.u_Park_Transform.n17982 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_5_lut_LC_11_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_5_lut_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_5_lut_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_5_lut_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__32089),
            .in2(N__34321),
            .in3(N__31942),
            .lcout(\foc.u_Park_Transform.n234_adj_2125 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17982 ),
            .carryout(\foc.u_Park_Transform.n17983 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_6_lut_LC_11_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_6_lut_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_6_lut_LC_11_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_6_lut_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__32093),
            .in2(N__34362),
            .in3(N__31930),
            .lcout(\foc.u_Park_Transform.n283_adj_2122 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17983 ),
            .carryout(\foc.u_Park_Transform.n17984 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_7_lut_LC_11_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_7_lut_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_7_lut_LC_11_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_7_lut_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__34356),
            .in2(N__32116),
            .in3(N__31903),
            .lcout(\foc.u_Park_Transform.n332_adj_2110 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17984 ),
            .carryout(\foc.u_Park_Transform.n17985 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_8_lut_LC_11_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_8_lut_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_8_lut_LC_11_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_573_8_lut_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__32404),
            .in2(N__34363),
            .in3(N__31900),
            .lcout(\foc.u_Park_Transform.n786_adj_2152 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17985 ),
            .carryout(\foc.u_Park_Transform.n787_adj_2149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n787_adj_2149_THRU_LUT4_0_LC_11_11_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n787_adj_2149_THRU_LUT4_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n787_adj_2149_THRU_LUT4_0_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n787_adj_2149_THRU_LUT4_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32143),
            .lcout(\foc.u_Park_Transform.n787_adj_2149_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i519_2_lut_LC_11_12_0 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i519_2_lut_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i519_2_lut_LC_11_12_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i519_2_lut_LC_11_12_0  (
            .in0(N__32194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i26_2_lut_LC_11_12_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i26_2_lut_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i26_2_lut_LC_11_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i26_2_lut_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32419),
            .lcout(\foc.u_Park_Transform.n625 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16567_2_lut_LC_11_12_2.C_ON=1'b0;
    defparam i16567_2_lut_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam i16567_2_lut_LC_11_12_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i16567_2_lut_LC_11_12_2 (
            .in0(N__40485),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44410),
            .lcout(),
            .ltout(n21486_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_11_12_3.C_ON=1'b0;
    defparam i7_4_lut_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_11_12_3.LUT_INIT=16'b0101100101101010;
    LogicCell40 i7_4_lut_LC_11_12_3 (
            .in0(N__44253),
            .in1(_gnd_net_),
            .in2(N__32050),
            .in3(N__40446),
            .lcout(n139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i14_2_lut_LC_11_12_4 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i14_2_lut_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i14_2_lut_LC_11_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i14_2_lut_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32205),
            .lcout(\foc.u_Park_Transform.n607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i516_2_lut_LC_11_12_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i516_2_lut_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i516_2_lut_LC_11_12_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i516_2_lut_LC_11_12_5  (
            .in0(N__32206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i11560_3_lut_LC_11_12_6 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i11560_3_lut_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i11560_3_lut_LC_11_12_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \foc.u_Park_Transform.i11560_3_lut_LC_11_12_6  (
            .in0(N__40484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44409),
            .lcout(\foc.u_Park_Transform.n90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i16_2_lut_LC_11_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i16_2_lut_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i16_2_lut_LC_11_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i16_2_lut_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32193),
            .lcout(\foc.u_Park_Transform.n610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_2_lut_LC_11_13_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_2_lut_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_2_lut_LC_11_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_2_lut_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__32641),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.Look_Up_Table_out1_1_2 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_3_lut_LC_11_13_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_3_lut_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_3_lut_LC_11_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_3_lut_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__33043),
            .in2(_gnd_net_),
            .in3(N__32215),
            .lcout(\foc.Look_Up_Table_out1_1_3 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15944 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_4_lut_LC_11_13_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_4_lut_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_4_lut_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_4_lut_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__33031),
            .in2(_gnd_net_),
            .in3(N__32212),
            .lcout(\foc.Look_Up_Table_out1_1_4 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15945 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_5_lut_LC_11_13_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_5_lut_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_5_lut_LC_11_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_5_lut_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__33013),
            .in2(_gnd_net_),
            .in3(N__32209),
            .lcout(\foc.Look_Up_Table_out1_1_5 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15946 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_6_lut_LC_11_13_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_6_lut_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_6_lut_LC_11_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_6_lut_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__32980),
            .in2(_gnd_net_),
            .in3(N__32197),
            .lcout(\foc.Look_Up_Table_out1_1_6 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15947 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_7_lut_LC_11_13_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_7_lut_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_7_lut_LC_11_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_7_lut_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__32950),
            .in2(_gnd_net_),
            .in3(N__32185),
            .lcout(\foc.Look_Up_Table_out1_1_7 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15948 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_8_lut_LC_11_13_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_8_lut_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_8_lut_LC_11_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_8_lut_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__32935),
            .in2(_gnd_net_),
            .in3(N__32173),
            .lcout(\foc.Look_Up_Table_out1_1_8 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15949 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_9_lut_LC_11_13_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_9_lut_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_9_lut_LC_11_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_9_lut_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__32914),
            .in2(_gnd_net_),
            .in3(N__32161),
            .lcout(\foc.Look_Up_Table_out1_1_9 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15950 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15951 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_10_lut_LC_11_14_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_10_lut_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_10_lut_LC_11_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_10_lut_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__32878),
            .in2(_gnd_net_),
            .in3(N__32146),
            .lcout(\foc.Look_Up_Table_out1_1_10 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_11_lut_LC_11_14_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_11_lut_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_11_lut_LC_11_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_11_lut_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__33262),
            .in2(_gnd_net_),
            .in3(N__32434),
            .lcout(\foc.Look_Up_Table_out1_1_11 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15952 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_12_lut_LC_11_14_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_12_lut_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_12_lut_LC_11_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_12_lut_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__33226),
            .in2(_gnd_net_),
            .in3(N__32431),
            .lcout(\foc.Look_Up_Table_out1_1_12 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15953 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_13_lut_LC_11_14_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_13_lut_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_13_lut_LC_11_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_13_lut_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__33181),
            .in2(_gnd_net_),
            .in3(N__32428),
            .lcout(Look_Up_Table_out1_1_13),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15954 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_14_lut_LC_11_14_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_14_lut_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_14_lut_LC_11_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_14_lut_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__33136),
            .in2(N__44860),
            .in3(N__32425),
            .lcout(Look_Up_Table_out1_1_14),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15955 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n15956 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_15_lut_LC_11_14_5 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_15_lut_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_15_lut_LC_11_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_551_15_lut_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__33091),
            .in2(_gnd_net_),
            .in3(N__32422),
            .lcout(Look_Up_Table_out1_1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i534_2_lut_LC_11_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i534_2_lut_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i534_2_lut_LC_11_14_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i534_2_lut_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32415),
            .lcout(\foc.u_Park_Transform.n785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_2_lut_LC_11_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_2_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_2_lut_LC_11_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_2_lut_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__32352),
            .in2(N__34276),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n75_adj_2123 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\foc.u_Park_Transform.n16948 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_3_lut_LC_11_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_3_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_3_lut_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_3_lut_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__32242),
            .in2(N__34277),
            .in3(N__32233),
            .lcout(\foc.u_Park_Transform.n124_adj_2090 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16948 ),
            .carryout(\foc.u_Park_Transform.n16949 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_4_lut_LC_11_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_4_lut_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_4_lut_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_4_lut_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__34249),
            .in2(N__32230),
            .in3(N__32218),
            .lcout(\foc.u_Park_Transform.n173_adj_2061 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16949 ),
            .carryout(\foc.u_Park_Transform.n16950 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_5_lut_LC_11_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_5_lut_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_5_lut_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_5_lut_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__34243),
            .in2(N__32578),
            .in3(N__32566),
            .lcout(\foc.u_Park_Transform.n222_adj_2049 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16950 ),
            .carryout(\foc.u_Park_Transform.n16951 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_6_lut_LC_11_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_6_lut_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_6_lut_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_6_lut_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__34250),
            .in2(N__32563),
            .in3(N__32551),
            .lcout(\foc.u_Park_Transform.n271_adj_2043 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16951 ),
            .carryout(\foc.u_Park_Transform.n16952 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_7_lut_LC_11_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_7_lut_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_7_lut_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_7_lut_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__34244),
            .in2(N__32548),
            .in3(N__32536),
            .lcout(\foc.u_Park_Transform.n320_adj_2036 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16952 ),
            .carryout(\foc.u_Park_Transform.n16953 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_8_lut_LC_11_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_8_lut_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_8_lut_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_8_lut_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__34251),
            .in2(N__32533),
            .in3(N__32521),
            .lcout(\foc.u_Park_Transform.n369_adj_2026 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16953 ),
            .carryout(\foc.u_Park_Transform.n16954 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_9_lut_LC_11_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_9_lut_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_9_lut_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_9_lut_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__34245),
            .in2(N__32518),
            .in3(N__32506),
            .lcout(\foc.u_Park_Transform.n418 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16954 ),
            .carryout(\foc.u_Park_Transform.n16955 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_10_lut_LC_11_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_10_lut_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_10_lut_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_10_lut_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__34280),
            .in2(N__32503),
            .in3(N__32488),
            .lcout(\foc.u_Park_Transform.n467 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\foc.u_Park_Transform.n16956 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_11_lut_LC_11_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_11_lut_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_11_lut_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_11_lut_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__32485),
            .in2(N__34292),
            .in3(N__32476),
            .lcout(\foc.u_Park_Transform.n516 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16956 ),
            .carryout(\foc.u_Park_Transform.n16957 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_12_lut_LC_11_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_12_lut_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_12_lut_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_12_lut_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__34284),
            .in2(N__32473),
            .in3(N__32461),
            .lcout(\foc.u_Park_Transform.n565_adj_2020 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16957 ),
            .carryout(\foc.u_Park_Transform.n16958 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_13_lut_LC_11_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_13_lut_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_13_lut_LC_11_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_13_lut_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__32458),
            .in2(N__34293),
            .in3(N__32449),
            .lcout(\foc.u_Park_Transform.n614 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16958 ),
            .carryout(\foc.u_Park_Transform.n16959 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_14_lut_LC_11_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_14_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_14_lut_LC_11_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_14_lut_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__32600),
            .in2(N__34294),
            .in3(N__32629),
            .lcout(\foc.u_Park_Transform.n663 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16959 ),
            .carryout(\foc.u_Park_Transform.n16960 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_15_lut_LC_11_16_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_15_lut_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_15_lut_LC_11_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_15_lut_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__34291),
            .in2(N__32607),
            .in3(N__32626),
            .lcout(\foc.u_Park_Transform.n712 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16960 ),
            .carryout(\foc.u_Park_Transform.n16961 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_16_lut_LC_11_16_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_16_lut_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_569_16_lut_LC_11_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_569_16_lut_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__32623),
            .in2(N__32608),
            .in3(N__32584),
            .lcout(\foc.u_Park_Transform.n770 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16961 ),
            .carryout(\foc.u_Park_Transform.n771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n771_THRU_LUT4_0_LC_11_16_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n771_THRU_LUT4_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n771_THRU_LUT4_0_LC_11_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n771_THRU_LUT4_0_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32581),
            .lcout(\foc.u_Park_Transform.n771_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_2_LC_11_17_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_2_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_2_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_2_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__36660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_3_LC_11_17_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_3_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_3_LC_11_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_3_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__32848),
            .in2(N__36415),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17358 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_4_LC_11_17_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_4_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_4_LC_11_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_4_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__36388),
            .in2(N__32861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17359 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_5_LC_11_17_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_5_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_5_LC_11_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_5_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__32852),
            .in2(N__36364),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17360 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_6_LC_11_17_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_6_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_6_LC_11_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_6_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__36334),
            .in2(N__32862),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17361 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_7_LC_11_17_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_7_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_7_LC_11_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_7_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__32856),
            .in2(N__36310),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17362 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_8_lut_LC_11_17_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_8_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_8_lut_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_8_lut_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__36286),
            .in2(N__32863),
            .in3(N__32866),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3008 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17363 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_9_lut_LC_11_17_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_9_lut_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_9_lut_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_9_lut_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__32860),
            .in2(N__36265),
            .in3(N__32824),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3108 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17364 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17365 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_10_lut_LC_11_18_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_10_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_10_lut_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5955_10_lut_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__36622),
            .in2(_gnd_net_),
            .in3(N__32821),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3211 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_LUT4_0_LC_11_18_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_LUT4_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_LUT4_0_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_LUT4_0_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32818),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3212_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_2_lut_LC_11_19_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_2_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_2_lut_LC_11_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_2_lut_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__32815),
            .in2(N__32804),
            .in3(_gnd_net_),
            .lcout(\foc.Look_Up_Table_out1_1_0 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_3_lut_LC_11_19_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_3_lut_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_3_lut_LC_11_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_3_lut_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__32659),
            .in2(_gnd_net_),
            .in3(N__32650),
            .lcout(\foc.Look_Up_Table_out1_1_1 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17490 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_4_lut_LC_11_19_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_4_lut_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_4_lut_LC_11_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_4_lut_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__32647),
            .in2(_gnd_net_),
            .in3(N__32632),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_34 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17491 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_5_lut_LC_11_19_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_5_lut_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_5_lut_LC_11_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_5_lut_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__36601),
            .in2(N__33052),
            .in3(N__33034),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_35 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17492 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_6_lut_LC_11_19_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_6_lut_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_6_lut_LC_11_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_6_lut_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__34837),
            .in2(N__36583),
            .in3(N__33022),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_36 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17493 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_7_lut_LC_11_19_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_7_lut_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_7_lut_LC_11_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_7_lut_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__33019),
            .in2(N__34825),
            .in3(N__33004),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_37 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17494 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_8_lut_LC_11_19_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_8_lut_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_8_lut_LC_11_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_8_lut_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__33001),
            .in2(N__32989),
            .in3(N__32968),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_38 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17495 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_9_lut_LC_11_19_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_9_lut_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_9_lut_LC_11_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_9_lut_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__33439),
            .in2(N__32965),
            .in3(N__32938),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_39 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17496 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17497 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_10_lut_LC_11_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_10_lut_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_10_lut_LC_11_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_10_lut_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__33376),
            .in2(N__33748),
            .in3(N__32926),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_40 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_11_lut_LC_11_20_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_11_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_11_lut_LC_11_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_11_lut_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__32923),
            .in2(N__33361),
            .in3(N__32905),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_41 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17498 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_12_lut_LC_11_20_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_12_lut_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_12_lut_LC_11_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_12_lut_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__32902),
            .in2(N__32890),
            .in3(N__32869),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_42 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17499 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_13_lut_LC_11_20_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_13_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_13_lut_LC_11_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_13_lut_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__33286),
            .in2(N__33277),
            .in3(N__33253),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_43 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17500 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_14_lut_LC_11_20_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_14_lut_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_14_lut_LC_11_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_14_lut_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__33250),
            .in2(N__33238),
            .in3(N__33214),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_44 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17501 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_15_lut_LC_11_20_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_15_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_15_lut_LC_11_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_15_lut_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__33211),
            .in2(N__33196),
            .in3(N__33169),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_45 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17502 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_16_lut_LC_11_20_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_16_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_16_lut_LC_11_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_16_lut_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__33166),
            .in2(N__33154),
            .in3(N__33124),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_46 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17503 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17504 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_17_lut_LC_11_20_7 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_17_lut_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_17_lut_LC_11_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_3098_17_lut_LC_11_20_7  (
            .in0(N__33121),
            .in1(N__33106),
            .in2(_gnd_net_),
            .in3(N__33094),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.Look_Up_Table_mul_temp1_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_2_lut_LC_11_21_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_2_lut_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_2_lut_LC_11_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_2_lut_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__33079),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2426 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_3_lut_LC_11_21_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_3_lut_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_3_lut_LC_11_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_3_lut_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__33327),
            .in2(N__33073),
            .in3(N__33064),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2526 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17412 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_4_lut_LC_11_21_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_4_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_4_lut_LC_11_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_4_lut_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__33061),
            .in2(N__33345),
            .in3(N__33055),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2626 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17413 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_5_lut_LC_11_21_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_5_lut_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_5_lut_LC_11_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_5_lut_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__33331),
            .in2(N__33430),
            .in3(N__33421),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2726 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17414 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_6_lut_LC_11_21_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_6_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_6_lut_LC_11_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_6_lut_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__33418),
            .in2(N__33346),
            .in3(N__33412),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2826 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17415 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_7_lut_LC_11_21_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_7_lut_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_7_lut_LC_11_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_7_lut_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__33409),
            .in2(N__33348),
            .in3(N__33403),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2926 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17416 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_8_lut_LC_11_21_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_8_lut_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_8_lut_LC_11_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_8_lut_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__33400),
            .in2(N__33347),
            .in3(N__33394),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3026 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17417 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_9_lut_LC_11_21_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_9_lut_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_9_lut_LC_11_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_9_lut_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__33391),
            .in2(N__33349),
            .in3(N__33385),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3126 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17418 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17419 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_10_lut_LC_11_22_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_10_lut_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_10_lut_LC_11_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5961_10_lut_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__33382),
            .in2(_gnd_net_),
            .in3(N__33367),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3235 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_LUT4_0_LC_11_22_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_LUT4_0_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_LUT4_0_LC_11_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_LUT4_0_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33364),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3236_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_2_lut_LC_11_23_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_2_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_2_lut_LC_11_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_2_lut_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__33344),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2423 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_3_lut_LC_11_23_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_3_lut_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_3_lut_LC_11_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_3_lut_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__33496),
            .in2(N__33652),
            .in3(N__33634),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2523 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17403 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_4_lut_LC_11_23_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_4_lut_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_4_lut_LC_11_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_4_lut_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__33631),
            .in2(N__33513),
            .in3(N__33613),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2623 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17404 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_5_lut_LC_11_23_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_5_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_5_lut_LC_11_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_5_lut_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__33500),
            .in2(N__33610),
            .in3(N__33592),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2723 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17405 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_6_lut_LC_11_23_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_6_lut_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_6_lut_LC_11_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_6_lut_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__33589),
            .in2(N__33514),
            .in3(N__33568),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2823 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17406 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_7_lut_LC_11_23_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_7_lut_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_7_lut_LC_11_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_7_lut_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__33565),
            .in2(N__33516),
            .in3(N__33550),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2923 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17407 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_8_lut_LC_11_23_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_8_lut_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_8_lut_LC_11_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_8_lut_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__33547),
            .in2(N__33515),
            .in3(N__33529),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3023 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17408 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_9_lut_LC_11_23_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_9_lut_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_9_lut_LC_11_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_9_lut_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(N__33526),
            .in2(N__33517),
            .in3(N__33451),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3123 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17409 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17410 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_10_lut_LC_11_24_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_10_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_10_lut_LC_11_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5960_10_lut_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__33448),
            .in2(_gnd_net_),
            .in3(N__33754),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3231 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_LUT4_0_LC_11_24_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_LUT4_0_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_LUT4_0_LC_11_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_LUT4_0_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33751),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3232_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_2_lut_LC_12_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_2_lut_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_2_lut_LC_12_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_2_lut_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__35813),
            .in2(N__36133),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n69 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\foc.u_Park_Transform.n17161 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_3_lut_LC_12_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_3_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_3_lut_LC_12_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_3_lut_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__36124),
            .in2(N__33736),
            .in3(N__33724),
            .lcout(\foc.u_Park_Transform.n118 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17161 ),
            .carryout(\foc.u_Park_Transform.n17162 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_4_lut_LC_12_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_4_lut_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_4_lut_LC_12_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_4_lut_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__36029),
            .in2(N__33721),
            .in3(N__33709),
            .lcout(\foc.u_Park_Transform.n167 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17162 ),
            .carryout(\foc.u_Park_Transform.n17163 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_5_lut_LC_12_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_5_lut_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_5_lut_LC_12_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_5_lut_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__33706),
            .in2(N__36082),
            .in3(N__33697),
            .lcout(\foc.u_Park_Transform.n216 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17163 ),
            .carryout(\foc.u_Park_Transform.n17164 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_6_lut_LC_12_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_6_lut_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_6_lut_LC_12_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_6_lut_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__36033),
            .in2(N__33694),
            .in3(N__33682),
            .lcout(\foc.u_Park_Transform.n265 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17164 ),
            .carryout(\foc.u_Park_Transform.n17165 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_7_lut_LC_12_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_7_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_7_lut_LC_12_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_7_lut_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__33679),
            .in2(N__36083),
            .in3(N__33670),
            .lcout(\foc.u_Park_Transform.n314 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17165 ),
            .carryout(\foc.u_Park_Transform.n17166 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_8_lut_LC_12_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_8_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_8_lut_LC_12_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_8_lut_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__36037),
            .in2(N__33667),
            .in3(N__33655),
            .lcout(\foc.u_Park_Transform.n363 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17166 ),
            .carryout(\foc.u_Park_Transform.n17167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_9_lut_LC_12_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_9_lut_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_9_lut_LC_12_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_9_lut_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__33862),
            .in2(N__36084),
            .in3(N__33853),
            .lcout(\foc.u_Park_Transform.n412 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17167 ),
            .carryout(\foc.u_Park_Transform.n17168 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_10_lut_LC_12_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_10_lut_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_10_lut_LC_12_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_10_lut_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__33850),
            .in2(N__36078),
            .in3(N__33838),
            .lcout(\foc.u_Park_Transform.n461 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\foc.u_Park_Transform.n17169 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_11_lut_LC_12_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_11_lut_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_11_lut_LC_12_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_11_lut_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__36018),
            .in2(N__33835),
            .in3(N__33823),
            .lcout(\foc.u_Park_Transform.n510_adj_2004 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17169 ),
            .carryout(\foc.u_Park_Transform.n17170 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_12_lut_LC_12_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_12_lut_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_12_lut_LC_12_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_12_lut_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__33820),
            .in2(N__36079),
            .in3(N__33811),
            .lcout(\foc.u_Park_Transform.n559_adj_2001 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17170 ),
            .carryout(\foc.u_Park_Transform.n17171 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_13_lut_LC_12_10_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_13_lut_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_13_lut_LC_12_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_13_lut_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__36022),
            .in2(N__33808),
            .in3(N__33796),
            .lcout(\foc.u_Park_Transform.n608 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17171 ),
            .carryout(\foc.u_Park_Transform.n17172 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_14_lut_LC_12_10_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_14_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_14_lut_LC_12_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_14_lut_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__33793),
            .in2(N__36080),
            .in3(N__33784),
            .lcout(\foc.u_Park_Transform.n657 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17172 ),
            .carryout(\foc.u_Park_Transform.n17173 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_15_lut_LC_12_10_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_15_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_15_lut_LC_12_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_15_lut_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__33781),
            .in2(N__36081),
            .in3(N__33772),
            .lcout(\foc.u_Park_Transform.n706 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17173 ),
            .carryout(\foc.u_Park_Transform.n17174 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_16_lut_LC_12_10_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_16_lut_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_16_lut_LC_12_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_567_16_lut_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__35934),
            .in2(N__33769),
            .in3(N__33757),
            .lcout(\foc.u_Park_Transform.n762 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17174 ),
            .carryout(\foc.u_Park_Transform.n763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n763_THRU_LUT4_0_LC_12_10_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n763_THRU_LUT4_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n763_THRU_LUT4_0_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n763_THRU_LUT4_0_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33961),
            .lcout(\foc.u_Park_Transform.n763_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_2_lut_LC_12_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_2_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_2_lut_LC_12_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_2_lut_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__35976),
            .in2(N__37759),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n66 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\foc.u_Park_Transform.n17176 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_3_lut_LC_12_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_3_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_3_lut_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_3_lut_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__37736),
            .in2(N__33958),
            .in3(N__33946),
            .lcout(\foc.u_Park_Transform.n115 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17176 ),
            .carryout(\foc.u_Park_Transform.n17177 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_4_lut_LC_12_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_4_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_4_lut_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_4_lut_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__37737),
            .in2(N__33943),
            .in3(N__33931),
            .lcout(\foc.u_Park_Transform.n164 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17177 ),
            .carryout(\foc.u_Park_Transform.n17178 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_5_lut_LC_12_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_5_lut_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_5_lut_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_5_lut_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__33928),
            .in2(N__37760),
            .in3(N__33919),
            .lcout(\foc.u_Park_Transform.n213 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17178 ),
            .carryout(\foc.u_Park_Transform.n17179 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_6_lut_LC_12_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_6_lut_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_6_lut_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_6_lut_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__37741),
            .in2(N__33916),
            .in3(N__33904),
            .lcout(\foc.u_Park_Transform.n262_adj_1996 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17179 ),
            .carryout(\foc.u_Park_Transform.n17180 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_7_lut_LC_12_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_7_lut_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_7_lut_LC_12_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_7_lut_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__33901),
            .in2(N__37761),
            .in3(N__33892),
            .lcout(\foc.u_Park_Transform.n311 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17180 ),
            .carryout(\foc.u_Park_Transform.n17181 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_8_lut_LC_12_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_8_lut_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_8_lut_LC_12_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_8_lut_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__37745),
            .in2(N__33889),
            .in3(N__33877),
            .lcout(\foc.u_Park_Transform.n360 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17181 ),
            .carryout(\foc.u_Park_Transform.n17182 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_9_lut_LC_12_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_9_lut_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_9_lut_LC_12_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_9_lut_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__33874),
            .in2(N__37762),
            .in3(N__33865),
            .lcout(\foc.u_Park_Transform.n409 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17182 ),
            .carryout(\foc.u_Park_Transform.n17183 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_10_lut_LC_12_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_10_lut_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_10_lut_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_10_lut_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__37643),
            .in2(N__34057),
            .in3(N__34045),
            .lcout(\foc.u_Park_Transform.n458 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\foc.u_Park_Transform.n17184 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_11_lut_LC_12_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_11_lut_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_11_lut_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_11_lut_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__34042),
            .in2(N__37713),
            .in3(N__34033),
            .lcout(\foc.u_Park_Transform.n507_adj_2165 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17184 ),
            .carryout(\foc.u_Park_Transform.n17185 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_12_lut_LC_12_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_12_lut_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_12_lut_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_12_lut_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__37647),
            .in2(N__34030),
            .in3(N__34018),
            .lcout(\foc.u_Park_Transform.n556_adj_2164 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17185 ),
            .carryout(\foc.u_Park_Transform.n17186 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_13_lut_LC_12_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_13_lut_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_13_lut_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_13_lut_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__34015),
            .in2(N__37714),
            .in3(N__34006),
            .lcout(\foc.u_Park_Transform.n605_adj_2163 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17186 ),
            .carryout(\foc.u_Park_Transform.n17187 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_14_lut_LC_12_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_14_lut_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_14_lut_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_14_lut_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__34003),
            .in2(N__37716),
            .in3(N__33994),
            .lcout(\foc.u_Park_Transform.n654_adj_2162 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17187 ),
            .carryout(\foc.u_Park_Transform.n17188 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_15_lut_LC_12_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_15_lut_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_15_lut_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_15_lut_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__33991),
            .in2(N__37715),
            .in3(N__33982),
            .lcout(\foc.u_Park_Transform.n703_adj_2160 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17188 ),
            .carryout(\foc.u_Park_Transform.n17189 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_16_lut_LC_12_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_16_lut_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_16_lut_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_566_16_lut_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__35541),
            .in2(N__33979),
            .in3(N__33967),
            .lcout(\foc.u_Park_Transform.n758_adj_2168 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17189 ),
            .carryout(\foc.u_Park_Transform.n759_adj_2166 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n759_adj_2166_THRU_LUT4_0_LC_12_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n759_adj_2166_THRU_LUT4_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n759_adj_2166_THRU_LUT4_0_LC_12_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n759_adj_2166_THRU_LUT4_0_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33964),
            .lcout(\foc.u_Park_Transform.n759_adj_2166_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i8_2_lut_LC_12_13_0 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i8_2_lut_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i8_2_lut_LC_12_13_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i8_2_lut_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__34083),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i507_2_lut_LC_12_13_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i507_2_lut_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i507_2_lut_LC_12_13_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i507_2_lut_LC_12_13_1  (
            .in0(N__34084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i510_2_lut_LC_12_13_2 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i510_2_lut_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i510_2_lut_LC_12_13_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i510_2_lut_LC_12_13_2  (
            .in0(N__34066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i504_2_lut_LC_12_13_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i504_2_lut_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i504_2_lut_LC_12_13_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i504_2_lut_LC_12_13_3  (
            .in0(N__42714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i513_2_lut_LC_12_13_4 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i513_2_lut_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i513_2_lut_LC_12_13_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i513_2_lut_LC_12_13_4  (
            .in0(N__34075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i12_2_lut_LC_12_13_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i12_2_lut_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i12_2_lut_LC_12_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i12_2_lut_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34074),
            .lcout(\foc.u_Park_Transform.n604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.u_29__I_0_71_inv_0_i4_1_lut_LC_12_13_6 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.u_29__I_0_71_inv_0_i4_1_lut_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.u_29__I_0_71_inv_0_i4_1_lut_LC_12_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.u_29__I_0_71_inv_0_i4_1_lut_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Amp25_out1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i10_2_lut_LC_12_13_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i10_2_lut_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i10_2_lut_LC_12_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i10_2_lut_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34065),
            .lcout(\foc.u_Park_Transform.n601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i498_2_lut_LC_12_14_0 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i498_2_lut_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i498_2_lut_LC_12_14_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i498_2_lut_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36568),
            .lcout(\foc.u_Park_Transform.n737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i2_4_lut_4_lut_LC_12_14_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i2_4_lut_4_lut_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i2_4_lut_4_lut_LC_12_14_1 .LUT_INIT=16'b0010010010110100;
    LogicCell40 \foc.u_Park_Transform.i2_4_lut_4_lut_LC_12_14_1  (
            .in0(N__44188),
            .in1(N__44317),
            .in2(_gnd_net_),
            .in3(N__44394),
            .lcout(\foc.u_Park_Transform.n790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11567_4_lut_4_lut_LC_12_14_2.C_ON=1'b0;
    defparam i11567_4_lut_4_lut_LC_12_14_2.SEQ_MODE=4'b0000;
    defparam i11567_4_lut_4_lut_LC_12_14_2.LUT_INIT=16'b1110110000000000;
    LogicCell40 i11567_4_lut_4_lut_LC_12_14_2 (
            .in0(N__44395),
            .in1(N__44240),
            .in2(_gnd_net_),
            .in3(N__40475),
            .lcout(n4),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_LC_12_14_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_LC_12_14_3 .LUT_INIT=16'b1000111000001100;
    LogicCell40 \foc.u_Park_Transform.i1_3_lut_4_lut_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__44315),
            .in2(N__34366),
            .in3(N__44392),
            .lcout(\foc.u_Park_Transform.n237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i2_2_lut_LC_12_14_6 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i2_2_lut_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i2_2_lut_LC_12_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i2_2_lut_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36567),
            .lcout(\foc.u_Park_Transform.dCurrent_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i2_3_lut_4_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i2_3_lut_4_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i2_3_lut_4_lut_LC_12_14_7 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \foc.u_Park_Transform.i2_3_lut_4_lut_LC_12_14_7  (
            .in0(N__42507),
            .in1(N__44316),
            .in2(_gnd_net_),
            .in3(N__44393),
            .lcout(\foc.u_Park_Transform.n188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_2_lut_LC_12_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_2_lut_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_2_lut_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_2_lut_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__34279),
            .in2(N__35883),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n72_adj_2062 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\foc.u_Park_Transform.n16963 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_3_lut_LC_12_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_3_lut_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_3_lut_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_3_lut_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__34126),
            .in2(N__35884),
            .in3(N__34120),
            .lcout(\foc.u_Park_Transform.n121_adj_2051 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16963 ),
            .carryout(\foc.u_Park_Transform.n16964 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_4_lut_LC_12_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_4_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_4_lut_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_4_lut_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__35838),
            .in2(N__34117),
            .in3(N__34108),
            .lcout(\foc.u_Park_Transform.n170_adj_2048 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16964 ),
            .carryout(\foc.u_Park_Transform.n16965 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_5_lut_LC_12_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_5_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_5_lut_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_5_lut_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__34105),
            .in2(N__35885),
            .in3(N__34099),
            .lcout(\foc.u_Park_Transform.n219_adj_2040 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16965 ),
            .carryout(\foc.u_Park_Transform.n16966 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_6_lut_LC_12_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_6_lut_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_6_lut_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_6_lut_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__35842),
            .in2(N__34096),
            .in3(N__34087),
            .lcout(\foc.u_Park_Transform.n268_adj_2027 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16966 ),
            .carryout(\foc.u_Park_Transform.n16967 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_7_lut_LC_12_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_7_lut_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_7_lut_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_7_lut_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__34453),
            .in2(N__35886),
            .in3(N__34447),
            .lcout(\foc.u_Park_Transform.n317_adj_2021 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16967 ),
            .carryout(\foc.u_Park_Transform.n16968 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_8_lut_LC_12_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_8_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_8_lut_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_8_lut_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__35846),
            .in2(N__34444),
            .in3(N__34435),
            .lcout(\foc.u_Park_Transform.n366_adj_2013 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16968 ),
            .carryout(\foc.u_Park_Transform.n16969 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_9_lut_LC_12_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_9_lut_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_9_lut_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_9_lut_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__34432),
            .in2(N__35887),
            .in3(N__34426),
            .lcout(\foc.u_Park_Transform.n415 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16969 ),
            .carryout(\foc.u_Park_Transform.n16970 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_10_lut_LC_12_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_10_lut_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_10_lut_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_10_lut_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__35850),
            .in2(N__34423),
            .in3(N__34414),
            .lcout(\foc.u_Park_Transform.n464 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\foc.u_Park_Transform.n16971 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_11_lut_LC_12_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_11_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_11_lut_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_11_lut_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__34411),
            .in2(N__35888),
            .in3(N__34405),
            .lcout(\foc.u_Park_Transform.n513 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16971 ),
            .carryout(\foc.u_Park_Transform.n16972 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_12_lut_LC_12_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_12_lut_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_12_lut_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_12_lut_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__35854),
            .in2(N__34402),
            .in3(N__34393),
            .lcout(\foc.u_Park_Transform.n562 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16972 ),
            .carryout(\foc.u_Park_Transform.n16973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_13_lut_LC_12_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_13_lut_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_13_lut_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_13_lut_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__34390),
            .in2(N__35889),
            .in3(N__34384),
            .lcout(\foc.u_Park_Transform.n611_adj_2107 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16973 ),
            .carryout(\foc.u_Park_Transform.n16974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_14_lut_LC_12_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_14_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_14_lut_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_14_lut_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__34381),
            .in2(N__35891),
            .in3(N__34375),
            .lcout(\foc.u_Park_Transform.n660_adj_2091 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16974 ),
            .carryout(\foc.u_Park_Transform.n16975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_15_lut_LC_12_16_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_15_lut_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_15_lut_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_15_lut_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__34372),
            .in2(N__35890),
            .in3(N__34507),
            .lcout(\foc.u_Park_Transform.n709_adj_2066 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16975 ),
            .carryout(\foc.u_Park_Transform.n16976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_16_lut_LC_12_16_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_16_lut_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_568_16_lut_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_568_16_lut_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__34504),
            .in2(N__34483),
            .in3(N__34474),
            .lcout(\foc.u_Park_Transform.n766_adj_2053 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16976 ),
            .carryout(\foc.u_Park_Transform.n767_adj_2041 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n767_adj_2041_THRU_LUT4_0_LC_12_16_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n767_adj_2041_THRU_LUT4_0_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n767_adj_2041_THRU_LUT4_0_LC_12_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n767_adj_2041_THRU_LUT4_0_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34471),
            .lcout(\foc.u_Park_Transform.n767_adj_2041_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_1_LC_12_17_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_1_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_1_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Park_Transform.add_1232_1_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__37989),
            .in2(N__37993),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\foc.u_Park_Transform.n16900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_2_lut_LC_12_17_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_2_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_2_lut_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_2_lut_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__40447),
            .in2(_gnd_net_),
            .in3(N__34468),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_15 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16900 ),
            .carryout(\foc.u_Park_Transform.n16901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_3_lut_LC_12_17_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_3_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_3_lut_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_3_lut_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__40141),
            .in2(N__37966),
            .in3(N__34465),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_16 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16901 ),
            .carryout(\foc.u_Park_Transform.n16902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_4_lut_LC_12_17_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_4_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_4_lut_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_4_lut_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__42763),
            .in2(N__40123),
            .in3(N__34462),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_17 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16902 ),
            .carryout(\foc.u_Park_Transform.n16903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_5_lut_LC_12_17_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_5_lut_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_5_lut_LC_12_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_5_lut_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__39931),
            .in2(N__42745),
            .in3(N__34459),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_18 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16903 ),
            .carryout(\foc.u_Park_Transform.n16904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_6_lut_LC_12_17_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_6_lut_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_6_lut_LC_12_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_6_lut_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__37813),
            .in2(N__40105),
            .in3(N__34456),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_19 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16904 ),
            .carryout(\foc.u_Park_Transform.n16905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_7_lut_LC_12_17_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_7_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_7_lut_LC_12_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_7_lut_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__35530),
            .in2(N__37795),
            .in3(N__34678),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_20 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16905 ),
            .carryout(\foc.u_Park_Transform.n16906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_8_lut_LC_12_17_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_8_lut_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_8_lut_LC_12_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_8_lut_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__35515),
            .in2(N__35908),
            .in3(N__34675),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_21 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16906 ),
            .carryout(\foc.u_Park_Transform.n16907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_9_lut_LC_12_18_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_9_lut_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_9_lut_LC_12_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_9_lut_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__34672),
            .in2(N__36487),
            .in3(N__34663),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_22 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\foc.u_Park_Transform.n16908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_10_lut_LC_12_18_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_10_lut_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_10_lut_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_10_lut_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__34660),
            .in2(N__34651),
            .in3(N__34639),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_23 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16908 ),
            .carryout(\foc.u_Park_Transform.n16909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_11_lut_LC_12_18_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_11_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_11_lut_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_11_lut_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__34636),
            .in2(N__34624),
            .in3(N__34612),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_24 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16909 ),
            .carryout(\foc.u_Park_Transform.n16910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_12_lut_LC_12_18_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_12_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_12_lut_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_12_lut_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__34609),
            .in2(N__34600),
            .in3(N__34585),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_25 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16910 ),
            .carryout(\foc.u_Park_Transform.n16911 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_13_lut_LC_12_18_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_13_lut_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_13_lut_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_13_lut_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__34582),
            .in2(N__34570),
            .in3(N__34558),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_26 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16911 ),
            .carryout(\foc.u_Park_Transform.n16912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_14_lut_LC_12_18_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_14_lut_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_14_lut_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_14_lut_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__34555),
            .in2(N__34543),
            .in3(N__34528),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_27 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16912 ),
            .carryout(\foc.u_Park_Transform.n16913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_15_lut_LC_12_18_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1232_15_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_15_lut_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1232_15_lut_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__35316),
            .in2(N__34525),
            .in3(N__34510),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_28 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16913 ),
            .carryout(\foc.u_Park_Transform.n16914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1232_16_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.add_1232_16_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1232_16_lut_LC_12_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Park_Transform.add_1232_16_lut_LC_12_18_7  (
            .in0(N__36537),
            .in1(N__44467),
            .in2(_gnd_net_),
            .in3(N__34801),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_2_lut_LC_12_19_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_2_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_2_lut_LC_12_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_2_lut_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__34798),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2414 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_3_lut_LC_12_19_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_3_lut_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_3_lut_LC_12_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_3_lut_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__36447),
            .in2(N__34756),
            .in3(N__34744),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2514 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17376 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_4_lut_LC_12_19_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_4_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_4_lut_LC_12_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_4_lut_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__34741),
            .in2(N__36467),
            .in3(N__34732),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2614 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17377 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_5_lut_LC_12_19_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_5_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_5_lut_LC_12_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_5_lut_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__36451),
            .in2(N__34729),
            .in3(N__34717),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2714 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17378 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_6_lut_LC_12_19_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_6_lut_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_6_lut_LC_12_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_6_lut_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__34714),
            .in2(N__36468),
            .in3(N__34705),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2814 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17379 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_7_lut_LC_12_19_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_7_lut_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_7_lut_LC_12_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_7_lut_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__34702),
            .in2(N__36470),
            .in3(N__34693),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2914 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17380 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_8_lut_LC_12_19_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_8_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_8_lut_LC_12_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_8_lut_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__34690),
            .in2(N__36469),
            .in3(N__34681),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3014 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17381 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_9_lut_LC_12_19_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_9_lut_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_9_lut_LC_12_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_9_lut_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__34861),
            .in2(N__36471),
            .in3(N__34852),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3114 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17382 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17383 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_10_lut_LC_12_20_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_10_lut_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_10_lut_LC_12_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5957_10_lut_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__34849),
            .in2(_gnd_net_),
            .in3(N__34831),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3219 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_LUT4_0_LC_12_20_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_LUT4_0_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_LUT4_0_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_LUT4_0_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34828),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3220_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_12_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__66260),
            .in2(N__66515),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n78_adj_617 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_12_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__36526),
            .in2(N__66517),
            .in3(N__34816),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n127_adj_615 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17656 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_12_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__66464),
            .in2(N__36517),
            .in3(N__34813),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n176_adj_613 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17657 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_12_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__36502),
            .in2(N__66518),
            .in3(N__34810),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n225_adj_611 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17658 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_12_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__66468),
            .in2(N__36802),
            .in3(N__34807),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n274_adj_609 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17659 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_12_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_12_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__36787),
            .in2(N__66519),
            .in3(N__34804),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n323_adj_607 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17660 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_12_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_12_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(N__36772),
            .in2(N__66516),
            .in3(N__34885),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n372 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17661 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_12_22_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_12_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__36760),
            .in2(N__66520),
            .in3(N__34882),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n421 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17662 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_12_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_12_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__36745),
            .in2(N__66574),
            .in3(N__34879),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n470 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_12_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__36733),
            .in2(N__66575),
            .in3(N__34876),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n519 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17664 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_12_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__66534),
            .in2(N__36720),
            .in3(N__34873),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n568 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17665 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_12_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__36716),
            .in2(N__66576),
            .in3(N__34870),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n617 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17666 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_12_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__45457),
            .in2(N__36721),
            .in3(N__34867),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n774 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17667 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_LUT4_0_LC_12_23_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_LUT4_0_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_LUT4_0_LC_12_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_LUT4_0_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34864),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_12_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_12_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__66538),
            .in2(N__66888),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n75_adj_618 ),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_12_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_12_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(N__34981),
            .in2(N__66923),
            .in3(N__34972),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n124_adj_616 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18107 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_12_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__34969),
            .in2(N__66889),
            .in3(N__34960),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n173_adj_614 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18108 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_12_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_12_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__34957),
            .in2(N__66924),
            .in3(N__34948),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n222_adj_612 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18109 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_12_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_12_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__34945),
            .in2(N__66890),
            .in3(N__34936),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n271_adj_610 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18110 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_12_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_12_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__34933),
            .in2(N__66925),
            .in3(N__34924),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n320_adj_608 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18111 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_12_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_12_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__34921),
            .in2(N__66891),
            .in3(N__34912),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n369_adj_606 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18112 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_12_24_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_12_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_12_24_7  (
            .in0(_gnd_net_),
            .in1(N__34909),
            .in2(N__66926),
            .in3(N__34900),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n418_adj_605 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18113 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_12_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_12_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__34897),
            .in2(N__66927),
            .in3(N__34888),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n467_adj_604 ),
            .ltout(),
            .carryin(bfn_12_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_12_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_12_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_12_25_1  (
            .in0(_gnd_net_),
            .in1(N__35053),
            .in2(N__66930),
            .in3(N__35044),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n516_adj_603 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18115 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_12_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_12_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__35041),
            .in2(N__66928),
            .in3(N__35032),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n565_adj_602 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18116 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18117 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_12_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_12_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(N__35029),
            .in2(N__66931),
            .in3(N__35020),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n614_adj_601 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18117 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18118 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_12_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_12_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(N__35003),
            .in2(N__66929),
            .in3(N__35017),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n663_adj_600 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18118 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18119 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_12_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_12_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(N__66913),
            .in2(N__35010),
            .in3(N__35014),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n712_adj_599 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18119 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18120 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_12_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_12_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__45484),
            .in2(N__35011),
            .in3(N__34987),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n770_adj_597 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18120 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_LUT4_0_LC_12_25_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_LUT4_0_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_LUT4_0_LC_12_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_LUT4_0_LC_12_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34984),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_adj_598_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i18_1_lut_LC_13_6_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i18_1_lut_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i18_1_lut_LC_13_6_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i18_1_lut_LC_13_6_0  (
            .in0(N__37354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i20_1_lut_LC_13_6_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i20_1_lut_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i20_1_lut_LC_13_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i20_1_lut_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37318),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n14_adj_517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i21_1_lut_LC_13_6_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i21_1_lut_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i21_1_lut_LC_13_6_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i21_1_lut_LC_13_6_3  (
            .in0(N__37300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i22_1_lut_LC_13_6_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i22_1_lut_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i22_1_lut_LC_13_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i22_1_lut_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37282),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n12_adj_516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i23_1_lut_LC_13_6_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i23_1_lut_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i23_1_lut_LC_13_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i23_1_lut_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37264),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i24_1_lut_LC_13_6_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i24_1_lut_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i24_1_lut_LC_13_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i24_1_lut_LC_13_6_6  (
            .in0(N__37246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i25_1_lut_LC_13_6_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i25_1_lut_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i25_1_lut_LC_13_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i25_1_lut_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37228),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_1_LC_13_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_1_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_1_LC_13_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_Park_Transform.add_1234_1_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__39645),
            .in2(N__39649),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\foc.u_Park_Transform.n17083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_2_lut_LC_13_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_2_lut_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_2_lut_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_2_lut_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__40462),
            .in2(_gnd_net_),
            .in3(N__35065),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_15 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17083 ),
            .carryout(\foc.u_Park_Transform.n17084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_3_lut_LC_13_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_3_lut_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_3_lut_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_3_lut_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__39907),
            .in2(N__39622),
            .in3(N__35062),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_16 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17084 ),
            .carryout(\foc.u_Park_Transform.n17085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_4_lut_LC_13_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_4_lut_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_4_lut_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_4_lut_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__37483),
            .in2(N__39889),
            .in3(N__35059),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_17 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17085 ),
            .carryout(\foc.u_Park_Transform.n17086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_5_lut_LC_13_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_5_lut_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_5_lut_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_5_lut_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__42256),
            .in2(N__37777),
            .in3(N__35056),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_18 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17086 ),
            .carryout(\foc.u_Park_Transform.n17087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_6_lut_LC_13_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_6_lut_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_6_lut_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_6_lut_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__35494),
            .in2(N__42238),
            .in3(N__35236),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_19 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17087 ),
            .carryout(\foc.u_Park_Transform.n17088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_7_lut_LC_13_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_7_lut_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_7_lut_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_7_lut_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__35233),
            .in2(N__35479),
            .in3(N__35221),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_20 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17088 ),
            .carryout(\foc.u_Park_Transform.n17089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_8_lut_LC_13_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_8_lut_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_8_lut_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_8_lut_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__35218),
            .in2(N__35206),
            .in3(N__35197),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_21 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17089 ),
            .carryout(\foc.u_Park_Transform.n17090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_9_lut_LC_13_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_9_lut_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_9_lut_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_9_lut_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__35194),
            .in2(N__35185),
            .in3(N__35176),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_22 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\foc.u_Park_Transform.n17091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_10_lut_LC_13_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_10_lut_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_10_lut_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_10_lut_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__35173),
            .in2(N__35161),
            .in3(N__35149),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_23 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17091 ),
            .carryout(\foc.u_Park_Transform.n17092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_11_lut_LC_13_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_11_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_11_lut_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_11_lut_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__35146),
            .in2(N__35134),
            .in3(N__35119),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_24 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17092 ),
            .carryout(\foc.u_Park_Transform.n17093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_12_lut_LC_13_10_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_12_lut_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_12_lut_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_12_lut_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__35116),
            .in2(N__35107),
            .in3(N__35092),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_25 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17093 ),
            .carryout(\foc.u_Park_Transform.n17094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_13_lut_LC_13_10_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_13_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_13_lut_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_13_lut_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__35089),
            .in2(N__35080),
            .in3(N__35068),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_26 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17094 ),
            .carryout(\foc.u_Park_Transform.n17095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_14_lut_LC_13_10_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_14_lut_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_14_lut_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_14_lut_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__35350),
            .in2(N__35338),
            .in3(N__35326),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_27 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17095 ),
            .carryout(\foc.u_Park_Transform.n17096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_15_lut_LC_13_10_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_1234_15_lut_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_15_lut_LC_13_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_1234_15_lut_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__35323),
            .in2(N__35302),
            .in3(N__35287),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_28 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17096 ),
            .carryout(\foc.u_Park_Transform.n17097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_1234_16_lut_LC_13_10_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.add_1234_16_lut_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_1234_16_lut_LC_13_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Park_Transform.add_1234_16_lut_LC_13_10_7  (
            .in0(N__44463),
            .in1(N__36544),
            .in2(_gnd_net_),
            .in3(N__35284),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_2_lut_LC_13_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_2_lut_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_2_lut_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_2_lut_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__37754),
            .in2(N__41690),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n63_adj_2158 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\foc.u_Park_Transform.n17191 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_3_lut_LC_13_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_3_lut_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_3_lut_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_3_lut_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__35281),
            .in2(N__41691),
            .in3(N__35275),
            .lcout(\foc.u_Park_Transform.n112_adj_2157 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17191 ),
            .carryout(\foc.u_Park_Transform.n17192 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_4_lut_LC_13_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_4_lut_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_4_lut_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_4_lut_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__41666),
            .in2(N__35272),
            .in3(N__35263),
            .lcout(\foc.u_Park_Transform.n161_adj_2156 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17192 ),
            .carryout(\foc.u_Park_Transform.n17193 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_5_lut_LC_13_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_5_lut_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_5_lut_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_5_lut_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__41660),
            .in2(N__35260),
            .in3(N__35251),
            .lcout(\foc.u_Park_Transform.n210_adj_2155 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17193 ),
            .carryout(\foc.u_Park_Transform.n17194 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_6_lut_LC_13_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_6_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_6_lut_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_6_lut_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__41667),
            .in2(N__35248),
            .in3(N__35239),
            .lcout(\foc.u_Park_Transform.n259_adj_2154 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17194 ),
            .carryout(\foc.u_Park_Transform.n17195 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_7_lut_LC_13_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_7_lut_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_7_lut_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_7_lut_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__41661),
            .in2(N__35449),
            .in3(N__35440),
            .lcout(\foc.u_Park_Transform.n308_adj_2153 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17195 ),
            .carryout(\foc.u_Park_Transform.n17196 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_8_lut_LC_13_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_8_lut_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_8_lut_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_8_lut_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__41668),
            .in2(N__35437),
            .in3(N__35428),
            .lcout(\foc.u_Park_Transform.n357_adj_2151 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17196 ),
            .carryout(\foc.u_Park_Transform.n17197 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_9_lut_LC_13_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_9_lut_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_9_lut_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_9_lut_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__41662),
            .in2(N__35425),
            .in3(N__35416),
            .lcout(\foc.u_Park_Transform.n406_adj_2150 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17197 ),
            .carryout(\foc.u_Park_Transform.n17198 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_10_lut_LC_13_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_10_lut_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_10_lut_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_10_lut_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__35413),
            .in2(N__41651),
            .in3(N__35407),
            .lcout(\foc.u_Park_Transform.n455_adj_2148 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\foc.u_Park_Transform.n17199 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_11_lut_LC_13_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_11_lut_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_11_lut_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_11_lut_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__41600),
            .in2(N__35404),
            .in3(N__35395),
            .lcout(\foc.u_Park_Transform.n504_adj_2147 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17199 ),
            .carryout(\foc.u_Park_Transform.n17200 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_12_lut_LC_13_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_12_lut_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_12_lut_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_12_lut_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__35392),
            .in2(N__41652),
            .in3(N__35386),
            .lcout(\foc.u_Park_Transform.n553_adj_2146 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17200 ),
            .carryout(\foc.u_Park_Transform.n17201 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_13_lut_LC_13_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_13_lut_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_13_lut_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_13_lut_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__41604),
            .in2(N__35383),
            .in3(N__35374),
            .lcout(\foc.u_Park_Transform.n602_adj_2144 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17201 ),
            .carryout(\foc.u_Park_Transform.n17202 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_14_lut_LC_13_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_14_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_14_lut_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_14_lut_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__35371),
            .in2(N__41653),
            .in3(N__35365),
            .lcout(\foc.u_Park_Transform.n651_adj_2143 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17202 ),
            .carryout(\foc.u_Park_Transform.n17203 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_15_lut_LC_13_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_15_lut_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_15_lut_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_15_lut_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__41608),
            .in2(N__35362),
            .in3(N__35353),
            .lcout(\foc.u_Park_Transform.n700_adj_2141 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17203 ),
            .carryout(\foc.u_Park_Transform.n17204 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_16_lut_LC_13_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_16_lut_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_16_lut_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_565_16_lut_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__37833),
            .in2(N__35503),
            .in3(N__35485),
            .lcout(\foc.u_Park_Transform.n754_adj_2159 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17204 ),
            .carryout(\foc.u_Park_Transform.n755_adj_2161 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n755_adj_2161_THRU_LUT4_0_LC_13_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n755_adj_2161_THRU_LUT4_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n755_adj_2161_THRU_LUT4_0_LC_13_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n755_adj_2161_THRU_LUT4_0_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35482),
            .lcout(\foc.u_Park_Transform.n755_adj_2161_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_2_lut_LC_13_13_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_2_lut_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_2_lut_LC_13_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_2_lut_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__36085),
            .in2(N__37755),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n66_adj_2033 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\foc.u_Park_Transform.n16993 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_3_lut_LC_13_13_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_3_lut_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_3_lut_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_3_lut_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__37720),
            .in2(N__35707),
            .in3(N__35467),
            .lcout(\foc.u_Park_Transform.n115_adj_2028 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16993 ),
            .carryout(\foc.u_Park_Transform.n16994 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_4_lut_LC_13_13_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_4_lut_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_4_lut_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_4_lut_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__37721),
            .in2(N__35689),
            .in3(N__35464),
            .lcout(\foc.u_Park_Transform.n164_adj_2014 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16994 ),
            .carryout(\foc.u_Park_Transform.n16995 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_5_lut_LC_13_13_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_5_lut_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_5_lut_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_5_lut_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__35665),
            .in2(N__37756),
            .in3(N__35461),
            .lcout(\foc.u_Park_Transform.n213_adj_1999 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16995 ),
            .carryout(\foc.u_Park_Transform.n16996 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_6_lut_LC_13_13_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_6_lut_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_6_lut_LC_13_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_6_lut_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__37725),
            .in2(N__35647),
            .in3(N__35458),
            .lcout(\foc.u_Park_Transform.n262 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16996 ),
            .carryout(\foc.u_Park_Transform.n16997 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_7_lut_LC_13_13_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_7_lut_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_7_lut_LC_13_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_7_lut_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__35623),
            .in2(N__37757),
            .in3(N__35455),
            .lcout(\foc.u_Park_Transform.n311_adj_2022 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16997 ),
            .carryout(\foc.u_Park_Transform.n16998 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_8_lut_LC_13_13_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_8_lut_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_8_lut_LC_13_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_8_lut_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__37729),
            .in2(N__35605),
            .in3(N__35452),
            .lcout(\foc.u_Park_Transform.n360_adj_2009 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16998 ),
            .carryout(\foc.u_Park_Transform.n16999 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_9_lut_LC_13_13_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_9_lut_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_9_lut_LC_13_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_9_lut_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__35581),
            .in2(N__37758),
            .in3(N__35563),
            .lcout(\foc.u_Park_Transform.n409_adj_1997 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16999 ),
            .carryout(\foc.u_Park_Transform.n17000 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_10_lut_LC_13_14_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_10_lut_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_10_lut_LC_13_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_10_lut_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__37696),
            .in2(N__36250),
            .in3(N__35560),
            .lcout(\foc.u_Park_Transform.n458_adj_2093 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\foc.u_Park_Transform.n17001 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_11_lut_LC_13_14_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_11_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_11_lut_LC_13_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_11_lut_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__36229),
            .in2(N__37750),
            .in3(N__35557),
            .lcout(\foc.u_Park_Transform.n507 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17001 ),
            .carryout(\foc.u_Park_Transform.n17002 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_12_lut_LC_13_14_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_12_lut_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_12_lut_LC_13_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_12_lut_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__37700),
            .in2(N__36211),
            .in3(N__35554),
            .lcout(\foc.u_Park_Transform.n556 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17002 ),
            .carryout(\foc.u_Park_Transform.n17003 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_13_lut_LC_13_14_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_13_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_13_lut_LC_13_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_13_lut_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__36187),
            .in2(N__37751),
            .in3(N__35551),
            .lcout(\foc.u_Park_Transform.n605 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17003 ),
            .carryout(\foc.u_Park_Transform.n17004 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_14_lut_LC_13_14_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_14_lut_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_14_lut_LC_13_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_14_lut_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__36169),
            .in2(N__37753),
            .in3(N__35548),
            .lcout(\foc.u_Park_Transform.n654 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17004 ),
            .carryout(\foc.u_Park_Transform.n17005 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_15_lut_LC_13_14_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_15_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_15_lut_LC_13_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_15_lut_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__36151),
            .in2(N__37752),
            .in3(N__35545),
            .lcout(\foc.u_Park_Transform.n703 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17005 ),
            .carryout(\foc.u_Park_Transform.n17006 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_16_lut_LC_13_14_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_16_lut_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_566_16_lut_LC_13_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_566_16_lut_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__35542),
            .in2(N__35956),
            .in3(N__35521),
            .lcout(\foc.u_Park_Transform.n758 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17006 ),
            .carryout(\foc.u_Park_Transform.n759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n759_THRU_LUT4_0_LC_13_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n759_THRU_LUT4_0_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n759_THRU_LUT4_0_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n759_THRU_LUT4_0_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35518),
            .lcout(\foc.u_Park_Transform.n759_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_2_lut_LC_13_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_2_lut_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_2_lut_LC_13_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_2_lut_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__36091),
            .in2(N__35892),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n69_adj_2059 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\foc.u_Park_Transform.n16978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_3_lut_LC_13_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_3_lut_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_3_lut_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_3_lut_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__35695),
            .in2(N__36125),
            .in3(N__35677),
            .lcout(\foc.u_Park_Transform.n118_adj_2037 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16978 ),
            .carryout(\foc.u_Park_Transform.n16979 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_4_lut_LC_13_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_4_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_4_lut_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_4_lut_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__36095),
            .in2(N__35674),
            .in3(N__35656),
            .lcout(\foc.u_Park_Transform.n167_adj_2029 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16979 ),
            .carryout(\foc.u_Park_Transform.n16980 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_5_lut_LC_13_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_5_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_5_lut_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_5_lut_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__35653),
            .in2(N__36126),
            .in3(N__35635),
            .lcout(\foc.u_Park_Transform.n216_adj_2025 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16980 ),
            .carryout(\foc.u_Park_Transform.n16981 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_6_lut_LC_13_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_6_lut_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_6_lut_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_6_lut_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__36099),
            .in2(N__35632),
            .in3(N__35614),
            .lcout(\foc.u_Park_Transform.n265_adj_2023 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16981 ),
            .carryout(\foc.u_Park_Transform.n16982 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_7_lut_LC_13_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_7_lut_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_7_lut_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_7_lut_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__35611),
            .in2(N__36127),
            .in3(N__35593),
            .lcout(\foc.u_Park_Transform.n314_adj_2010 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16982 ),
            .carryout(\foc.u_Park_Transform.n16983 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_8_lut_LC_13_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_8_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_8_lut_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_8_lut_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__36103),
            .in2(N__35590),
            .in3(N__35572),
            .lcout(\foc.u_Park_Transform.n363_adj_1998 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16983 ),
            .carryout(\foc.u_Park_Transform.n16984 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_9_lut_LC_13_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_9_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_9_lut_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_9_lut_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__35569),
            .in2(N__36128),
            .in3(N__36241),
            .lcout(\foc.u_Park_Transform.n412_adj_1995 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16984 ),
            .carryout(\foc.u_Park_Transform.n16985 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_10_lut_LC_13_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_10_lut_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_10_lut_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_10_lut_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__36107),
            .in2(N__36238),
            .in3(N__36220),
            .lcout(\foc.u_Park_Transform.n461_adj_2007 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\foc.u_Park_Transform.n16986 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_11_lut_LC_13_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_11_lut_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_11_lut_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_11_lut_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__36217),
            .in2(N__36129),
            .in3(N__36199),
            .lcout(\foc.u_Park_Transform.n510 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16986 ),
            .carryout(\foc.u_Park_Transform.n16987 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_12_lut_LC_13_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_12_lut_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_12_lut_LC_13_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_12_lut_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__36111),
            .in2(N__36196),
            .in3(N__36178),
            .lcout(\foc.u_Park_Transform.n559 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16987 ),
            .carryout(\foc.u_Park_Transform.n16988 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_13_lut_LC_13_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_13_lut_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_13_lut_LC_13_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_13_lut_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__36175),
            .in2(N__36130),
            .in3(N__36160),
            .lcout(\foc.u_Park_Transform.n608_adj_2067 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16988 ),
            .carryout(\foc.u_Park_Transform.n16989 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_14_lut_LC_13_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_14_lut_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_14_lut_LC_13_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_14_lut_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__36157),
            .in2(N__36132),
            .in3(N__36142),
            .lcout(\foc.u_Park_Transform.n657_adj_2064 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16989 ),
            .carryout(\foc.u_Park_Transform.n16990 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_15_lut_LC_13_16_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_15_lut_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_15_lut_LC_13_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_15_lut_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__36139),
            .in2(N__36131),
            .in3(N__35944),
            .lcout(\foc.u_Park_Transform.n706_adj_2044 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16990 ),
            .carryout(\foc.u_Park_Transform.n16991 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_16_lut_LC_13_16_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_16_lut_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_567_16_lut_LC_13_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_567_16_lut_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__35941),
            .in2(N__35920),
            .in3(N__35899),
            .lcout(\foc.u_Park_Transform.n762_adj_2065 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n16991 ),
            .carryout(\foc.u_Park_Transform.n763_adj_2054 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n763_adj_2054_THRU_LUT4_0_LC_13_16_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n763_adj_2054_THRU_LUT4_0_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n763_adj_2054_THRU_LUT4_0_LC_13_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n763_adj_2054_THRU_LUT4_0_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36490),
            .lcout(\foc.u_Park_Transform.n763_adj_2054_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_2_lut_LC_13_17_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_2_lut_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_2_lut_LC_13_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_2_lut_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__36472),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2411 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_3_lut_LC_13_17_1 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_3_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_3_lut_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_3_lut_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__36661),
            .in2(N__36400),
            .in3(N__36379),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2511 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17367 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_4_lut_LC_13_17_2 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_4_lut_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_4_lut_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__36376),
            .in2(N__36678),
            .in3(N__36349),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2611 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17368 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_5_lut_LC_13_17_3 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_5_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_5_lut_LC_13_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_5_lut_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__36665),
            .in2(N__36346),
            .in3(N__36322),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2711 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17369 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_6_lut_LC_13_17_4 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_6_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_6_lut_LC_13_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_6_lut_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__36319),
            .in2(N__36679),
            .in3(N__36298),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2811 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17370 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_7_lut_LC_13_17_5 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_7_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_7_lut_LC_13_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_7_lut_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__36295),
            .in2(N__36681),
            .in3(N__36277),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n2911 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17371 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_8_lut_LC_13_17_6 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_8_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_8_lut_LC_13_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_8_lut_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__36274),
            .in2(N__36680),
            .in3(N__36253),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3011 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17372 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_9_lut_LC_13_17_7 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_9_lut_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_9_lut_LC_13_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_9_lut_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__36691),
            .in2(N__36682),
            .in3(N__36610),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3111 ),
            .ltout(),
            .carryin(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17373 ),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n17374 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_10_lut_LC_13_18_0 .C_ON=1'b1;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_10_lut_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_10_lut_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.add_5956_10_lut_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__36607),
            .in2(_gnd_net_),
            .in3(N__36589),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3215 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_LUT4_0_LC_13_18_1 .C_ON=1'b0;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_LUT4_0_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_LUT4_0_LC_13_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_LUT4_0_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36586),
            .lcout(\foc.u_Sine_Cosine.u_Sine_Cosine_LUT.n3216_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i1_1_lut_2_lut_LC_13_18_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i1_1_lut_2_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i1_1_lut_2_lut_LC_13_18_2 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i1_1_lut_2_lut_LC_13_18_2  (
            .in0(N__36561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_13_18_7.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_13_18_7.LUT_INIT=16'b1000100011111000;
    LogicCell40 i1_3_lut_4_lut_LC_13_18_7 (
            .in0(N__44894),
            .in1(N__40458),
            .in2(_gnd_net_),
            .in3(N__40497),
            .lcout(n794),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_13_20_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_13_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__66056),
            .in2(N__66217),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n81_adj_750 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17856 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_13_20_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_13_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__66180),
            .in2(N__38416),
            .in3(N__36505),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n130_adj_748 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17856 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17857 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_13_20_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_13_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__38407),
            .in2(N__66218),
            .in3(N__36493),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n179_adj_746 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17857 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17858 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_13_20_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_13_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__66184),
            .in2(N__38398),
            .in3(N__36790),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n228_adj_742 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17858 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17859 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_13_20_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_13_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__38386),
            .in2(N__66219),
            .in3(N__36775),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n277_adj_741 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17859 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17860 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_13_20_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_13_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__66188),
            .in2(N__38536),
            .in3(N__36763),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n326 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17860 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17861 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_13_20_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_13_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__38524),
            .in2(N__66220),
            .in3(N__36748),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n375 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17861 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17862 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_13_20_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_13_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__66192),
            .in2(N__38515),
            .in3(N__36736),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n424 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17862 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17863 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_13_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_13_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__38495),
            .in2(N__66293),
            .in3(N__36724),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n473 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17864 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_13_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_13_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__66259),
            .in2(N__38502),
            .in3(N__36700),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n522 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17864 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17865 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_13_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_13_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__45426),
            .in2(N__38503),
            .in3(N__36697),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n778_adj_737 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17865 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_LUT4_0_LC_13_21_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_LUT4_0_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_LUT4_0_LC_13_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_LUT4_0_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36694),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_adj_736_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_1_LC_13_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_1_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_1_LC_13_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_1_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__43245),
            .in2(N__43249),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17957 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_2_lut_LC_13_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_2_lut_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_2_lut_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_2_lut_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__48968),
            .in2(_gnd_net_),
            .in3(N__36826),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17957 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17958 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_3_lut_LC_13_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_3_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_3_lut_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_3_lut_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__43759),
            .in2(N__43222),
            .in3(N__36823),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17958 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17959 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_4_lut_LC_13_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_4_lut_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_4_lut_LC_13_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_4_lut_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__43510),
            .in2(N__43741),
            .in3(N__36820),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17959 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17960 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_5_lut_LC_13_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_5_lut_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_5_lut_LC_13_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_5_lut_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__38794),
            .in2(N__43489),
            .in3(N__36817),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17960 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17961 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_6_lut_LC_13_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_6_lut_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_6_lut_LC_13_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_6_lut_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__38629),
            .in2(N__38776),
            .in3(N__36814),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17961 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17962 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_7_lut_LC_13_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_7_lut_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_7_lut_LC_13_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_7_lut_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__41017),
            .in2(N__38614),
            .in3(N__36811),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17962 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17963 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_8_lut_LC_13_22_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_8_lut_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_8_lut_LC_13_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_8_lut_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__41284),
            .in2(N__40999),
            .in3(N__36808),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17963 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17964 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_9_lut_LC_13_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_9_lut_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_9_lut_LC_13_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_9_lut_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__37009),
            .in2(N__41266),
            .in3(N__36805),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_22 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17965 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_10_lut_LC_13_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_10_lut_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_10_lut_LC_13_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_10_lut_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__36994),
            .in2(N__36910),
            .in3(N__36898),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_23 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17965 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17966 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_11_lut_LC_13_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_11_lut_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_11_lut_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_11_lut_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__36895),
            .in2(N__36889),
            .in3(N__36877),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17966 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17967 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_12_lut_LC_13_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_12_lut_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_12_lut_LC_13_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_12_lut_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__36874),
            .in2(N__36865),
            .in3(N__36856),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17967 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17968 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_13_lut_LC_13_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_13_lut_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_13_lut_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_13_lut_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__38479),
            .in2(N__36853),
            .in3(N__36841),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17968 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17969 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_14_lut_LC_13_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_14_lut_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_14_lut_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_14_lut_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__40651),
            .in2(N__38467),
            .in3(N__36838),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17969 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17970 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_15_lut_LC_13_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_15_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_15_lut_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_15_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__40633),
            .in2(N__40789),
            .in3(N__36835),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17970 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17971 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_16_lut_LC_13_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_16_lut_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_16_lut_LC_13_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_16_lut_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__40774),
            .in2(N__40819),
            .in3(N__36832),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17971 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17972 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_17_lut_LC_13_24_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_17_lut_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_17_lut_LC_13_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4258_17_lut_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__49011),
            .in2(_gnd_net_),
            .in3(N__36829),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_13_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_13_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__66822),
            .in2(N__63111),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n72_adj_634 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_13_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_13_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__36985),
            .in2(N__63132),
            .in3(N__36979),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n121_adj_633 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18092 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_13_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_13_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__36976),
            .in2(N__63112),
            .in3(N__36970),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n170_adj_632 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18093 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_13_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_13_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(N__36967),
            .in2(N__63133),
            .in3(N__36961),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n219_adj_631 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18094 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_13_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_13_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__36958),
            .in2(N__63113),
            .in3(N__36952),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n268_adj_630 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18095 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_13_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_13_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__36949),
            .in2(N__63134),
            .in3(N__36943),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n317_adj_629 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18096 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_13_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_13_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__36940),
            .in2(N__63114),
            .in3(N__36934),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n366_adj_628 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18097 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_13_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_13_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(N__36931),
            .in2(N__63135),
            .in3(N__36925),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n415_adj_627 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18098 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_13_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__36922),
            .in2(N__63096),
            .in3(N__36913),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n464_adj_626 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_13_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__63044),
            .in2(N__37072),
            .in3(N__37063),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n513_adj_625 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18100 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_13_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__37060),
            .in2(N__63097),
            .in3(N__37054),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n562_adj_624 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18101 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_13_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__63048),
            .in2(N__37051),
            .in3(N__37042),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n611_adj_623 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18102 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_13_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__37039),
            .in2(N__63098),
            .in3(N__37033),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n660_adj_622 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18103 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_13_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__63052),
            .in2(N__37030),
            .in3(N__37021),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n709_adj_621 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18104 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_13_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__45169),
            .in2(N__37018),
            .in3(N__37000),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n766_adj_619 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18105 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_LUT4_0_LC_13_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_LUT4_0_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_LUT4_0_LC_13_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_LUT4_0_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36997),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_adj_620_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i9_1_lut_LC_14_5_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i9_1_lut_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i9_1_lut_LC_14_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i9_1_lut_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37084),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i19_1_lut_LC_14_5_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i19_1_lut_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i19_1_lut_LC_14_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i19_1_lut_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37336),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15_adj_518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i6_1_lut_LC_14_5_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i6_1_lut_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i6_1_lut_LC_14_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i6_1_lut_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37120),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i26_1_lut_LC_14_5_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i26_1_lut_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i26_1_lut_LC_14_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i26_1_lut_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37429),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i5_1_lut_LC_14_5_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i5_1_lut_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i5_1_lut_LC_14_5_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i5_1_lut_LC_14_5_4  (
            .in0(N__37129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i8_1_lut_LC_14_5_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i8_1_lut_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i8_1_lut_LC_14_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i8_1_lut_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37096),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i4_1_lut_LC_14_5_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i4_1_lut_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i4_1_lut_LC_14_5_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i4_1_lut_LC_14_5_6  (
            .in0(N__39151),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i7_1_lut_LC_14_5_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i7_1_lut_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i7_1_lut_LC_14_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i7_1_lut_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37108),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i17_1_lut_LC_14_6_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i17_1_lut_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i17_1_lut_LC_14_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i17_1_lut_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37141),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i14_1_lut_LC_14_6_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i14_1_lut_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i14_1_lut_LC_14_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i14_1_lut_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37177),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i11_1_lut_LC_14_6_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i11_1_lut_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i11_1_lut_LC_14_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i11_1_lut_LC_14_6_2  (
            .in0(N__37207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i16_1_lut_LC_14_6_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i16_1_lut_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i16_1_lut_LC_14_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i16_1_lut_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37153),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i10_1_lut_LC_14_6_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i10_1_lut_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i10_1_lut_LC_14_6_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i10_1_lut_LC_14_6_4  (
            .in0(N__37216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i13_1_lut_LC_14_6_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i13_1_lut_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i13_1_lut_LC_14_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i13_1_lut_LC_14_6_5  (
            .in0(N__37189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i15_1_lut_LC_14_6_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i15_1_lut_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i15_1_lut_LC_14_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i15_1_lut_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37165),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i12_1_lut_LC_14_6_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i12_1_lut_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i12_1_lut_LC_14_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i12_1_lut_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37198),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_2_lut_LC_14_7_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_2_lut_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_2_lut_LC_14_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_2_lut_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__39139),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.dCurrent_4 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\foc.u_Park_Transform.n17277 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_3_lut_LC_14_7_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_3_lut_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_3_lut_LC_14_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_3_lut_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__39127),
            .in2(_gnd_net_),
            .in3(N__37111),
            .lcout(\foc.dCurrent_5 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17277 ),
            .carryout(\foc.u_Park_Transform.n17278 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_4_lut_LC_14_7_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_4_lut_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_4_lut_LC_14_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_4_lut_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__39115),
            .in2(_gnd_net_),
            .in3(N__37099),
            .lcout(\foc.dCurrent_6 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17278 ),
            .carryout(\foc.u_Park_Transform.n17279 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_5_lut_LC_14_7_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_5_lut_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_5_lut_LC_14_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_5_lut_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__39103),
            .in2(_gnd_net_),
            .in3(N__37087),
            .lcout(\foc.dCurrent_7 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17279 ),
            .carryout(\foc.u_Park_Transform.n17280 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_6_lut_LC_14_7_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_6_lut_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_6_lut_LC_14_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_6_lut_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__39091),
            .in2(_gnd_net_),
            .in3(N__37075),
            .lcout(\foc.dCurrent_8 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17280 ),
            .carryout(\foc.u_Park_Transform.n17281 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_7_lut_LC_14_7_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_7_lut_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_7_lut_LC_14_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_7_lut_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__39484),
            .in2(_gnd_net_),
            .in3(N__37210),
            .lcout(\foc.dCurrent_9 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17281 ),
            .carryout(\foc.u_Park_Transform.n17282 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_8_lut_LC_14_7_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_8_lut_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_8_lut_LC_14_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_8_lut_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__39472),
            .in2(_gnd_net_),
            .in3(N__37201),
            .lcout(\foc.dCurrent_10 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17282 ),
            .carryout(\foc.u_Park_Transform.n17283 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_9_lut_LC_14_7_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_9_lut_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_9_lut_LC_14_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_9_lut_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__39457),
            .in2(_gnd_net_),
            .in3(N__37192),
            .lcout(\foc.dCurrent_11 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17283 ),
            .carryout(\foc.u_Park_Transform.n17284 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_10_lut_LC_14_8_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_10_lut_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_10_lut_LC_14_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_10_lut_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__39442),
            .in2(_gnd_net_),
            .in3(N__37180),
            .lcout(\foc.dCurrent_12 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\foc.u_Park_Transform.n17285 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_11_lut_LC_14_8_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_11_lut_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_11_lut_LC_14_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_11_lut_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__39427),
            .in2(_gnd_net_),
            .in3(N__37168),
            .lcout(\foc.dCurrent_13 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17285 ),
            .carryout(\foc.u_Park_Transform.n17286 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_12_lut_LC_14_8_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_12_lut_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_12_lut_LC_14_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_12_lut_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__39415),
            .in2(_gnd_net_),
            .in3(N__37156),
            .lcout(\foc.dCurrent_14 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17286 ),
            .carryout(\foc.u_Park_Transform.n17287 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_13_lut_LC_14_8_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_13_lut_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_13_lut_LC_14_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_13_lut_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__39403),
            .in2(_gnd_net_),
            .in3(N__37144),
            .lcout(\foc.dCurrent_15 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17287 ),
            .carryout(\foc.u_Park_Transform.n17288 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_14_lut_LC_14_8_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_14_lut_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_14_lut_LC_14_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_14_lut_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__39211),
            .in2(_gnd_net_),
            .in3(N__37132),
            .lcout(\foc.dCurrent_16 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17288 ),
            .carryout(\foc.u_Park_Transform.n17289 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_15_lut_LC_14_8_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_15_lut_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_15_lut_LC_14_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_15_lut_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__37360),
            .in2(_gnd_net_),
            .in3(N__37345),
            .lcout(\foc.dCurrent_17 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17289 ),
            .carryout(\foc.u_Park_Transform.n17290 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_16_lut_LC_14_8_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_16_lut_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_16_lut_LC_14_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_16_lut_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__37342),
            .in2(_gnd_net_),
            .in3(N__37327),
            .lcout(\foc.dCurrent_18 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17290 ),
            .carryout(\foc.u_Park_Transform.n17291 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_17_lut_LC_14_8_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_17_lut_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_17_lut_LC_14_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_17_lut_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__37324),
            .in2(_gnd_net_),
            .in3(N__37309),
            .lcout(\foc.dCurrent_19 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17291 ),
            .carryout(\foc.u_Park_Transform.n17292 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_18_lut_LC_14_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_18_lut_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_18_lut_LC_14_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_18_lut_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__37306),
            .in2(_gnd_net_),
            .in3(N__37291),
            .lcout(\foc.dCurrent_20 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\foc.u_Park_Transform.n17293 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_19_lut_LC_14_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_19_lut_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_19_lut_LC_14_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_19_lut_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__37288),
            .in2(_gnd_net_),
            .in3(N__37273),
            .lcout(\foc.dCurrent_21 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17293 ),
            .carryout(\foc.u_Park_Transform.n17294 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_20_lut_LC_14_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_20_lut_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_20_lut_LC_14_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_20_lut_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__37270),
            .in2(_gnd_net_),
            .in3(N__37255),
            .lcout(\foc.dCurrent_22 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17294 ),
            .carryout(\foc.u_Park_Transform.n17295 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_21_lut_LC_14_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_21_lut_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_21_lut_LC_14_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_21_lut_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__37252),
            .in2(_gnd_net_),
            .in3(N__37237),
            .lcout(\foc.dCurrent_23 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17295 ),
            .carryout(\foc.u_Park_Transform.n17296 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_22_lut_LC_14_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_22_lut_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_22_lut_LC_14_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_22_lut_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__37234),
            .in2(_gnd_net_),
            .in3(N__37219),
            .lcout(\foc.dCurrent_24 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17296 ),
            .carryout(\foc.u_Park_Transform.n17297 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_23_lut_LC_14_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_23_lut_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_23_lut_LC_14_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_23_lut_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__37435),
            .in2(_gnd_net_),
            .in3(N__37420),
            .lcout(\foc.dCurrent_25 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17297 ),
            .carryout(\foc.u_Park_Transform.n17298 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_24_lut_LC_14_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_24_lut_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_24_lut_LC_14_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_24_lut_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__37417),
            .in2(_gnd_net_),
            .in3(N__37411),
            .lcout(\foc.dCurrent_26 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17298 ),
            .carryout(\foc.u_Park_Transform.n17299 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_25_lut_LC_14_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_25_lut_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_25_lut_LC_14_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_25_lut_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__37408),
            .in2(_gnd_net_),
            .in3(N__37402),
            .lcout(\foc.dCurrent_27 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17299 ),
            .carryout(\foc.u_Park_Transform.n17300 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_26_lut_LC_14_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_26_lut_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_26_lut_LC_14_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_26_lut_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__37399),
            .in2(_gnd_net_),
            .in3(N__37393),
            .lcout(\foc.dCurrent_28 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\foc.u_Park_Transform.n17301 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_27_lut_LC_14_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_27_lut_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_27_lut_LC_14_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_27_lut_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__37390),
            .in2(_gnd_net_),
            .in3(N__37384),
            .lcout(\foc.dCurrent_29 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17301 ),
            .carryout(\foc.u_Park_Transform.n17302 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_28_lut_LC_14_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.add_8094_28_lut_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_28_lut_LC_14_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_28_lut_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__37381),
            .in2(_gnd_net_),
            .in3(N__37375),
            .lcout(\foc.dCurrent_30 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17302 ),
            .carryout(\foc.u_Park_Transform.n17303 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.add_8094_29_lut_LC_14_10_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.add_8094_29_lut_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.add_8094_29_lut_LC_14_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.add_8094_29_lut_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__37372),
            .in2(_gnd_net_),
            .in3(N__37366),
            .lcout(),
            .ltout(\foc.dCurrent_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i32_1_lut_LC_14_10_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i32_1_lut_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i32_1_lut_LC_14_10_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i32_1_lut_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37363),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i30_1_lut_LC_14_10_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i30_1_lut_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i30_1_lut_LC_14_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i30_1_lut_LC_14_10_5  (
            .in0(N__37468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n4_adj_515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i29_1_lut_LC_14_10_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i29_1_lut_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i29_1_lut_LC_14_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i29_1_lut_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37462),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i31_1_lut_LC_14_10_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i31_1_lut_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i31_1_lut_LC_14_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i31_1_lut_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37456),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_2_lut_LC_14_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_2_lut_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_2_lut_LC_14_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_2_lut_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__42182),
            .in2(N__42700),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n57_adj_2116 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\foc.u_Park_Transform.n17221 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_3_lut_LC_14_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_3_lut_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_3_lut_LC_14_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_3_lut_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__42683),
            .in2(N__41542),
            .in3(N__37450),
            .lcout(\foc.u_Park_Transform.n106_adj_2115 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17221 ),
            .carryout(\foc.u_Park_Transform.n17222 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_4_lut_LC_14_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_4_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_4_lut_LC_14_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_4_lut_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__42684),
            .in2(N__41521),
            .in3(N__37447),
            .lcout(\foc.u_Park_Transform.n155_adj_2114 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17222 ),
            .carryout(\foc.u_Park_Transform.n17223 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_5_lut_LC_14_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_5_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_5_lut_LC_14_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_5_lut_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__41494),
            .in2(N__42701),
            .in3(N__37444),
            .lcout(\foc.u_Park_Transform.n204_adj_2113 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17223 ),
            .carryout(\foc.u_Park_Transform.n17224 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_6_lut_LC_14_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_6_lut_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_6_lut_LC_14_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_6_lut_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__42688),
            .in2(N__41473),
            .in3(N__37441),
            .lcout(\foc.u_Park_Transform.n253_adj_2112 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17224 ),
            .carryout(\foc.u_Park_Transform.n17225 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_7_lut_LC_14_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_7_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_7_lut_LC_14_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_7_lut_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__41446),
            .in2(N__42702),
            .in3(N__37438),
            .lcout(\foc.u_Park_Transform.n302_adj_2111 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17225 ),
            .carryout(\foc.u_Park_Transform.n17226 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_8_lut_LC_14_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_8_lut_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_8_lut_LC_14_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_8_lut_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__42692),
            .in2(N__41422),
            .in3(N__37507),
            .lcout(\foc.u_Park_Transform.n351_adj_2108 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17226 ),
            .carryout(\foc.u_Park_Transform.n17227 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_9_lut_LC_14_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_9_lut_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_9_lut_LC_14_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_9_lut_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__41917),
            .in2(N__42703),
            .in3(N__37504),
            .lcout(\foc.u_Park_Transform.n400_adj_2106 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17227 ),
            .carryout(\foc.u_Park_Transform.n17228 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_10_lut_LC_14_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_10_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_10_lut_LC_14_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_10_lut_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__42666),
            .in2(N__41896),
            .in3(N__37501),
            .lcout(\foc.u_Park_Transform.n449_adj_2103 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\foc.u_Park_Transform.n17229 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_11_lut_LC_14_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_11_lut_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_11_lut_LC_14_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_11_lut_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__41863),
            .in2(N__42696),
            .in3(N__37498),
            .lcout(\foc.u_Park_Transform.n498_adj_2102 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17229 ),
            .carryout(\foc.u_Park_Transform.n17230 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_12_lut_LC_14_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_12_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_12_lut_LC_14_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_12_lut_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__42670),
            .in2(N__41842),
            .in3(N__37495),
            .lcout(\foc.u_Park_Transform.n547_adj_2100 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17230 ),
            .carryout(\foc.u_Park_Transform.n17231 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_13_lut_LC_14_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_13_lut_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_13_lut_LC_14_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_13_lut_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__41815),
            .in2(N__42697),
            .in3(N__37492),
            .lcout(\foc.u_Park_Transform.n596_adj_2099 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17231 ),
            .carryout(\foc.u_Park_Transform.n17232 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_14_lut_LC_14_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_14_lut_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_14_lut_LC_14_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_14_lut_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__41791),
            .in2(N__42699),
            .in3(N__37489),
            .lcout(\foc.u_Park_Transform.n645_adj_2098 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17232 ),
            .carryout(\foc.u_Park_Transform.n17233 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_15_lut_LC_14_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_15_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_15_lut_LC_14_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_15_lut_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__41770),
            .in2(N__42698),
            .in3(N__37486),
            .lcout(\foc.u_Park_Transform.n694_adj_2097 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17233 ),
            .carryout(\foc.u_Park_Transform.n17234 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_16_lut_LC_14_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_16_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_16_lut_LC_14_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_563_16_lut_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__42789),
            .in2(N__41749),
            .in3(N__37471),
            .lcout(\foc.u_Park_Transform.n746 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17234 ),
            .carryout(\foc.u_Park_Transform.n747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n747_THRU_LUT4_0_LC_14_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n747_THRU_LUT4_0_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n747_THRU_LUT4_0_LC_14_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n747_THRU_LUT4_0_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37780),
            .lcout(\foc.u_Park_Transform.n747_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_2_lut_LC_14_13_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_2_lut_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_2_lut_LC_14_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_2_lut_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__37749),
            .in2(N__41685),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n63 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\foc.u_Park_Transform.n17008 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_3_lut_LC_14_13_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_3_lut_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_3_lut_LC_14_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_3_lut_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__41638),
            .in2(N__37582),
            .in3(N__37573),
            .lcout(\foc.u_Park_Transform.n112 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17008 ),
            .carryout(\foc.u_Park_Transform.n17009 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_4_lut_LC_14_13_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_4_lut_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_4_lut_LC_14_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_4_lut_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__41639),
            .in2(N__37570),
            .in3(N__37561),
            .lcout(\foc.u_Park_Transform.n161 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17009 ),
            .carryout(\foc.u_Park_Transform.n17010 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_5_lut_LC_14_13_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_5_lut_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_5_lut_LC_14_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_5_lut_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__37558),
            .in2(N__41686),
            .in3(N__37552),
            .lcout(\foc.u_Park_Transform.n210 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17010 ),
            .carryout(\foc.u_Park_Transform.n17011 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_6_lut_LC_14_13_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_6_lut_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_6_lut_LC_14_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_6_lut_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__41643),
            .in2(N__37549),
            .in3(N__37540),
            .lcout(\foc.u_Park_Transform.n259 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17011 ),
            .carryout(\foc.u_Park_Transform.n17012 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_7_lut_LC_14_13_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_7_lut_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_7_lut_LC_14_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_7_lut_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__37537),
            .in2(N__41687),
            .in3(N__37531),
            .lcout(\foc.u_Park_Transform.n308 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17012 ),
            .carryout(\foc.u_Park_Transform.n17013 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_8_lut_LC_14_13_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_8_lut_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_8_lut_LC_14_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_8_lut_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__41647),
            .in2(N__37528),
            .in3(N__37519),
            .lcout(\foc.u_Park_Transform.n357 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17013 ),
            .carryout(\foc.u_Park_Transform.n17014 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_9_lut_LC_14_13_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_9_lut_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_9_lut_LC_14_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_9_lut_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__37516),
            .in2(N__41688),
            .in3(N__37510),
            .lcout(\foc.u_Park_Transform.n406 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17014 ),
            .carryout(\foc.u_Park_Transform.n17015 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_10_lut_LC_14_14_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_10_lut_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_10_lut_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_10_lut_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__41692),
            .in2(N__37903),
            .in3(N__37894),
            .lcout(\foc.u_Park_Transform.n455 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\foc.u_Park_Transform.n17016 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_11_lut_LC_14_14_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_11_lut_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_11_lut_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_11_lut_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__37891),
            .in2(N__41707),
            .in3(N__37885),
            .lcout(\foc.u_Park_Transform.n504 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17016 ),
            .carryout(\foc.u_Park_Transform.n17017 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_12_lut_LC_14_14_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_12_lut_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_12_lut_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_12_lut_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__41696),
            .in2(N__37882),
            .in3(N__37873),
            .lcout(\foc.u_Park_Transform.n553 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17017 ),
            .carryout(\foc.u_Park_Transform.n17018 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_13_lut_LC_14_14_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_13_lut_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_13_lut_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_13_lut_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__37870),
            .in2(N__41708),
            .in3(N__37864),
            .lcout(\foc.u_Park_Transform.n602 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17018 ),
            .carryout(\foc.u_Park_Transform.n17019 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_14_lut_LC_14_14_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_14_lut_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_14_lut_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_14_lut_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__41700),
            .in2(N__37861),
            .in3(N__37852),
            .lcout(\foc.u_Park_Transform.n651 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17019 ),
            .carryout(\foc.u_Park_Transform.n17020 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_15_lut_LC_14_14_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_15_lut_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_15_lut_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_15_lut_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__37849),
            .in2(N__41709),
            .in3(N__37843),
            .lcout(\foc.u_Park_Transform.n700 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17020 ),
            .carryout(\foc.u_Park_Transform.n17021 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_16_lut_LC_14_14_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_16_lut_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_565_16_lut_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_565_16_lut_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__37840),
            .in2(N__37822),
            .in3(N__37801),
            .lcout(\foc.u_Park_Transform.n754 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17021 ),
            .carryout(\foc.u_Park_Transform.n755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n755_THRU_LUT4_0_LC_14_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n755_THRU_LUT4_0_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n755_THRU_LUT4_0_LC_14_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n755_THRU_LUT4_0_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37798),
            .lcout(\foc.u_Park_Transform.n755_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_2_lut_LC_14_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_2_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_2_lut_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_2_lut_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__40313),
            .in2(N__39313),
            .in3(_gnd_net_),
            .lcout(\foc.qCurrent_3 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\foc.u_Park_Transform.n17068 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_3_lut_LC_14_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_3_lut_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_3_lut_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_3_lut_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__39274),
            .in2(N__40090),
            .in3(N__37927),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_2 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17068 ),
            .carryout(\foc.u_Park_Transform.n17069 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_4_lut_LC_14_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_4_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_4_lut_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_4_lut_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__40081),
            .in2(N__39314),
            .in3(N__37924),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_3 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17069 ),
            .carryout(\foc.u_Park_Transform.n17070 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_5_lut_LC_14_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_5_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_5_lut_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_5_lut_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__39278),
            .in2(N__40072),
            .in3(N__37921),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_4 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17070 ),
            .carryout(\foc.u_Park_Transform.n17071 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_6_lut_LC_14_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_6_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_6_lut_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_6_lut_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__40060),
            .in2(N__39315),
            .in3(N__37918),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_5 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17071 ),
            .carryout(\foc.u_Park_Transform.n17072 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_7_lut_LC_14_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_7_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_7_lut_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_7_lut_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__39282),
            .in2(N__40051),
            .in3(N__37915),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_6 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17072 ),
            .carryout(\foc.u_Park_Transform.n17073 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_8_lut_LC_14_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_8_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_8_lut_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_8_lut_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__40039),
            .in2(N__39316),
            .in3(N__37912),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_7 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17073 ),
            .carryout(\foc.u_Park_Transform.n17074 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_9_lut_LC_14_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_9_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_9_lut_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_9_lut_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__39286),
            .in2(N__40030),
            .in3(N__37909),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_8 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17074 ),
            .carryout(\foc.u_Park_Transform.n17075 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_10_lut_LC_14_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_10_lut_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_10_lut_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_10_lut_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__40018),
            .in2(N__39348),
            .in3(N__37906),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_9 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\foc.u_Park_Transform.n17076 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_11_lut_LC_14_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_11_lut_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_11_lut_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_11_lut_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__40198),
            .in2(N__39351),
            .in3(N__38008),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_10 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17076 ),
            .carryout(\foc.u_Park_Transform.n17077 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_12_lut_LC_14_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_12_lut_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_12_lut_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_12_lut_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__40189),
            .in2(N__39349),
            .in3(N__38005),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_11 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17077 ),
            .carryout(\foc.u_Park_Transform.n17078 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_13_lut_LC_14_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_13_lut_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_13_lut_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_13_lut_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__40180),
            .in2(N__39352),
            .in3(N__38002),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_12 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17078 ),
            .carryout(\foc.u_Park_Transform.n17079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_14_lut_LC_14_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_14_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_14_lut_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_14_lut_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__40171),
            .in2(N__39350),
            .in3(N__37999),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_13 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17079 ),
            .carryout(\foc.u_Park_Transform.n17080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_15_lut_LC_14_16_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_15_lut_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_15_lut_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_15_lut_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__40162),
            .in2(N__39353),
            .in3(N__37996),
            .lcout(\foc.u_Park_Transform.Product4_mul_temp_14 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17080 ),
            .carryout(\foc.u_Park_Transform.n17081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_16_lut_LC_14_16_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_16_lut_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_561_16_lut_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_561_16_lut_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__39195),
            .in2(N__40153),
            .in3(N__37972),
            .lcout(\foc.u_Park_Transform.n738_adj_2003 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17081 ),
            .carryout(\foc.u_Park_Transform.n739_adj_2006 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n739_adj_2006_THRU_LUT4_0_LC_14_16_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n739_adj_2006_THRU_LUT4_0_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n739_adj_2006_THRU_LUT4_0_LC_14_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n739_adj_2006_THRU_LUT4_0_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37969),
            .lcout(\foc.u_Park_Transform.n739_adj_2006_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_2_lut_LC_14_17_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_2_lut_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_2_lut_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_2_lut_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__37951),
            .in2(N__44893),
            .in3(N__37942),
            .lcout(\foc.qCurrent_4 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\foc.u_Park_Transform.n15748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_3_lut_LC_14_17_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_3_lut_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_3_lut_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_3_lut_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__37939),
            .in2(N__68390),
            .in3(N__37930),
            .lcout(\foc.qCurrent_5 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15748 ),
            .carryout(\foc.u_Park_Transform.n15749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_4_lut_LC_14_17_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_4_lut_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_4_lut_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_4_lut_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__38107),
            .in2(N__68393),
            .in3(N__38098),
            .lcout(\foc.qCurrent_6 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15749 ),
            .carryout(\foc.u_Park_Transform.n15750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_5_lut_LC_14_17_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_5_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_5_lut_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_5_lut_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__38095),
            .in2(N__68391),
            .in3(N__38086),
            .lcout(\foc.qCurrent_7 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15750 ),
            .carryout(\foc.u_Park_Transform.n15751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_6_lut_LC_14_17_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_6_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_6_lut_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_6_lut_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__38083),
            .in2(N__68394),
            .in3(N__38074),
            .lcout(\foc.qCurrent_8 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15751 ),
            .carryout(\foc.u_Park_Transform.n15752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_7_lut_LC_14_17_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_7_lut_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_7_lut_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_7_lut_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__38071),
            .in2(N__68392),
            .in3(N__38062),
            .lcout(\foc.qCurrent_9 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15752 ),
            .carryout(\foc.u_Park_Transform.n15753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_8_lut_LC_14_17_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_8_lut_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_8_lut_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_8_lut_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__38059),
            .in2(N__68395),
            .in3(N__38050),
            .lcout(\foc.qCurrent_10 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15753 ),
            .carryout(\foc.u_Park_Transform.n15754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_9_lut_LC_14_17_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_9_lut_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_9_lut_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_9_lut_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__68332),
            .in2(N__38047),
            .in3(N__38038),
            .lcout(\foc.qCurrent_11 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15754 ),
            .carryout(\foc.u_Park_Transform.n15755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_10_lut_LC_14_18_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_10_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_10_lut_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_10_lut_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__38035),
            .in2(N__68396),
            .in3(N__38026),
            .lcout(\foc.qCurrent_12 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\foc.u_Park_Transform.n15756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_11_lut_LC_14_18_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_11_lut_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_11_lut_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_11_lut_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__68336),
            .in2(N__38023),
            .in3(N__38011),
            .lcout(\foc.qCurrent_13 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15756 ),
            .carryout(\foc.u_Park_Transform.n15757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_12_lut_LC_14_18_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_12_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_12_lut_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_12_lut_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__38245),
            .in2(N__68397),
            .in3(N__38236),
            .lcout(\foc.qCurrent_14 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15757 ),
            .carryout(\foc.u_Park_Transform.n15758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_13_lut_LC_14_18_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_13_lut_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_13_lut_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_13_lut_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__68340),
            .in2(N__38233),
            .in3(N__38221),
            .lcout(\foc.qCurrent_15 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15758 ),
            .carryout(\foc.u_Park_Transform.n15759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_14_lut_LC_14_18_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_14_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_14_lut_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_14_lut_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(N__68398),
            .in3(N__38209),
            .lcout(\foc.qCurrent_16 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15759 ),
            .carryout(\foc.u_Park_Transform.n15760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_15_lut_LC_14_18_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_15_lut_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_15_lut_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_15_lut_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__68344),
            .in2(N__38206),
            .in3(N__38191),
            .lcout(\foc.qCurrent_17 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15760 ),
            .carryout(\foc.u_Park_Transform.n15761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_16_lut_LC_14_18_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_16_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_16_lut_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_16_lut_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__38188),
            .in2(N__68399),
            .in3(N__38176),
            .lcout(\foc.qCurrent_18 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15761 ),
            .carryout(\foc.u_Park_Transform.n15762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_17_lut_LC_14_18_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_17_lut_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_17_lut_LC_14_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_17_lut_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__68348),
            .in2(N__38173),
            .in3(N__38158),
            .lcout(\foc.qCurrent_19 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15762 ),
            .carryout(\foc.u_Park_Transform.n15763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_18_lut_LC_14_19_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_18_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_18_lut_LC_14_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_18_lut_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__38155),
            .in2(N__68400),
            .in3(N__38143),
            .lcout(\foc.qCurrent_20 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\foc.u_Park_Transform.n15764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_19_lut_LC_14_19_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_19_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_19_lut_LC_14_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_19_lut_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__68352),
            .in2(N__38140),
            .in3(N__38125),
            .lcout(\foc.qCurrent_21 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15764 ),
            .carryout(\foc.u_Park_Transform.n15765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_20_lut_LC_14_19_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_20_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_20_lut_LC_14_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_20_lut_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__38122),
            .in2(N__68401),
            .in3(N__38110),
            .lcout(\foc.qCurrent_22 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15765 ),
            .carryout(\foc.u_Park_Transform.n15766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_21_lut_LC_14_19_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_21_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_21_lut_LC_14_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_21_lut_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__68356),
            .in2(N__38377),
            .in3(N__38362),
            .lcout(\foc.qCurrent_23 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15766 ),
            .carryout(\foc.u_Park_Transform.n15767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_22_lut_LC_14_19_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_22_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_22_lut_LC_14_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_22_lut_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__38359),
            .in2(N__68402),
            .in3(N__38347),
            .lcout(\foc.qCurrent_24 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15767 ),
            .carryout(\foc.u_Park_Transform.n15768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_23_lut_LC_14_19_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_23_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_23_lut_LC_14_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_23_lut_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__68360),
            .in2(N__38344),
            .in3(N__38329),
            .lcout(\foc.qCurrent_25 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15768 ),
            .carryout(\foc.u_Park_Transform.n15769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_24_lut_LC_14_19_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_24_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_24_lut_LC_14_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_24_lut_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__38326),
            .in2(N__68403),
            .in3(N__38314),
            .lcout(\foc.qCurrent_26 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15769 ),
            .carryout(\foc.u_Park_Transform.n15770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_25_lut_LC_14_19_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_25_lut_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_25_lut_LC_14_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_25_lut_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__68364),
            .in2(N__38311),
            .in3(N__38296),
            .lcout(\foc.qCurrent_27 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15770 ),
            .carryout(\foc.u_Park_Transform.n15771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_26_lut_LC_14_20_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_26_lut_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_26_lut_LC_14_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_26_lut_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__38293),
            .in2(N__68426),
            .in3(N__38281),
            .lcout(\foc.qCurrent_28 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\foc.u_Park_Transform.n15772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_27_lut_LC_14_20_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_27_lut_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_27_lut_LC_14_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_27_lut_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__68407),
            .in2(N__38278),
            .in3(N__38263),
            .lcout(\foc.qCurrent_29 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15772 ),
            .carryout(\foc.u_Park_Transform.n15773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_28_lut_LC_14_20_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.sub_65_add_2_28_lut_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_28_lut_LC_14_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_28_lut_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__38260),
            .in2(N__68427),
            .in3(N__38248),
            .lcout(\foc.qCurrent_30 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n15773 ),
            .carryout(\foc.u_Park_Transform.n15774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.sub_65_add_2_29_lut_LC_14_20_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.sub_65_add_2_29_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.sub_65_add_2_29_lut_LC_14_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_Park_Transform.sub_65_add_2_29_lut_LC_14_20_3  (
            .in0(N__38455),
            .in1(N__68411),
            .in2(_gnd_net_),
            .in3(N__38443),
            .lcout(\foc.qCurrent_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i20_1_lut_LC_14_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i20_1_lut_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i20_1_lut_LC_14_20_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i20_1_lut_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__38440),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i28_1_lut_LC_14_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i28_1_lut_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i28_1_lut_LC_14_20_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i28_1_lut_LC_14_20_5  (
            .in0(N__38434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i22_1_lut_LC_14_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i22_1_lut_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i22_1_lut_LC_14_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i22_1_lut_LC_14_20_6  (
            .in0(N__38428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i29_1_lut_LC_14_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i29_1_lut_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i29_1_lut_LC_14_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i29_1_lut_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38422),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_14_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_14_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__65739),
            .in2(N__66028),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n84_adj_749 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_14_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__40723),
            .in2(N__66031),
            .in3(N__38401),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n133_adj_747 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17727 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_14_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__40717),
            .in2(N__66029),
            .in3(N__38389),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n182_adj_745 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17728 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_14_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__65975),
            .in2(N__40708),
            .in3(N__38380),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n231_adj_744 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17729 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_14_21_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__40696),
            .in2(N__66030),
            .in3(N__38527),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n280_adj_743 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17730 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_14_21_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__65979),
            .in2(N__40687),
            .in3(N__38518),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n329_adj_740 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17731 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_14_21_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__65983),
            .in2(N__40674),
            .in3(N__38506),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n378_adj_739 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17732 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_14_21_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_14_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__40670),
            .in2(N__66032),
            .in3(N__38482),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n427_adj_738 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17733 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_14_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_14_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__45399),
            .in2(N__40675),
            .in3(N__38473),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n782_adj_735 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_LUT4_0_LC_14_22_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_LUT4_0_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_LUT4_0_LC_14_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_LUT4_0_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38470),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_adj_734_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_14_22_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_14_22_4 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_14_22_4  (
            .in0(N__48967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_14_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_14_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__63607),
            .in2(N__63889),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n63_adj_682 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18047 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_14_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_14_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__40762),
            .in2(N__63893),
            .in3(N__38458),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n112_adj_681 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18047 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18048 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_14_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_14_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__40756),
            .in2(N__63890),
            .in3(N__38563),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n161_adj_680 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18048 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18049 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_14_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_14_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__40747),
            .in2(N__63894),
            .in3(N__38560),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n210_adj_679 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18049 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18050 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_14_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_14_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__40738),
            .in2(N__63891),
            .in3(N__38557),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n259_adj_678 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18050 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18051 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_14_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_14_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__40900),
            .in2(N__63895),
            .in3(N__38554),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n308_adj_677 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18051 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18052 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_14_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_14_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__40891),
            .in2(N__63892),
            .in3(N__38551),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n357_adj_676 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18052 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18053 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_14_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_14_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__40882),
            .in2(N__63896),
            .in3(N__38548),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n406_adj_675 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18053 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18054 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_14_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_14_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__40873),
            .in2(N__63946),
            .in3(N__38545),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n455_adj_674 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18055 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_14_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_14_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__40864),
            .in2(N__63949),
            .in3(N__38542),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n504_adj_673 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18055 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18056 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_14_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_14_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__40855),
            .in2(N__63947),
            .in3(N__38539),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n553_adj_672 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18056 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18057 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_14_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_14_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__40846),
            .in2(N__63950),
            .in3(N__38638),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n602_adj_671 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18057 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18058 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_14_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_14_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__40837),
            .in2(N__63948),
            .in3(N__38635),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n651_adj_670 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18058 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18059 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_14_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_14_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__41038),
            .in2(N__63951),
            .in3(N__38632),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n700_adj_669 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18059 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18060 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_14_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_14_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__45241),
            .in2(N__41029),
            .in3(N__38620),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n754_adj_667 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18060 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_LUT4_0_LC_14_24_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_LUT4_0_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_LUT4_0_LC_14_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_LUT4_0_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38617),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_adj_668_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_14_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_14_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__63875),
            .in2(N__64237),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n60_adj_698 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18032 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_14_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_14_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__64207),
            .in2(N__38602),
            .in3(N__38590),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n109_adj_697 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18032 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18033 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_14_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_14_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__38587),
            .in2(N__64238),
            .in3(N__38578),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n158_adj_696 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18033 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18034 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_14_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_14_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__64211),
            .in2(N__38575),
            .in3(N__38749),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n207_adj_695 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18034 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18035 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_14_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_14_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__38746),
            .in2(N__64239),
            .in3(N__38737),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n256_adj_694 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18035 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18036 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_14_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_14_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__64215),
            .in2(N__38734),
            .in3(N__38722),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n305_adj_693 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18036 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18037 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_14_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_14_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__38719),
            .in2(N__64240),
            .in3(N__38710),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n354_adj_692 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18037 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18038 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_14_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_14_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__64219),
            .in2(N__38707),
            .in3(N__38695),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n403_adj_691 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18038 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18039 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_14_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_14_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__38692),
            .in2(N__64233),
            .in3(N__38683),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n452_adj_690 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18040 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_14_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_14_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__64192),
            .in2(N__38680),
            .in3(N__38668),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n501_adj_689 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18040 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18041 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_14_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_14_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__38665),
            .in2(N__64234),
            .in3(N__38656),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n550_adj_688 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18041 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18042 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_14_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_14_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__64196),
            .in2(N__38653),
            .in3(N__38641),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n599_adj_687 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18042 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18043 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_14_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_14_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__38833),
            .in2(N__64235),
            .in3(N__38824),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n648_adj_686 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18043 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18044 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_14_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_14_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__64200),
            .in2(N__38821),
            .in3(N__38809),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n697_adj_685 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18044 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18045 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_14_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_14_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__45268),
            .in2(N__38806),
            .in3(N__38782),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n750_adj_683 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18045 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_LUT4_0_LC_14_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_LUT4_0_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_LUT4_0_LC_14_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_LUT4_0_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38779),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_adj_684_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_2_LC_15_5_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_2_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_2_LC_15_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_2_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__68435),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_3_LC_15_5_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_3_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_3_LC_15_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_3_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(N__42856),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15775 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_4_LC_15_5_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_4_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_4_LC_15_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_4_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(N__38761),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15776 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_5_LC_15_5_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_5_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_5_LC_15_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_5_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(N__38755),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15777 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_6_LC_15_5_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_6_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_6_LC_15_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_6_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(N__38887),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15778 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_7_LC_15_5_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_7_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_7_LC_15_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_7_LC_15_5_5  (
            .in0(_gnd_net_),
            .in1(N__38881),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15779 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_8_LC_15_5_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_8_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_8_LC_15_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_8_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(N__38875),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15780 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_9_LC_15_5_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_9_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_9_LC_15_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_9_LC_15_5_7  (
            .in0(_gnd_net_),
            .in1(N__38869),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15781 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_10_LC_15_6_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_10_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_10_LC_15_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_10_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__38863),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_11_LC_15_6_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_11_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_11_LC_15_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_11_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(N__38857),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15783 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_12_LC_15_6_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_12_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_12_LC_15_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_12_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__38851),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15784 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_13_LC_15_6_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_13_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_13_LC_15_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_13_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__38845),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15785 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_14_LC_15_6_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_14_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_14_LC_15_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_14_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(N__38839),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15786 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_15_LC_15_6_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_15_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_15_LC_15_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_15_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__38980),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15787 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_16_LC_15_6_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_16_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_16_LC_15_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_16_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(N__38974),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15788 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_17_lut_LC_15_6_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_17_lut_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_17_lut_LC_15_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_17_lut_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(N__38968),
            .in2(_gnd_net_),
            .in3(N__38962),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15789 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_18_lut_LC_15_7_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_18_lut_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_18_lut_LC_15_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_18_lut_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__38959),
            .in2(_gnd_net_),
            .in3(N__38947),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_17 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_19_lut_LC_15_7_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_19_lut_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_19_lut_LC_15_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_19_lut_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__38944),
            .in2(_gnd_net_),
            .in3(N__38935),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15791 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_20_lut_LC_15_7_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_20_lut_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_20_lut_LC_15_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_20_lut_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__38932),
            .in2(_gnd_net_),
            .in3(N__38920),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15792 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_21_lut_LC_15_7_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_21_lut_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_21_lut_LC_15_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_21_lut_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__38917),
            .in2(_gnd_net_),
            .in3(N__38905),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15793 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_22_lut_LC_15_7_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_22_lut_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_22_lut_LC_15_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_22_lut_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__38902),
            .in2(_gnd_net_),
            .in3(N__38890),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15794 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_23_lut_LC_15_7_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_23_lut_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_23_lut_LC_15_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_23_lut_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__39079),
            .in2(_gnd_net_),
            .in3(N__39067),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_22 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15795 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_24_lut_LC_15_7_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_24_lut_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_24_lut_LC_15_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_24_lut_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__39064),
            .in2(_gnd_net_),
            .in3(N__39052),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_23 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15796 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_25_lut_LC_15_7_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_25_lut_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_25_lut_LC_15_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_25_lut_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__39049),
            .in2(_gnd_net_),
            .in3(N__39037),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15797 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_26_lut_LC_15_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_26_lut_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_26_lut_LC_15_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_26_lut_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__39034),
            .in2(_gnd_net_),
            .in3(N__39025),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_25 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_27_lut_LC_15_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_27_lut_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_27_lut_LC_15_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_27_lut_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__39157),
            .in2(_gnd_net_),
            .in3(N__39022),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15799 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_28_lut_LC_15_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_28_lut_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_28_lut_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_28_lut_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__41722),
            .in2(_gnd_net_),
            .in3(N__39019),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15800 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_29_lut_LC_15_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_29_lut_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_29_lut_LC_15_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_29_lut_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__39016),
            .in2(_gnd_net_),
            .in3(N__39007),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15801 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_30_lut_LC_15_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_30_lut_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_30_lut_LC_15_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_30_lut_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__39004),
            .in2(_gnd_net_),
            .in3(N__38995),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15802 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_31_lut_LC_15_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_31_lut_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_31_lut_LC_15_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_31_lut_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__38992),
            .in2(_gnd_net_),
            .in3(N__38983),
            .lcout(Error_sub_temp_30),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15803 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_32_lut_LC_15_8_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_32_lut_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_32_lut_LC_15_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_307_32_lut_LC_15_8_6  (
            .in0(N__39175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39166),
            .lcout(Error_sub_temp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i27_1_lut_LC_15_8_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i27_1_lut_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i27_1_lut_LC_15_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i27_1_lut_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39163),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_2_lut_LC_15_9_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_2_lut_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_2_lut_LC_15_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_2_lut_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__40390),
            .in2(N__39387),
            .in3(_gnd_net_),
            .lcout(\foc.dCurrent_3 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\foc.u_Park_Transform.n17251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_3_lut_LC_15_9_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_3_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_3_lut_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_3_lut_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__39607),
            .in2(N__39391),
            .in3(N__39130),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_2 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17251 ),
            .carryout(\foc.u_Park_Transform.n17252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_4_lut_LC_15_9_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_4_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_4_lut_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_4_lut_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__39589),
            .in2(N__39388),
            .in3(N__39118),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_3 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17252 ),
            .carryout(\foc.u_Park_Transform.n17253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_5_lut_LC_15_9_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_5_lut_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_5_lut_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_5_lut_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__39372),
            .in2(N__39568),
            .in3(N__39106),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_4 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17253 ),
            .carryout(\foc.u_Park_Transform.n17254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_6_lut_LC_15_9_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_6_lut_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_6_lut_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_6_lut_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__39547),
            .in2(N__39389),
            .in3(N__39094),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_5 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17254 ),
            .carryout(\foc.u_Park_Transform.n17255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_7_lut_LC_15_9_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_7_lut_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_7_lut_LC_15_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_7_lut_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__39376),
            .in2(N__39526),
            .in3(N__39082),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_6 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17255 ),
            .carryout(\foc.u_Park_Transform.n17256 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_8_lut_LC_15_9_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_8_lut_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_8_lut_LC_15_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_8_lut_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__39505),
            .in2(N__39390),
            .in3(N__39475),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_7 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17256 ),
            .carryout(\foc.u_Park_Transform.n17257 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_9_lut_LC_15_9_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_9_lut_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_9_lut_LC_15_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_9_lut_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__39380),
            .in2(N__39808),
            .in3(N__39460),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_8 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17257 ),
            .carryout(\foc.u_Park_Transform.n17258 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_10_lut_LC_15_10_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_10_lut_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_10_lut_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_10_lut_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__39787),
            .in2(N__39384),
            .in3(N__39445),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_9 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\foc.u_Park_Transform.n17259 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_11_lut_LC_15_10_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_11_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_11_lut_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_11_lut_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__39357),
            .in2(N__39769),
            .in3(N__39430),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_10 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17259 ),
            .carryout(\foc.u_Park_Transform.n17260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_12_lut_LC_15_10_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_12_lut_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_12_lut_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_12_lut_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__39748),
            .in2(N__39385),
            .in3(N__39418),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_11 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17260 ),
            .carryout(\foc.u_Park_Transform.n17261 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_13_lut_LC_15_10_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_13_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_13_lut_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_13_lut_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__39361),
            .in2(N__39727),
            .in3(N__39406),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_12 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17261 ),
            .carryout(\foc.u_Park_Transform.n17262 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_14_lut_LC_15_10_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_14_lut_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_14_lut_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_14_lut_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__39706),
            .in2(N__39386),
            .in3(N__39394),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_13 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17262 ),
            .carryout(\foc.u_Park_Transform.n17263 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_15_lut_LC_15_10_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_15_lut_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_15_lut_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_15_lut_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__39365),
            .in2(N__39685),
            .in3(N__39202),
            .lcout(\foc.u_Park_Transform.Product1_mul_temp_14 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17263 ),
            .carryout(\foc.u_Park_Transform.n17264 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_16_lut_LC_15_10_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_16_lut_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_16_lut_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_561_16_lut_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__39199),
            .in2(N__39664),
            .in3(N__39628),
            .lcout(\foc.u_Park_Transform.n738 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17264 ),
            .carryout(\foc.u_Park_Transform.n739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n739_THRU_LUT4_0_LC_15_10_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n739_THRU_LUT4_0_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n739_THRU_LUT4_0_LC_15_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n739_THRU_LUT4_0_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39625),
            .lcout(\foc.u_Park_Transform.n739_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_2_lut_LC_15_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_2_lut_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_2_lut_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_2_lut_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__42633),
            .in2(N__40386),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n54_adj_2095 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\foc.u_Park_Transform.n17236 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_3_lut_LC_15_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_3_lut_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_3_lut_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_3_lut_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__40367),
            .in2(N__39598),
            .in3(N__39580),
            .lcout(\foc.u_Park_Transform.n103_adj_2092 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17236 ),
            .carryout(\foc.u_Park_Transform.n17237 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_4_lut_LC_15_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_4_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_4_lut_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_4_lut_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__40368),
            .in2(N__39577),
            .in3(N__39556),
            .lcout(\foc.u_Park_Transform.n152_adj_2088 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17237 ),
            .carryout(\foc.u_Park_Transform.n17238 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_5_lut_LC_15_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_5_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_5_lut_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_5_lut_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__39553),
            .in2(N__40387),
            .in3(N__39538),
            .lcout(\foc.u_Park_Transform.n201_adj_2085 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17238 ),
            .carryout(\foc.u_Park_Transform.n17239 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_6_lut_LC_15_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_6_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_6_lut_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_6_lut_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__40372),
            .in2(N__39535),
            .in3(N__39514),
            .lcout(\foc.u_Park_Transform.n250_adj_2084 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17239 ),
            .carryout(\foc.u_Park_Transform.n17240 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_7_lut_LC_15_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_7_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_7_lut_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_7_lut_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__39511),
            .in2(N__40388),
            .in3(N__39496),
            .lcout(\foc.u_Park_Transform.n299_adj_2083 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17240 ),
            .carryout(\foc.u_Park_Transform.n17241 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_8_lut_LC_15_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_8_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_8_lut_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_8_lut_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__40376),
            .in2(N__39493),
            .in3(N__39796),
            .lcout(\foc.u_Park_Transform.n348_adj_2082 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17241 ),
            .carryout(\foc.u_Park_Transform.n17242 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_9_lut_LC_15_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_9_lut_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_9_lut_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_9_lut_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__39793),
            .in2(N__40389),
            .in3(N__39781),
            .lcout(\foc.u_Park_Transform.n397_adj_2081 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17242 ),
            .carryout(\foc.u_Park_Transform.n17243 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_10_lut_LC_15_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_10_lut_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_10_lut_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_10_lut_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__40352),
            .in2(N__39778),
            .in3(N__39757),
            .lcout(\foc.u_Park_Transform.n446_adj_2079 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\foc.u_Park_Transform.n17244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_11_lut_LC_15_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_11_lut_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_11_lut_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_11_lut_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__39754),
            .in2(N__40383),
            .in3(N__39739),
            .lcout(\foc.u_Park_Transform.n495_adj_2077 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17244 ),
            .carryout(\foc.u_Park_Transform.n17245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_12_lut_LC_15_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_12_lut_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_12_lut_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_12_lut_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__40356),
            .in2(N__39736),
            .in3(N__39715),
            .lcout(\foc.u_Park_Transform.n544_adj_2074 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17245 ),
            .carryout(\foc.u_Park_Transform.n17246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_13_lut_LC_15_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_13_lut_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_13_lut_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_13_lut_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__39712),
            .in2(N__40384),
            .in3(N__39697),
            .lcout(\foc.u_Park_Transform.n593_adj_2073 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17246 ),
            .carryout(\foc.u_Park_Transform.n17247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_14_lut_LC_15_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_14_lut_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_14_lut_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_14_lut_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__40360),
            .in2(N__39694),
            .in3(N__39673),
            .lcout(\foc.u_Park_Transform.n642_adj_2072 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17247 ),
            .carryout(\foc.u_Park_Transform.n17248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_15_lut_LC_15_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_15_lut_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_15_lut_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_15_lut_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__39670),
            .in2(N__40385),
            .in3(N__39652),
            .lcout(\foc.u_Park_Transform.n691_adj_2071 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17248 ),
            .carryout(\foc.u_Park_Transform.n17249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_16_lut_LC_15_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_16_lut_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_16_lut_LC_15_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_562_16_lut_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__40516),
            .in2(N__39916),
            .in3(N__39895),
            .lcout(\foc.u_Park_Transform.n742 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17249 ),
            .carryout(\foc.u_Park_Transform.n743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n743_THRU_LUT4_0_LC_15_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n743_THRU_LUT4_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n743_THRU_LUT4_0_LC_15_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n743_THRU_LUT4_0_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39892),
            .lcout(\foc.u_Park_Transform.n743_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_2_lut_LC_15_13_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_2_lut_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_2_lut_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_2_lut_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__42091),
            .in2(N__41689),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n60 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\foc.u_Park_Transform.n17023 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_3_lut_LC_15_13_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_3_lut_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_3_lut_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_3_lut_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__39874),
            .in2(N__42134),
            .in3(N__39868),
            .lcout(\foc.u_Park_Transform.n109 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17023 ),
            .carryout(\foc.u_Park_Transform.n17024 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_4_lut_LC_15_13_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_4_lut_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_4_lut_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_4_lut_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__42095),
            .in2(N__39865),
            .in3(N__39856),
            .lcout(\foc.u_Park_Transform.n158 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17024 ),
            .carryout(\foc.u_Park_Transform.n17025 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_5_lut_LC_15_13_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_5_lut_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_5_lut_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_5_lut_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__39853),
            .in2(N__42135),
            .in3(N__39847),
            .lcout(\foc.u_Park_Transform.n207 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17025 ),
            .carryout(\foc.u_Park_Transform.n17026 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_6_lut_LC_15_13_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_6_lut_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_6_lut_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_6_lut_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__42099),
            .in2(N__39844),
            .in3(N__39835),
            .lcout(\foc.u_Park_Transform.n256 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17026 ),
            .carryout(\foc.u_Park_Transform.n17027 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_7_lut_LC_15_13_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_7_lut_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_7_lut_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_7_lut_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__39832),
            .in2(N__42136),
            .in3(N__39826),
            .lcout(\foc.u_Park_Transform.n305 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17027 ),
            .carryout(\foc.u_Park_Transform.n17028 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_8_lut_LC_15_13_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_8_lut_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_8_lut_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_8_lut_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__42103),
            .in2(N__39823),
            .in3(N__39811),
            .lcout(\foc.u_Park_Transform.n354 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17028 ),
            .carryout(\foc.u_Park_Transform.n17029 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_9_lut_LC_15_13_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_9_lut_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_9_lut_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_9_lut_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__40012),
            .in2(N__42137),
            .in3(N__40006),
            .lcout(\foc.u_Park_Transform.n403 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17029 ),
            .carryout(\foc.u_Park_Transform.n17030 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_10_lut_LC_15_14_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_10_lut_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_10_lut_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_10_lut_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__42138),
            .in2(N__40003),
            .in3(N__39994),
            .lcout(\foc.u_Park_Transform.n452 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\foc.u_Park_Transform.n17031 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_11_lut_LC_15_14_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_11_lut_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_11_lut_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_11_lut_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__39991),
            .in2(N__42183),
            .in3(N__39985),
            .lcout(\foc.u_Park_Transform.n501 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17031 ),
            .carryout(\foc.u_Park_Transform.n17032 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_12_lut_LC_15_14_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_12_lut_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_12_lut_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_12_lut_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__42142),
            .in2(N__39982),
            .in3(N__39973),
            .lcout(\foc.u_Park_Transform.n550 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17032 ),
            .carryout(\foc.u_Park_Transform.n17033 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_13_lut_LC_15_14_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_13_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_13_lut_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_13_lut_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__39970),
            .in2(N__42184),
            .in3(N__39964),
            .lcout(\foc.u_Park_Transform.n599 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17033 ),
            .carryout(\foc.u_Park_Transform.n17034 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_14_lut_LC_15_14_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_14_lut_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_14_lut_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_14_lut_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__42146),
            .in2(N__39961),
            .in3(N__39952),
            .lcout(\foc.u_Park_Transform.n648 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17034 ),
            .carryout(\foc.u_Park_Transform.n17035 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_15_lut_LC_15_14_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_15_lut_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_15_lut_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_15_lut_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__39949),
            .in2(N__42185),
            .in3(N__39943),
            .lcout(\foc.u_Park_Transform.n697 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17035 ),
            .carryout(\foc.u_Park_Transform.n17036 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_16_lut_LC_15_14_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_16_lut_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_564_16_lut_LC_15_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_564_16_lut_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__42291),
            .in2(N__39940),
            .in3(N__39919),
            .lcout(\foc.u_Park_Transform.n750_adj_2117 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17036 ),
            .carryout(\foc.u_Park_Transform.n751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n751_THRU_LUT4_0_LC_15_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n751_THRU_LUT4_0_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n751_THRU_LUT4_0_LC_15_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n751_THRU_LUT4_0_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40108),
            .lcout(\foc.u_Park_Transform.n751_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_2_lut_LC_15_15_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_2_lut_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_2_lut_LC_15_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_2_lut_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__40303),
            .in2(N__42593),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n54 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\foc.u_Park_Transform.n17053 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_3_lut_LC_15_15_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_3_lut_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_3_lut_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_3_lut_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__42040),
            .in2(N__40350),
            .in3(N__40075),
            .lcout(\foc.u_Park_Transform.n103 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17053 ),
            .carryout(\foc.u_Park_Transform.n17054 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_4_lut_LC_15_15_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_4_lut_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_4_lut_LC_15_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_4_lut_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__40307),
            .in2(N__42025),
            .in3(N__40063),
            .lcout(\foc.u_Park_Transform.n152 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17054 ),
            .carryout(\foc.u_Park_Transform.n17055 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_5_lut_LC_15_15_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_5_lut_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_5_lut_LC_15_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_5_lut_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__41998),
            .in2(N__40351),
            .in3(N__40054),
            .lcout(\foc.u_Park_Transform.n201 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17055 ),
            .carryout(\foc.u_Park_Transform.n17056 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_6_lut_LC_15_15_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_6_lut_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_6_lut_LC_15_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_6_lut_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__40311),
            .in2(N__41980),
            .in3(N__40042),
            .lcout(\foc.u_Park_Transform.n250 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17056 ),
            .carryout(\foc.u_Park_Transform.n17057 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_7_lut_LC_15_15_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_7_lut_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_7_lut_LC_15_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_7_lut_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__40348),
            .in2(N__41956),
            .in3(N__40033),
            .lcout(\foc.u_Park_Transform.n299 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17057 ),
            .carryout(\foc.u_Park_Transform.n17058 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_8_lut_LC_15_15_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_8_lut_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_8_lut_LC_15_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_8_lut_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__40312),
            .in2(N__41935),
            .in3(N__40021),
            .lcout(\foc.u_Park_Transform.n348 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17058 ),
            .carryout(\foc.u_Park_Transform.n17059 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_9_lut_LC_15_15_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_9_lut_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_9_lut_LC_15_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_9_lut_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__40349),
            .in2(N__42469),
            .in3(N__40201),
            .lcout(\foc.u_Park_Transform.n397 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17059 ),
            .carryout(\foc.u_Park_Transform.n17060 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_10_lut_LC_15_16_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_10_lut_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_10_lut_LC_15_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_10_lut_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__40261),
            .in2(N__42448),
            .in3(N__40192),
            .lcout(\foc.u_Park_Transform.n446 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\foc.u_Park_Transform.n17061 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_11_lut_LC_15_16_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_11_lut_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_11_lut_LC_15_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_11_lut_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__42421),
            .in2(N__40301),
            .in3(N__40183),
            .lcout(\foc.u_Park_Transform.n495 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17061 ),
            .carryout(\foc.u_Park_Transform.n17062 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_12_lut_LC_15_16_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_12_lut_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_12_lut_LC_15_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_12_lut_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__40265),
            .in2(N__42403),
            .in3(N__40174),
            .lcout(\foc.u_Park_Transform.n544 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17062 ),
            .carryout(\foc.u_Park_Transform.n17063 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_13_lut_LC_15_16_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_13_lut_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_13_lut_LC_15_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_13_lut_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__42376),
            .in2(N__40302),
            .in3(N__40165),
            .lcout(\foc.u_Park_Transform.n593 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17063 ),
            .carryout(\foc.u_Park_Transform.n17064 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_14_lut_LC_15_16_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_14_lut_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_14_lut_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_14_lut_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__40269),
            .in2(N__42358),
            .in3(N__40156),
            .lcout(\foc.u_Park_Transform.n642 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17064 ),
            .carryout(\foc.u_Park_Transform.n17065 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_15_lut_LC_15_16_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_15_lut_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_15_lut_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_15_lut_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__40270),
            .in2(N__42334),
            .in3(N__40144),
            .lcout(\foc.u_Park_Transform.n691 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17065 ),
            .carryout(\foc.u_Park_Transform.n17066 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_16_lut_LC_15_16_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_16_lut_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_562_16_lut_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_562_16_lut_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__40512),
            .in2(N__42313),
            .in3(N__40129),
            .lcout(\foc.u_Park_Transform.n742_adj_2086 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17066 ),
            .carryout(\foc.u_Park_Transform.n743_adj_2096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n743_adj_2096_THRU_LUT4_0_LC_15_16_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n743_adj_2096_THRU_LUT4_0_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n743_adj_2096_THRU_LUT4_0_LC_15_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n743_adj_2096_THRU_LUT4_0_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40126),
            .lcout(\foc.u_Park_Transform.n743_adj_2096_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i5_1_lut_LC_15_17_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i5_1_lut_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i5_1_lut_LC_15_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i5_1_lut_LC_15_17_0  (
            .in0(N__40522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n27_adj_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_i501_2_lut_LC_15_17_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i501_2_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_i501_2_lut_LC_15_17_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_i501_2_lut_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40405),
            .lcout(\foc.u_Park_Transform.n741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_15_17_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_15_17_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_15_17_3.LUT_INIT=16'b1110110010100000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_15_17_3 (
            .in0(N__40501),
            .in1(N__40457),
            .in2(_gnd_net_),
            .in3(N__44912),
            .lcout(n142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i7_1_lut_LC_15_17_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i7_1_lut_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i7_1_lut_LC_15_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i7_1_lut_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40411),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i4_2_lut_LC_15_17_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i4_2_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i4_2_lut_LC_15_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i4_2_lut_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40404),
            .lcout(\foc.u_Park_Transform.n592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i2_1_lut_LC_15_17_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i2_1_lut_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i2_1_lut_LC_15_17_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i2_1_lut_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__40228),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i17_1_lut_LC_15_18_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i17_1_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i17_1_lut_LC_15_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i17_1_lut_LC_15_18_0  (
            .in0(N__40219),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i18_1_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i18_1_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i18_1_lut_LC_15_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i18_1_lut_LC_15_18_2  (
            .in0(N__40213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i12_1_lut_LC_15_18_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i12_1_lut_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i12_1_lut_LC_15_18_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i12_1_lut_LC_15_18_3  (
            .in0(N__40207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i15_1_lut_LC_15_18_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i15_1_lut_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i15_1_lut_LC_15_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i15_1_lut_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40576),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i13_1_lut_LC_15_18_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i13_1_lut_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i13_1_lut_LC_15_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i13_1_lut_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40570),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i3_1_lut_LC_15_18_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i3_1_lut_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i3_1_lut_LC_15_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i3_1_lut_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40564),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i10_1_lut_LC_15_18_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i10_1_lut_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i10_1_lut_LC_15_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i10_1_lut_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40558),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i14_1_lut_LC_15_19_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i14_1_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i14_1_lut_LC_15_19_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i14_1_lut_LC_15_19_0  (
            .in0(N__40552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i21_1_lut_LC_15_19_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i21_1_lut_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i21_1_lut_LC_15_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i21_1_lut_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40546),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i16_1_lut_LC_15_19_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i16_1_lut_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i16_1_lut_LC_15_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i16_1_lut_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40540),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i23_1_lut_LC_15_19_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i23_1_lut_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i23_1_lut_LC_15_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i23_1_lut_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40534),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i26_1_lut_LC_15_19_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i26_1_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i26_1_lut_LC_15_19_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i26_1_lut_LC_15_19_4  (
            .in0(N__40528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i25_1_lut_LC_15_19_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i25_1_lut_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i25_1_lut_LC_15_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i25_1_lut_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40621),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i11_1_lut_LC_15_19_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i11_1_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i11_1_lut_LC_15_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i11_1_lut_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40615),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n21_adj_752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_272_LC_15_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_272_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_272_LC_15_20_0 .LUT_INIT=16'b1110101011100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_272_LC_15_20_0  (
            .in0(N__65508),
            .in1(N__44687),
            .in2(N__44832),
            .in3(N__44668),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18_adj_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i27_1_lut_LC_15_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i27_1_lut_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i27_1_lut_LC_15_20_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i27_1_lut_LC_15_20_1  (
            .in0(N__40609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i19_1_lut_LC_15_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i19_1_lut_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i19_1_lut_LC_15_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i19_1_lut_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40603),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_271_LC_15_20_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_271_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_271_LC_15_20_3 .LUT_INIT=16'b1110111011000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_271_LC_15_20_3  (
            .in0(N__44667),
            .in1(N__65507),
            .in2(N__44689),
            .in3(N__44823),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_757_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_LC_15_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_LC_15_20_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_LC_15_20_4  (
            .in0(N__65510),
            .in1(N__44688),
            .in2(N__40597),
            .in3(N__44828),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19841_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_273_LC_15_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_273_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_273_LC_15_20_5 .LUT_INIT=16'b1110111011000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_273_LC_15_20_5  (
            .in0(N__40594),
            .in1(N__65509),
            .in2(N__40585),
            .in3(N__44827),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n26_adj_759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i30_1_lut_LC_15_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i30_1_lut_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i30_1_lut_LC_15_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i30_1_lut_LC_15_20_6  (
            .in0(N__40582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i24_1_lut_LC_15_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i24_1_lut_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i24_1_lut_LC_15_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i24_1_lut_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40729),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_15_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_15_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__65467),
            .in2(N__65734),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n87_adj_730 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_15_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__40828),
            .in2(N__65737),
            .in3(N__40711),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n136_adj_728 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17973 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_15_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__44779),
            .in2(N__65735),
            .in3(N__40699),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n185_adj_726 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17974 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_15_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__43048),
            .in2(N__65738),
            .in3(N__40690),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n234_adj_724 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17975 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_15_21_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__43034),
            .in2(N__65736),
            .in3(N__40678),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n283_adj_723 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17976 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17977 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_15_21_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__65697),
            .in2(N__43041),
            .in3(N__40654),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n332_adj_722 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17977 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_15_21_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__45375),
            .in2(N__43042),
            .in3(N__40639),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n786_adj_719 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17978 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_LUT4_0_LC_15_21_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_LUT4_0_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_LUT4_0_LC_15_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_LUT4_0_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40636),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_adj_721_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12078_3_lut_LC_15_22_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12078_3_lut_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12078_3_lut_LC_15_22_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i12078_3_lut_LC_15_22_0  (
            .in0(N__45049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45124),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n90_adj_729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_291_LC_15_22_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_291_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_291_LC_15_22_2 .LUT_INIT=16'b1111101011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_291_LC_15_22_2  (
            .in0(N__40802),
            .in1(N__65118),
            .in2(_gnd_net_),
            .in3(N__65284),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n7_adj_760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_274_LC_15_22_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_274_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_274_LC_15_22_3 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_274_LC_15_22_3  (
            .in0(N__45125),
            .in1(N__40803),
            .in2(N__40822),
            .in3(N__65511),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791_adj_732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_4_lut_LC_15_22_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_4_lut_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_4_lut_LC_15_22_4 .LUT_INIT=16'b0010010010110100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_4_lut_LC_15_22_4  (
            .in0(N__40804),
            .in1(N__44833),
            .in2(_gnd_net_),
            .in3(N__45126),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n790_adj_733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12680_3_lut_LC_15_22_6.C_ON=1'b0;
    defparam i12680_3_lut_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam i12680_3_lut_LC_15_22_6.LUT_INIT=16'b0011001101000100;
    LogicCell40 i12680_3_lut_LC_15_22_6 (
            .in0(N__45050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65119),
            .lcout(n794_adj_2425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_15_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__63180),
            .in2(N__63632),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n66_adj_666 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18062 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_15_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__63587),
            .in2(N__40984),
            .in3(N__40750),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n115_adj_665 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18062 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18063 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_15_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__40960),
            .in2(N__63633),
            .in3(N__40741),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n164_adj_664 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18063 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18064 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_15_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__63591),
            .in2(N__40939),
            .in3(N__40732),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n213_adj_663 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18064 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18065 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_15_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__40912),
            .in2(N__63634),
            .in3(N__40894),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n262_adj_662 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18065 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18066 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_15_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__63595),
            .in2(N__41221),
            .in3(N__40885),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n311_adj_661 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18066 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18067 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_15_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__41194),
            .in2(N__63635),
            .in3(N__40876),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n360_adj_660 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18067 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18068 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_15_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__63599),
            .in2(N__41170),
            .in3(N__40867),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n409_adj_659 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18068 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18069 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_15_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__41146),
            .in2(N__63622),
            .in3(N__40858),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n458_adj_658 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18070 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_15_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__63561),
            .in2(N__41125),
            .in3(N__40849),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n507_adj_657 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18070 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18071 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_15_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__41098),
            .in2(N__63623),
            .in3(N__40840),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n556_adj_656 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18071 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18072 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_15_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__63565),
            .in2(N__41077),
            .in3(N__40831),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n605_adj_655 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18072 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18073 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_15_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_15_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__41050),
            .in2(N__63624),
            .in3(N__41032),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n654_adj_654 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18073 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18074 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_15_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_15_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__41335),
            .in2(N__63625),
            .in3(N__41020),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n703_adj_653 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18074 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18075 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_15_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_15_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__45217),
            .in2(N__41311),
            .in3(N__41005),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n758_adj_651 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18075 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_LUT4_0_LC_15_24_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_LUT4_0_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_LUT4_0_LC_15_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_LUT4_0_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41002),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_adj_652_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_15_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_15_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__62999),
            .in2(N__63284),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n69_adj_650 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18077 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_15_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_15_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_15_25_1  (
            .in0(_gnd_net_),
            .in1(N__63229),
            .in2(N__40972),
            .in3(N__40951),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n118_adj_649 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18077 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18078 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_15_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_15_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__40948),
            .in2(N__63285),
            .in3(N__40927),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n167_adj_648 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18078 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_15_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_15_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(N__63233),
            .in2(N__40924),
            .in3(N__40903),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n216_adj_647 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18079 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_15_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_15_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_15_25_4  (
            .in0(_gnd_net_),
            .in1(N__41230),
            .in2(N__63286),
            .in3(N__41209),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n265_adj_646 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18080 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_15_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_15_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__63237),
            .in2(N__41206),
            .in3(N__41185),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n314_adj_645 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18081 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18082 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_15_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_15_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__63280),
            .in2(N__41182),
            .in3(N__41158),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n363_adj_644 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18082 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_15_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_15_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_15_25_7  (
            .in0(_gnd_net_),
            .in1(N__41155),
            .in2(N__63336),
            .in3(N__41140),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n412_adj_643 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18083 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_15_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_15_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__41137),
            .in2(N__63358),
            .in3(N__41113),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n461_adj_642 ),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_15_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_15_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__63311),
            .in2(N__41110),
            .in3(N__41089),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n510_adj_641 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18085 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_15_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_15_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__41086),
            .in2(N__63359),
            .in3(N__41065),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n559_adj_640 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18086 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_15_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_15_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(N__63315),
            .in2(N__41062),
            .in3(N__41041),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n608_adj_639 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18087 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_15_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_15_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__41344),
            .in2(N__63360),
            .in3(N__41326),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n657_adj_638 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18088 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_15_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_15_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_15_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__63319),
            .in2(N__41323),
            .in3(N__41299),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n706_adj_637 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18089 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_15_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_15_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(N__45193),
            .in2(N__41296),
            .in3(N__41272),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n762_adj_635 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18090 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_LUT4_0_LC_15_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_LUT4_0_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_LUT4_0_LC_15_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_LUT4_0_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41269),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_adj_636_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_16_7_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_16_7_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_16_7_0  (
            .in0(N__41241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_7_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_7_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__41391),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_16_7_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_16_7_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_16_7_6  (
            .in0(N__41251),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_7_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41250),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_16_8_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_16_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41242),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_8_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41380),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_16_8_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_16_8_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_16_8_3  (
            .in0(N__41367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11954_3_lut_LC_16_8_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11954_3_lut_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11954_3_lut_LC_16_8_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i11954_3_lut_LC_16_8_4  (
            .in0(N__50342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44114),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_16_8_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_16_8_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_16_8_5  (
            .in0(N__41392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_8_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_8_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41379),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_16_9_0.C_ON=1'b0;
    defparam i1_2_lut_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_16_9_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_LC_16_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50343),
            .lcout(n141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_16_9_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_16_9_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_16_9_2  (
            .in0(N__41356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_16_9_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_16_9_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_16_9_3  (
            .in0(N__41371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_16_9_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_16_9_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_16_9_4  (
            .in0(N__41355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_128_LC_16_9_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_128_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_128_LC_16_9_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_128_LC_16_9_5  (
            .in0(N__44115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i28_1_lut_LC_16_10_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i28_1_lut_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i28_1_lut_LC_16_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.sub_76_inv_0_i28_1_lut_LC_16_10_6  (
            .in0(N__41734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_2_lut_LC_16_11_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_2_lut_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_2_lut_LC_16_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_2_lut_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__41710),
            .in2(N__42215),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n60_adj_2140 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\foc.u_Park_Transform.n17206 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_3_lut_LC_16_11_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_3_lut_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_3_lut_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_3_lut_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__41530),
            .in2(N__42220),
            .in3(N__41509),
            .lcout(\foc.u_Park_Transform.n109_adj_2139 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17206 ),
            .carryout(\foc.u_Park_Transform.n17207 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_4_lut_LC_16_11_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_4_lut_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_4_lut_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_4_lut_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__42203),
            .in2(N__41506),
            .in3(N__41485),
            .lcout(\foc.u_Park_Transform.n158_adj_2137 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17207 ),
            .carryout(\foc.u_Park_Transform.n17208 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_5_lut_LC_16_11_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_5_lut_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_5_lut_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_5_lut_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__41482),
            .in2(N__42221),
            .in3(N__41461),
            .lcout(\foc.u_Park_Transform.n207_adj_2136 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17208 ),
            .carryout(\foc.u_Park_Transform.n17209 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_6_lut_LC_16_11_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_6_lut_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_6_lut_LC_16_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_6_lut_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__42207),
            .in2(N__41458),
            .in3(N__41434),
            .lcout(\foc.u_Park_Transform.n256_adj_2135 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17209 ),
            .carryout(\foc.u_Park_Transform.n17210 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_7_lut_LC_16_11_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_7_lut_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_7_lut_LC_16_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_7_lut_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__41431),
            .in2(N__42222),
            .in3(N__41407),
            .lcout(\foc.u_Park_Transform.n305_adj_2134 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17210 ),
            .carryout(\foc.u_Park_Transform.n17211 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_8_lut_LC_16_11_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_8_lut_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_8_lut_LC_16_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_8_lut_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__42211),
            .in2(N__41404),
            .in3(N__41908),
            .lcout(\foc.u_Park_Transform.n354_adj_2133 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17211 ),
            .carryout(\foc.u_Park_Transform.n17212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_9_lut_LC_16_11_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_9_lut_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_9_lut_LC_16_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_9_lut_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__41905),
            .in2(N__42223),
            .in3(N__41881),
            .lcout(\foc.u_Park_Transform.n403_adj_2132 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17212 ),
            .carryout(\foc.u_Park_Transform.n17213 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_10_lut_LC_16_12_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_10_lut_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_10_lut_LC_16_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_10_lut_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__42186),
            .in2(N__41878),
            .in3(N__41854),
            .lcout(\foc.u_Park_Transform.n452_adj_2131 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\foc.u_Park_Transform.n17214 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_11_lut_LC_16_12_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_11_lut_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_11_lut_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_11_lut_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__41851),
            .in2(N__42216),
            .in3(N__41830),
            .lcout(\foc.u_Park_Transform.n501_adj_2130 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17214 ),
            .carryout(\foc.u_Park_Transform.n17215 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_12_lut_LC_16_12_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_12_lut_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_12_lut_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_12_lut_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__42190),
            .in2(N__41827),
            .in3(N__41803),
            .lcout(\foc.u_Park_Transform.n550_adj_2129 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17215 ),
            .carryout(\foc.u_Park_Transform.n17216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_13_lut_LC_16_12_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_13_lut_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_13_lut_LC_16_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_13_lut_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__41800),
            .in2(N__42217),
            .in3(N__41782),
            .lcout(\foc.u_Park_Transform.n599_adj_2128 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17216 ),
            .carryout(\foc.u_Park_Transform.n17217 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_14_lut_LC_16_12_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_14_lut_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_14_lut_LC_16_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_14_lut_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__41779),
            .in2(N__42219),
            .in3(N__41761),
            .lcout(\foc.u_Park_Transform.n648_adj_2124 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17217 ),
            .carryout(\foc.u_Park_Transform.n17218 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_15_lut_LC_16_12_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_15_lut_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_15_lut_LC_16_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_15_lut_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__41758),
            .in2(N__42218),
            .in3(N__41737),
            .lcout(\foc.u_Park_Transform.n697_adj_2121 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17218 ),
            .carryout(\foc.u_Park_Transform.n17219 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_16_lut_LC_16_12_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_16_lut_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_16_lut_LC_16_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_add_564_16_lut_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__42295),
            .in2(N__42268),
            .in3(N__42244),
            .lcout(\foc.u_Park_Transform.n750 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17219 ),
            .carryout(\foc.u_Park_Transform.n751_adj_2142 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n751_adj_2142_THRU_LUT4_0_LC_16_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n751_adj_2142_THRU_LUT4_0_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n751_adj_2142_THRU_LUT4_0_LC_16_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n751_adj_2142_THRU_LUT4_0_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42241),
            .lcout(\foc.u_Park_Transform.n751_adj_2142_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_2_lut_LC_16_13_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_2_lut_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_2_lut_LC_16_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_2_lut_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__42130),
            .in2(N__42628),
            .in3(_gnd_net_),
            .lcout(\foc.u_Park_Transform.n57 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\foc.u_Park_Transform.n17038 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_3_lut_LC_16_13_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_3_lut_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_3_lut_LC_16_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_3_lut_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__42031),
            .in2(N__42629),
            .in3(N__42010),
            .lcout(\foc.u_Park_Transform.n106 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17038 ),
            .carryout(\foc.u_Park_Transform.n17039 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_4_lut_LC_16_13_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_4_lut_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_4_lut_LC_16_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_4_lut_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__42603),
            .in2(N__42007),
            .in3(N__41989),
            .lcout(\foc.u_Park_Transform.n155 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17039 ),
            .carryout(\foc.u_Park_Transform.n17040 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_5_lut_LC_16_13_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_5_lut_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_5_lut_LC_16_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_5_lut_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__41986),
            .in2(N__42630),
            .in3(N__41968),
            .lcout(\foc.u_Park_Transform.n204 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17040 ),
            .carryout(\foc.u_Park_Transform.n17041 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_6_lut_LC_16_13_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_6_lut_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_6_lut_LC_16_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_6_lut_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__42607),
            .in2(N__41965),
            .in3(N__41944),
            .lcout(\foc.u_Park_Transform.n253 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17041 ),
            .carryout(\foc.u_Park_Transform.n17042 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_7_lut_LC_16_13_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_7_lut_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_7_lut_LC_16_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_7_lut_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__41941),
            .in2(N__42631),
            .in3(N__41920),
            .lcout(\foc.u_Park_Transform.n302 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17042 ),
            .carryout(\foc.u_Park_Transform.n17043 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_8_lut_LC_16_13_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_8_lut_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_8_lut_LC_16_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_8_lut_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__42611),
            .in2(N__42478),
            .in3(N__42457),
            .lcout(\foc.u_Park_Transform.n351 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17043 ),
            .carryout(\foc.u_Park_Transform.n17044 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_9_lut_LC_16_13_7 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_9_lut_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_9_lut_LC_16_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_9_lut_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__42454),
            .in2(N__42632),
            .in3(N__42433),
            .lcout(\foc.u_Park_Transform.n400 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17044 ),
            .carryout(\foc.u_Park_Transform.n17045 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_10_lut_LC_16_14_0 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_10_lut_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_10_lut_LC_16_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_10_lut_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__42555),
            .in2(N__42430),
            .in3(N__42412),
            .lcout(\foc.u_Park_Transform.n449 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\foc.u_Park_Transform.n17046 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_11_lut_LC_16_14_1 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_11_lut_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_11_lut_LC_16_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_11_lut_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__42409),
            .in2(N__42594),
            .in3(N__42388),
            .lcout(\foc.u_Park_Transform.n498 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17046 ),
            .carryout(\foc.u_Park_Transform.n17047 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_12_lut_LC_16_14_2 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_12_lut_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_12_lut_LC_16_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_12_lut_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__42559),
            .in2(N__42385),
            .in3(N__42367),
            .lcout(\foc.u_Park_Transform.n547 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17047 ),
            .carryout(\foc.u_Park_Transform.n17048 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_13_lut_LC_16_14_3 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_13_lut_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_13_lut_LC_16_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_13_lut_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__42364),
            .in2(N__42595),
            .in3(N__42346),
            .lcout(\foc.u_Park_Transform.n596 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17048 ),
            .carryout(\foc.u_Park_Transform.n17049 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_14_lut_LC_16_14_4 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_14_lut_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_14_lut_LC_16_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_14_lut_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__42563),
            .in2(N__42343),
            .in3(N__42322),
            .lcout(\foc.u_Park_Transform.n645 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17049 ),
            .carryout(\foc.u_Park_Transform.n17050 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_15_lut_LC_16_14_5 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_15_lut_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_15_lut_LC_16_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_15_lut_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__42319),
            .in2(N__42596),
            .in3(N__42298),
            .lcout(\foc.u_Park_Transform.n694 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17050 ),
            .carryout(\foc.u_Park_Transform.n17051 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_16_lut_LC_16_14_6 .C_ON=1'b1;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_16_lut_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Beta_15__I_0_add_563_16_lut_LC_16_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_Park_Transform.Beta_15__I_0_add_563_16_lut_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__42796),
            .in2(N__42772),
            .in3(N__42751),
            .lcout(\foc.u_Park_Transform.n746_adj_2011 ),
            .ltout(),
            .carryin(\foc.u_Park_Transform.n17051 ),
            .carryout(\foc.u_Park_Transform.n747_adj_2012 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.n747_adj_2012_THRU_LUT4_0_LC_16_14_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.n747_adj_2012_THRU_LUT4_0_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.n747_adj_2012_THRU_LUT4_0_LC_16_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_Park_Transform.n747_adj_2012_THRU_LUT4_0_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42748),
            .lcout(\foc.u_Park_Transform.n747_adj_2012_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_3_lut_3_lut_4_lut_LC_16_15_0 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_3_lut_3_lut_4_lut_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_3_lut_3_lut_4_lut_LC_16_15_0 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \foc.u_Park_Transform.i1_3_lut_3_lut_4_lut_LC_16_15_0  (
            .in0(N__44292),
            .in1(N__44436),
            .in2(_gnd_net_),
            .in3(N__42517),
            .lcout(),
            .ltout(\foc.u_Park_Transform.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_adj_308_LC_16_15_1 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_adj_308_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_3_lut_4_lut_adj_308_LC_16_15_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \foc.u_Park_Transform.i1_3_lut_4_lut_adj_308_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__44339),
            .in2(N__42727),
            .in3(N__44435),
            .lcout(\foc.u_Park_Transform.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i6_2_lut_LC_16_15_2 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i6_2_lut_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i6_2_lut_LC_16_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i6_2_lut_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42724),
            .lcout(\foc.u_Park_Transform.n595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_2_lut_4_lut_4_lut_LC_16_15_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_2_lut_4_lut_4_lut_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_2_lut_4_lut_4_lut_LC_16_15_3 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \foc.u_Park_Transform.i1_2_lut_4_lut_4_lut_LC_16_15_3  (
            .in0(N__42516),
            .in1(N__44291),
            .in2(_gnd_net_),
            .in3(N__44434),
            .lcout(\foc.u_Park_Transform.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_16_15_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_16_15_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_16_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i9_1_lut_LC_16_17_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i9_1_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i9_1_lut_LC_16_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i9_1_lut_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42496),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i6_1_lut_LC_16_17_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i6_1_lut_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i6_1_lut_LC_16_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i6_1_lut_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42487),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i4_1_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i4_1_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i4_1_lut_LC_16_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i4_1_lut_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42880),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i8_1_lut_LC_16_17_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i8_1_lut_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i8_1_lut_LC_16_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.sub_81_inv_0_i8_1_lut_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42871),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_2_LC_16_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_2_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_2_LC_16_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_2_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__42862),
            .in2(N__42849),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15720 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_3_LC_16_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_3_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_3_LC_16_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_3_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__42826),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15720 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_4_LC_16_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_4_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_4_LC_16_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_4_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__42820),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15721 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15722 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_5_LC_16_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_5_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_5_LC_16_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_5_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__42814),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15722 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_6_LC_16_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_6_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_6_LC_16_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_6_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__42808),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15723 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15724 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_7_LC_16_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_7_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_7_LC_16_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_7_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__42802),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15724 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15725 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_8_LC_16_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_8_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_8_LC_16_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_8_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__42940),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15725 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15726 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_9_LC_16_18_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_9_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_9_LC_16_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_9_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__42934),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15726 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_10_LC_16_19_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_10_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_10_LC_16_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_10_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__42928),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_11_LC_16_19_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_11_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_11_LC_16_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_11_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__42922),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15728 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_12_LC_16_19_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_12_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_12_LC_16_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_12_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__42916),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15729 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_13_LC_16_19_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_13_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_13_LC_16_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_13_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__42910),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15730 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_14_LC_16_19_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_14_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_14_LC_16_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_14_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__42904),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15731 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_15_lut_LC_16_19_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_15_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_15_lut_LC_16_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_15_lut_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__42898),
            .in2(_gnd_net_),
            .in3(N__42892),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15732 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_16_lut_LC_16_19_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_16_lut_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_16_lut_LC_16_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_16_lut_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__42889),
            .in2(_gnd_net_),
            .in3(N__42883),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15733 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_17_lut_LC_16_19_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_17_lut_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_17_lut_LC_16_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_17_lut_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__43021),
            .in2(_gnd_net_),
            .in3(N__43015),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15734 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15735 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_18_lut_LC_16_20_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_18_lut_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_18_lut_LC_16_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_18_lut_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__43012),
            .in2(_gnd_net_),
            .in3(N__43003),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_19 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_19_lut_LC_16_20_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_19_lut_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_19_lut_LC_16_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_19_lut_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__43000),
            .in2(_gnd_net_),
            .in3(N__42994),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15736 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_20_lut_LC_16_20_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_20_lut_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_20_lut_LC_16_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_20_lut_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__42991),
            .in2(_gnd_net_),
            .in3(N__42982),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15737 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_21_lut_LC_16_20_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_21_lut_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_21_lut_LC_16_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_21_lut_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__42979),
            .in2(_gnd_net_),
            .in3(N__42973),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_22 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15738 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_22_lut_LC_16_20_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_22_lut_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_22_lut_LC_16_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_22_lut_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__42970),
            .in2(_gnd_net_),
            .in3(N__42961),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_23 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15739 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_23_lut_LC_16_20_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_23_lut_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_23_lut_LC_16_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_23_lut_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__42958),
            .in2(_gnd_net_),
            .in3(N__42952),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15740 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_24_lut_LC_16_20_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_24_lut_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_24_lut_LC_16_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_24_lut_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__42949),
            .in2(_gnd_net_),
            .in3(N__42943),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15741 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_25_lut_LC_16_20_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_25_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_25_lut_LC_16_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_25_lut_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__43120),
            .in2(_gnd_net_),
            .in3(N__43114),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15742 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_26_lut_LC_16_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_26_lut_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_26_lut_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_26_lut_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__43111),
            .in2(_gnd_net_),
            .in3(N__43099),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_27 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_27_lut_LC_16_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_27_lut_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_27_lut_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_27_lut_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__43096),
            .in2(_gnd_net_),
            .in3(N__43090),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15744 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_28_lut_LC_16_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_28_lut_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_28_lut_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_28_lut_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__43087),
            .in2(_gnd_net_),
            .in3(N__43075),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15745 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_29_lut_LC_16_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_29_lut_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_29_lut_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_29_lut_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__43072),
            .in2(_gnd_net_),
            .in3(N__43060),
            .lcout(Error_sub_temp_30_adj_2385),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15746 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_30_lut_LC_16_21_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_30_lut_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_30_lut_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_308_30_lut_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__43057),
            .in2(_gnd_net_),
            .in3(N__43051),
            .lcout(Error_sub_temp_31_adj_2384),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_3_lut_4_lut_LC_16_21_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_3_lut_4_lut_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_3_lut_4_lut_LC_16_21_5 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_3_lut_4_lut_LC_16_21_5  (
            .in0(N__44822),
            .in1(N__44767),
            .in2(_gnd_net_),
            .in3(N__45120),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n188_adj_725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_21_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_21_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i35_2_lut_LC_16_21_6  (
            .in0(N__45018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_LC_16_21_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_LC_16_21_7 .LUT_INIT=16'b1011001000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_LC_16_21_7  (
            .in0(N__44821),
            .in1(N__44766),
            .in2(_gnd_net_),
            .in3(N__45119),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n237_adj_720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_22_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_22_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i53_2_lut_LC_16_22_0  (
            .in0(N__43144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_16_22_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_16_22_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_16_22_1  (
            .in0(N__43152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_16_22_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_16_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43153),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_22_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_22_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i39_2_lut_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45072),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_16_22_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_16_22_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43131),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_22_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_22_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i525_2_lut_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43143),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_16_22_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_16_22_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_16_22_6  (
            .in0(N__46554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_16_22_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_16_22_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_16_22_7  (
            .in0(N__43132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_16_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_16_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__64947),
            .in2(N__64638),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_1 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17987 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_16_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_16_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__64588),
            .in2(N__43471),
            .in3(N__43180),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_2 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17987 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17988 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_16_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_16_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__43444),
            .in2(N__64639),
            .in3(N__43177),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_3 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17988 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17989 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_16_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_16_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__64592),
            .in2(N__43423),
            .in3(N__43174),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_4 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17989 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17990 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_16_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_16_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(N__43399),
            .in2(N__64640),
            .in3(N__43171),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_5 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17990 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17991 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_16_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_16_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__43708),
            .in2(N__64641),
            .in3(N__43168),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_6 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17991 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17992 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_16_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_16_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(N__64599),
            .in2(N__43687),
            .in3(N__43165),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_7 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17992 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17993 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_16_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_16_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__43663),
            .in2(N__64642),
            .in3(N__43162),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_8 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17993 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17994 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_16_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_16_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__43642),
            .in2(N__64643),
            .in3(N__43159),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_9 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17995 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_16_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_16_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__43621),
            .in2(N__64646),
            .in3(N__43156),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_10 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17995 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17996 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_16_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_16_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__43600),
            .in2(N__64644),
            .in3(N__43261),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_11 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17996 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17997 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_16_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_16_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__43579),
            .in2(N__64647),
            .in3(N__43258),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_12 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17997 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17998 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_16_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_16_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__43558),
            .in2(N__64645),
            .in3(N__43255),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17998 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17999 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_16_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_16_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__64612),
            .in2(N__43810),
            .in3(N__43252),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Proportional_Gain_mul_temp_14 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n17999 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18000 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_16_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_16_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_16_24_6  (
            .in0(_gnd_net_),
            .in1(N__43786),
            .in2(N__45325),
            .in3(N__43228),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n738_adj_718 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18000 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_LUT4_0_LC_16_24_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_LUT4_0_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_LUT4_0_LC_16_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_LUT4_0_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43225),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n739_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_16_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_16_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__64091),
            .in2(N__64381),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n57_adj_714 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18017 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_16_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_16_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__64323),
            .in2(N__43207),
            .in3(N__43195),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n106_adj_713 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18017 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18018 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_16_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_16_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__43192),
            .in2(N__64382),
            .in3(N__43183),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n155_adj_712 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18018 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18019 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_16_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_16_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_16_25_3  (
            .in0(_gnd_net_),
            .in1(N__64327),
            .in2(N__43387),
            .in3(N__43375),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n204_adj_711 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18019 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18020 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_16_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_16_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(N__43372),
            .in2(N__64383),
            .in3(N__43363),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n253_adj_710 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18020 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18021 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_16_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_16_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_16_25_5  (
            .in0(_gnd_net_),
            .in1(N__64331),
            .in2(N__43360),
            .in3(N__43348),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n302_adj_709 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18021 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18022 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_16_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_16_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_16_25_6  (
            .in0(_gnd_net_),
            .in1(N__43345),
            .in2(N__64384),
            .in3(N__43336),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n351_adj_708 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18022 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18023 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_16_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_16_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__64335),
            .in2(N__43333),
            .in3(N__43321),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n400_adj_707 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18023 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18024 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_16_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_16_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_16_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_16_26_0  (
            .in0(_gnd_net_),
            .in1(N__43318),
            .in2(N__64437),
            .in3(N__43306),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n449_adj_706 ),
            .ltout(),
            .carryin(bfn_16_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18025 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_16_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_16_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__64388),
            .in2(N__43303),
            .in3(N__43291),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n498_adj_705 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18025 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18026 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_16_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_16_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_16_26_2  (
            .in0(_gnd_net_),
            .in1(N__43288),
            .in2(N__64438),
            .in3(N__43279),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n547_adj_704 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18026 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18027 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_16_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_16_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_16_26_3  (
            .in0(_gnd_net_),
            .in1(N__64392),
            .in2(N__43276),
            .in3(N__43264),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n596_adj_703 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18027 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18028 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_16_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_16_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_16_26_4  (
            .in0(_gnd_net_),
            .in1(N__43546),
            .in2(N__64439),
            .in3(N__43537),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n645_adj_702 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18028 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18029 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_16_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_16_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_16_26_5  (
            .in0(_gnd_net_),
            .in1(N__64396),
            .in2(N__43534),
            .in3(N__43522),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n694_adj_701 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18029 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18030 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_16_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_16_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_16_26_6  (
            .in0(_gnd_net_),
            .in1(N__43519),
            .in2(N__45289),
            .in3(N__43495),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n746_adj_699 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18030 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_LUT4_0_LC_16_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_LUT4_0_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_LUT4_0_LC_16_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_LUT4_0_LC_16_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43492),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_adj_700_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_16_27_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_16_27_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_16_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_16_27_0  (
            .in0(_gnd_net_),
            .in1(N__64453),
            .in2(N__65004),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n54 ),
            .ltout(),
            .carryin(bfn_16_27_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18002 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_16_27_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_16_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_16_27_1  (
            .in0(_gnd_net_),
            .in1(N__64964),
            .in2(N__43456),
            .in3(N__43435),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n103 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18002 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18003 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_16_27_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_16_27_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_16_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_16_27_2  (
            .in0(_gnd_net_),
            .in1(N__43432),
            .in2(N__65005),
            .in3(N__43411),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n152 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18003 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18004 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_16_27_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_16_27_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_16_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(N__43408),
            .in2(N__65014),
            .in3(N__43390),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n201 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18004 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18005 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_16_27_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_16_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_16_27_4  (
            .in0(_gnd_net_),
            .in1(N__43717),
            .in2(N__65006),
            .in3(N__43699),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n250 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18005 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18006 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_16_27_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_16_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_16_27_5  (
            .in0(_gnd_net_),
            .in1(N__43696),
            .in2(N__65015),
            .in3(N__43675),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n299 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18006 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18007 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_16_27_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_16_27_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_16_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_16_27_6  (
            .in0(_gnd_net_),
            .in1(N__43672),
            .in2(N__65007),
            .in3(N__43654),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n348 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18007 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18008 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_16_27_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_16_27_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_16_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_16_27_7  (
            .in0(_gnd_net_),
            .in1(N__43651),
            .in2(N__65016),
            .in3(N__43633),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n397 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18008 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18009 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_16_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_16_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_16_28_0  (
            .in0(_gnd_net_),
            .in1(N__43630),
            .in2(N__65008),
            .in3(N__43612),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n446 ),
            .ltout(),
            .carryin(bfn_16_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18010 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_16_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_16_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_16_28_1  (
            .in0(_gnd_net_),
            .in1(N__43609),
            .in2(N__65011),
            .in3(N__43591),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n495 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18010 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18011 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_16_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_16_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_16_28_2  (
            .in0(_gnd_net_),
            .in1(N__43588),
            .in2(N__65009),
            .in3(N__43570),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n544 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18011 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18012 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_16_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_16_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_16_28_3  (
            .in0(_gnd_net_),
            .in1(N__43567),
            .in2(N__65012),
            .in3(N__43549),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n593 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18012 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18013 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_16_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_16_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_16_28_4  (
            .in0(_gnd_net_),
            .in1(N__43819),
            .in2(N__65010),
            .in3(N__43798),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n642 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18013 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18014 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_16_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_16_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_16_28_5  (
            .in0(_gnd_net_),
            .in1(N__43795),
            .in2(N__65013),
            .in3(N__43774),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n691_adj_717 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18014 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18015 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_16_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_16_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_16_28_6  (
            .in0(_gnd_net_),
            .in1(N__45310),
            .in2(N__43771),
            .in3(N__43747),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n742_adj_715 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18015 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_LUT4_0_LC_16_28_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_LUT4_0_LC_16_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_LUT4_0_LC_16_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_LUT4_0_LC_16_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43744),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_adj_716_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_17_5_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_17_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_2_lut_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(N__55663),
            .in2(N__55872),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n84 ),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18135 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_17_5_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_17_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_3_lut_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__55823),
            .in2(N__43912),
            .in3(N__43726),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n133 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18135 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18136 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_17_5_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_17_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_17_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_4_lut_LC_17_5_2  (
            .in0(_gnd_net_),
            .in1(N__43891),
            .in2(N__55873),
            .in3(N__43723),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n182 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18136 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18137 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_17_5_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_17_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_5_lut_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(N__55827),
            .in2(N__43879),
            .in3(N__43720),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n231 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18137 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18138 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_17_5_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_17_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_6_lut_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__43864),
            .in2(N__55874),
            .in3(N__43852),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n280 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18138 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18139 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_17_5_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_17_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_7_lut_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(N__55831),
            .in2(N__44023),
            .in3(N__43849),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n329 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18139 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18140 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_17_5_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_17_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_17_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_8_lut_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__44003),
            .in2(N__55875),
            .in3(N__43846),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n378 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18140 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18141 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_17_5_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_17_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_17_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_9_lut_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(N__55835),
            .in2(N__44008),
            .in3(N__43843),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n427 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18141 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18142 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_17_6_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_17_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_572_10_lut_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__45654),
            .in2(N__44007),
            .in3(N__43840),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n782_adj_351 ),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_LUT4_0_LC_17_6_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_LUT4_0_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_LUT4_0_LC_17_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_LUT4_0_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43837),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_adj_349_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_17_7_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_17_7_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_17_7_0  (
            .in0(N__43834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_17_7_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_17_7_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i531_2_lut_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43938),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_17_7_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_17_7_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i528_2_lut_LC_17_7_2  (
            .in0(N__43833),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_17_7_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_17_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i47_2_lut_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45582),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_17_7_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_17_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43923),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_17_7_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_17_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i57_2_lut_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43939),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_7_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_7_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43924),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_7_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_7_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_7_7  (
            .in0(N__45609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_17_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_17_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_2_lut_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__55233),
            .in2(N__55616),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n87_adj_400 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_17_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_17_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_3_lut_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__43897),
            .in2(N__55619),
            .in3(N__43882),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n136_adj_399 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18167 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18168 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_17_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_17_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_4_lut_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__43966),
            .in2(N__55617),
            .in3(N__43867),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n185_adj_398 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18168 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18169 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_17_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_17_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_5_lut_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__43975),
            .in2(N__55620),
            .in3(N__43855),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n234_adj_397 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18169 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18170 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_17_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_17_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_6_lut_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__43952),
            .in2(N__55618),
            .in3(N__44011),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n283 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18170 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18171 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_17_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_17_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_7_lut_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__55582),
            .in2(N__43959),
            .in3(N__43984),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n332 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18171 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18172 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_17_8_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_17_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_573_8_lut_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__45774),
            .in2(N__43960),
            .in3(N__43981),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n786_adj_348 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18172 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_LUT4_0_LC_17_8_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_LUT4_0_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_LUT4_0_LC_17_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_LUT4_0_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43978),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_3_lut_4_lut_LC_17_9_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_3_lut_4_lut_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_3_lut_4_lut_LC_17_9_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i2_3_lut_4_lut_LC_17_9_1  (
            .in0(N__44152),
            .in1(N__44141),
            .in2(_gnd_net_),
            .in3(N__44058),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_9_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44140),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n138 ),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_LC_17_9_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_LC_17_9_3 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_LC_17_9_3  (
            .in0(N__44139),
            .in1(N__55073),
            .in2(N__43969),
            .in3(N__54969),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_315_LC_17_9_4.C_ON=1'b0;
    defparam i1_2_lut_adj_315_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_315_LC_17_9_4.LUT_INIT=16'b0000000010101010;
    LogicCell40 i1_2_lut_adj_315_LC_17_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50362),
            .lcout(n793),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_9_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_9_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_9_5  (
            .in0(N__44166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_4_lut_LC_17_9_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_4_lut_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_4_lut_LC_17_9_6 .LUT_INIT=16'b1011001000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_4_lut_LC_17_9_6  (
            .in0(N__44057),
            .in1(N__44151),
            .in2(_gnd_net_),
            .in3(N__44138),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_17_9_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_17_9_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_17_9_7  (
            .in0(N__44167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_17_10_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_17_10_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 i1_2_lut_3_lut_LC_17_10_2 (
            .in0(N__51127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50364),
            .lcout(n142_adj_2419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11961_4_lut_LC_17_10_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11961_4_lut_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i11961_4_lut_LC_17_10_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i11961_4_lut_LC_17_10_4  (
            .in0(N__55089),
            .in1(N__44142),
            .in2(N__55266),
            .in3(N__50363),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n4 ),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_4_lut_4_lut_4_lut_LC_17_10_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_4_lut_4_lut_4_lut_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_4_lut_4_lut_4_lut_LC_17_10_5 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_4_lut_4_lut_4_lut_LC_17_10_5  (
            .in0(N__44143),
            .in1(_gnd_net_),
            .in2(N__44098),
            .in3(N__44056),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_3_lut_LC_17_11_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_3_lut_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_3_lut_LC_17_11_0 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_3_lut_LC_17_11_0  (
            .in0(N__44059),
            .in1(N__55267),
            .in2(N__44091),
            .in3(N__44087),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19269 ),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_adj_135_LC_17_11_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_adj_135_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_adj_135_LC_17_11_1 .LUT_INIT=16'b1100100100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i2_4_lut_adj_135_LC_17_11_1  (
            .in0(N__44068),
            .in1(N__45756),
            .in2(N__44095),
            .in3(N__44062),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_LC_17_11_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_LC_17_11_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_3_lut_LC_17_11_5  (
            .in0(N__55268),
            .in1(N__44060),
            .in2(N__44092),
            .in3(N__44086),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19273 ),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_129_LC_17_11_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_129_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_129_LC_17_11_6 .LUT_INIT=16'b1110110010101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_129_LC_17_11_6  (
            .in0(N__44061),
            .in1(N__45755),
            .in2(N__44032),
            .in3(N__44029),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_12_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_12_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51128),
            .lcout(n146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_3_lut_LC_17_12_6 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_3_lut_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_3_lut_LC_17_12_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \foc.u_Park_Transform.i1_3_lut_LC_17_12_6  (
            .in0(N__44323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44186),
            .lcout(),
            .ltout(\foc.u_Park_Transform.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_4_lut_adj_307_LC_17_12_7 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_307_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_307_LC_17_12_7 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \foc.u_Park_Transform.i1_4_lut_adj_307_LC_17_12_7  (
            .in0(N__44187),
            .in1(N__44239),
            .in2(N__44470),
            .in3(N__44437),
            .lcout(\foc.u_Park_Transform.n791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_4_lut_LC_17_13_3 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_4_lut_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_4_lut_LC_17_13_3 .LUT_INIT=16'b1111101010001000;
    LogicCell40 \foc.u_Park_Transform.i1_4_lut_LC_17_13_3  (
            .in0(N__44318),
            .in1(N__44368),
            .in2(N__44350),
            .in3(N__44225),
            .lcout(),
            .ltout(\foc.u_Park_Transform.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i2_4_lut_LC_17_13_4 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i2_4_lut_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i2_4_lut_LC_17_13_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \foc.u_Park_Transform.i2_4_lut_LC_17_13_4  (
            .in0(N__44226),
            .in1(N__44349),
            .in2(N__44440),
            .in3(N__44319),
            .lcout(\foc.u_Park_Transform.n19845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i28_2_lut_LC_17_14_4 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i28_2_lut_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.Alpha_15__I_0_11_i28_2_lut_LC_17_14_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_Park_Transform.Alpha_15__I_0_11_i28_2_lut_LC_17_14_4  (
            .in0(N__44422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n628),
            .ltout(n628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_4_lut_adj_305_LC_17_14_5 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_305_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_305_LC_17_14_5 .LUT_INIT=16'b1110110011100000;
    LogicCell40 \foc.u_Park_Transform.i1_4_lut_adj_305_LC_17_14_5  (
            .in0(N__44364),
            .in1(N__44313),
            .in2(N__44353),
            .in3(N__44340),
            .lcout(),
            .ltout(\foc.u_Park_Transform.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_Park_Transform.i1_4_lut_adj_306_LC_17_14_6 .C_ON=1'b0;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_306_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_Park_Transform.i1_4_lut_adj_306_LC_17_14_6 .LUT_INIT=16'b1110110010101000;
    LogicCell40 \foc.u_Park_Transform.i1_4_lut_adj_306_LC_17_14_6  (
            .in0(N__44314),
            .in1(N__44224),
            .in2(N__44197),
            .in3(N__44194),
            .lcout(\foc.u_Park_Transform.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_17_15_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_17_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__60856),
            .in2(N__67442),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n66_adj_433 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_17_15_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_17_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__44503),
            .in2(N__58905),
            .in3(N__44497),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n112 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17781 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_17_15_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_17_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__48322),
            .in2(N__54806),
            .in3(N__44494),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n161 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17782 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_17_15_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_17_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__48301),
            .in2(N__54516),
            .in3(N__44491),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n210 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17783 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_17_15_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_17_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__48277),
            .in2(N__54248),
            .in3(N__44488),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n259 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17784 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_17_15_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_17_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__48256),
            .in2(N__53990),
            .in3(N__44485),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n308_adj_368 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17785 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_17_15_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_17_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__53680),
            .in2(N__48235),
            .in3(N__44482),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n357_adj_366 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17786 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_17_15_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_17_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__53316),
            .in2(N__48211),
            .in3(N__44479),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n406_adj_363 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17787 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_17_16_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_17_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__48187),
            .in2(N__53140),
            .in3(N__44476),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n455_adj_350 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_17_16_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_17_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__48472),
            .in2(N__56182),
            .in3(N__44473),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n504 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17789 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_17_16_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_17_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__48451),
            .in2(N__55944),
            .in3(N__44542),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n553 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17790 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_17_16_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_17_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__48430),
            .in2(N__55723),
            .in3(N__44539),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n602 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17791 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_17_16_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_17_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__48409),
            .in2(N__55348),
            .in3(N__44536),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n651_adj_474 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17792 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_17_16_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_17_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__55181),
            .in2(N__48388),
            .in3(N__44533),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n700_adj_455 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17793 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_17_16_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_17_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__54946),
            .in2(N__48361),
            .in3(N__44530),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n754 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17794 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_LUT4_0_LC_17_16_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_LUT4_0_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_LUT4_0_LC_17_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_LUT4_0_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44527),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_17_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_17_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__60966),
            .in2(N__67397),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n63_adj_384 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_17_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_17_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__44524),
            .in2(N__58907),
            .in3(N__44518),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n109_adj_383 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17766 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_17_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_17_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__44515),
            .in2(N__54813),
            .in3(N__44506),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n158_adj_375 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17767 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_17_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_17_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__44656),
            .in2(N__54530),
            .in3(N__44647),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n207 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17768 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_17_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_17_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__44644),
            .in2(N__54250),
            .in3(N__44635),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n256 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17769 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_17_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_17_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__44632),
            .in2(N__54000),
            .in3(N__44623),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n305 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17770 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_17_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_17_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__44620),
            .in2(N__53722),
            .in3(N__44611),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n354_adj_367 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17771 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_17_18_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_17_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__53426),
            .in2(N__44608),
            .in3(N__44596),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n403_adj_365 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17772 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_17_19_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_17_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__44593),
            .in2(N__53210),
            .in3(N__44584),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n452_adj_362 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_17_19_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_17_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__44581),
            .in2(N__56204),
            .in3(N__44572),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n501 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17774 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_17_19_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_17_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__55960),
            .in2(N__44569),
            .in3(N__44557),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n550 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17775 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_17_19_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_17_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__44554),
            .in2(N__55738),
            .in3(N__44545),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n599 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17776 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_17_19_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_17_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__44737),
            .in2(N__55337),
            .in3(N__44728),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n648_adj_347 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17777 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_17_19_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_17_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__55182),
            .in2(N__44725),
            .in3(N__44713),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n697 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17778 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_17_19_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_17_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__54958),
            .in2(N__44710),
            .in3(N__44698),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n750 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17779 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_LUT4_0_LC_17_19_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_LUT4_0_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_LUT4_0_LC_17_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_LUT4_0_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44695),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_17_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_17_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44748),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_17_20_1.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_17_20_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_17_20_1.LUT_INIT=16'b1110110010100000;
    LogicCell40 i1_2_lut_4_lut_LC_17_20_1 (
            .in0(N__48940),
            .in1(_gnd_net_),
            .in2(N__44956),
            .in3(N__45051),
            .lcout(n142_adj_2422),
            .ltout(n142_adj_2422_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_3_lut_4_lut_LC_17_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_3_lut_4_lut_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_3_lut_4_lut_LC_17_20_2 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_3_lut_4_lut_LC_17_20_2  (
            .in0(N__44765),
            .in1(_gnd_net_),
            .in2(N__44692),
            .in3(N__45129),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755 ),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n10_adj_755_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_292_LC_17_20_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_292_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_292_LC_17_20_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_4_lut_adj_292_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__44785),
            .in2(N__44671),
            .in3(N__45128),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n14_adj_756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i49_2_lut_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44997),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i66_2_lut_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__48939),
            .in2(_gnd_net_),
            .in3(N__44942),
            .lcout(n146_adj_2423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_3_lut_4_lut_LC_17_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_3_lut_4_lut_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_3_lut_4_lut_LC_17_20_7 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_3_lut_4_lut_LC_17_20_7  (
            .in0(N__44807),
            .in1(N__44764),
            .in2(_gnd_net_),
            .in3(N__45127),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n6_adj_763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_adj_275_LC_17_21_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_adj_275_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_adj_275_LC_17_21_0 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i2_4_lut_adj_275_LC_17_21_0  (
            .in0(N__45122),
            .in1(N__65438),
            .in2(N__65264),
            .in3(N__65061),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n139_adj_727 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_21_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_21_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i61_2_lut_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45123),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_312_LC_17_21_2.C_ON=1'b0;
    defparam i1_2_lut_adj_312_LC_17_21_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_312_LC_17_21_2.LUT_INIT=16'b1000100010001000;
    LogicCell40 i1_2_lut_adj_312_LC_17_21_2 (
            .in0(N__45048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n141_adj_2421),
            .ltout(n141_adj_2421_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12085_4_lut_LC_17_21_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12085_4_lut_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i12085_4_lut_LC_17_21_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i12085_4_lut_LC_17_21_3  (
            .in0(N__65437),
            .in1(N__45121),
            .in2(N__44770),
            .in3(N__45047),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n4_adj_761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_220_LC_17_21_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_220_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_220_LC_17_21_5 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_220_LC_17_21_5  (
            .in0(N__50922),
            .in1(N__52785),
            .in2(N__50708),
            .in3(N__44983),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_17_21_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_17_21_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44749),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_21_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_21_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i534_2_lut_LC_17_21_7  (
            .in0(N__46785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_218_LC_17_22_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_218_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_218_LC_17_22_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_218_LC_17_22_0  (
            .in0(N__44971),
            .in1(N__59181),
            .in2(N__51009),
            .in3(N__51042),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_219_LC_17_22_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_219_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_219_LC_17_22_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_219_LC_17_22_1  (
            .in0(N__51190),
            .in1(N__59466),
            .in2(N__44986),
            .in3(N__52641),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_216_LC_17_22_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_216_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_216_LC_17_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_216_LC_17_22_5  (
            .in0(N__46621),
            .in1(N__46651),
            .in2(N__46687),
            .in3(N__46747),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_217_LC_17_22_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_217_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_217_LC_17_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_217_LC_17_22_6  (
            .in0(N__46716),
            .in1(N__46591),
            .in2(N__44977),
            .in3(N__46774),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1213_4_lut_LC_17_22_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1213_4_lut_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1213_4_lut_LC_17_22_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1213_4_lut_LC_17_22_7  (
            .in0(N__48840),
            .in1(N__48819),
            .in2(N__44974),
            .in3(N__48867),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_211_LC_17_23_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_211_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_211_LC_17_23_0 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_211_LC_17_23_0  (
            .in0(N__44962),
            .in1(N__59465),
            .in2(N__51197),
            .in3(N__52640),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19827_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_212_LC_17_23_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_212_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_212_LC_17_23_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_212_LC_17_23_1  (
            .in0(N__50915),
            .in1(N__52772),
            .in2(N__44965),
            .in3(N__50693),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_210_LC_17_23_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_210_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_210_LC_17_23_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_210_LC_17_23_3  (
            .in0(N__48839),
            .in1(N__51041),
            .in2(N__51008),
            .in3(N__59180),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_17_23_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_17_23_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i510_2_lut_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45148),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_17_23_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_17_23_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i522_2_lut_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46573),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_23_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_23_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i513_2_lut_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46518),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_17_23_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_17_23_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i43_2_lut_LC_17_23_7  (
            .in0(N__45147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i537_2_lut_LC_17_24_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i537_2_lut_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i537_2_lut_LC_17_24_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i537_2_lut_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45133),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_17_24_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_17_24_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i504_2_lut_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45076),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_313_LC_17_24_2.C_ON=1'b0;
    defparam i1_2_lut_adj_313_LC_17_24_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_313_LC_17_24_2.LUT_INIT=16'b0100010001000100;
    LogicCell40 i1_2_lut_adj_313_LC_17_24_2 (
            .in0(N__45055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n793_adj_2424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_17_24_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_17_24_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i498_2_lut_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45022),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i31_LC_17_24_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i31_LC_17_24_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i31_LC_17_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i31_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58367),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62112),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_17_24_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_17_24_6 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__45004),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_17_24_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_17_24_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i501_2_lut_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51082),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_17_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_17_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__45321),
            .in2(N__65017),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n93 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18369 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_17_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_17_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_17_25_1  (
            .in0(_gnd_net_),
            .in1(N__45303),
            .in2(N__64452),
            .in3(N__45292),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n142 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18369 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18370 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_17_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_17_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(N__45282),
            .in2(N__64090),
            .in3(N__45271),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n191 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18370 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18371 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_17_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_17_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_17_25_3  (
            .in0(_gnd_net_),
            .in1(N__45258),
            .in2(N__63929),
            .in3(N__45244),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n240 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18371 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18372 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_17_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_17_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_17_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(N__45237),
            .in2(N__63626),
            .in3(N__45220),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n289 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18372 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18373 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_17_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_17_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_17_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__45213),
            .in2(N__63279),
            .in3(N__45196),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n338 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18373 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18374 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_17_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_17_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_17_25_6  (
            .in0(_gnd_net_),
            .in1(N__45189),
            .in2(N__62959),
            .in3(N__45172),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n387 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18374 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18375 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_17_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_17_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(N__45162),
            .in2(N__66876),
            .in3(N__45151),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n436 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18375 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18376 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_17_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_17_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__45477),
            .in2(N__66604),
            .in3(N__45460),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n485 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18377 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_17_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_17_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__45456),
            .in2(N__66345),
            .in3(N__45433),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n534 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18377 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18378 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_17_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_17_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_17_26_2  (
            .in0(_gnd_net_),
            .in1(N__45430),
            .in2(N__66063),
            .in3(N__45406),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n583 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18378 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18379 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_17_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_17_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_17_26_3  (
            .in0(_gnd_net_),
            .in1(N__45403),
            .in2(N__65808),
            .in3(N__45382),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n632 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18379 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18380 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_17_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_17_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__65492),
            .in2(N__45379),
            .in3(N__45358),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n681 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18380 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18381 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_17_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_17_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_17_26_5  (
            .in0(_gnd_net_),
            .in1(N__65313),
            .in2(N__45355),
            .in3(N__45343),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n730 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18381 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18382 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_17_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_17_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_17_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_17_26_6  (
            .in0(_gnd_net_),
            .in1(N__45340),
            .in2(N__65152),
            .in3(N__45331),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n794 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18382 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_LUT4_0_LC_17_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_LUT4_0_LC_17_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_LUT4_0_LC_17_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_LUT4_0_LC_17_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45328),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n795_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_18_5_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_18_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_18_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_2_lut_LC_18_5_0  (
            .in0(_gnd_net_),
            .in1(N__55839),
            .in2(N__56145),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n81 ),
            .ltout(),
            .carryin(bfn_18_5_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17266 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_18_5_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_18_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_18_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_3_lut_LC_18_5_1  (
            .in0(_gnd_net_),
            .in1(N__56094),
            .in2(N__45562),
            .in3(N__45553),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n130 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17266 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_18_5_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_18_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_18_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_4_lut_LC_18_5_2  (
            .in0(_gnd_net_),
            .in1(N__45550),
            .in2(N__56146),
            .in3(N__45544),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n179 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17267 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_18_5_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_18_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_18_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_5_lut_LC_18_5_3  (
            .in0(_gnd_net_),
            .in1(N__56098),
            .in2(N__45541),
            .in3(N__45532),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n228 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17268 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_18_5_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_18_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_18_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_6_lut_LC_18_5_4  (
            .in0(_gnd_net_),
            .in1(N__45529),
            .in2(N__56147),
            .in3(N__45523),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n277 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17269 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_18_5_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_18_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_18_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_7_lut_LC_18_5_5  (
            .in0(_gnd_net_),
            .in1(N__56102),
            .in2(N__45520),
            .in3(N__45511),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n326 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17270 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17271 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_18_5_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_18_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_18_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_8_lut_LC_18_5_6  (
            .in0(_gnd_net_),
            .in1(N__45508),
            .in2(N__56148),
            .in3(N__45502),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n375 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17271 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17272 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_18_5_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_18_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_18_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_9_lut_LC_18_5_7  (
            .in0(_gnd_net_),
            .in1(N__56106),
            .in2(N__45499),
            .in3(N__45490),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n424 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17272 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17273 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_18_6_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_18_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_10_lut_LC_18_6_0  (
            .in0(_gnd_net_),
            .in1(N__45632),
            .in2(N__56038),
            .in3(N__45487),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n473 ),
            .ltout(),
            .carryin(bfn_18_6_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17274 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_18_6_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_18_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_11_lut_LC_18_6_1  (
            .in0(_gnd_net_),
            .in1(N__56013),
            .in2(N__45639),
            .in3(N__45643),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n522 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17274 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17275 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_18_6_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_18_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_571_12_lut_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(N__45672),
            .in2(N__45640),
            .in3(N__45619),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n778_adj_356 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17275 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_LUT4_0_LC_18_6_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_LUT4_0_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_LUT4_0_LC_18_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_LUT4_0_LC_18_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45616),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_adj_352_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_18_7_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_18_7_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i507_2_lut_LC_18_7_0  (
            .in0(N__45595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_18_7_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_18_7_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i519_2_lut_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45613),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_18_7_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_18_7_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i41_2_lut_LC_18_7_2  (
            .in0(N__45594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_18_7_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_18_7_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i516_2_lut_LC_18_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45583),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_18_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_18_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_2_lut_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__61236),
            .in2(N__60862),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n93 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_18_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_18_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_3_lut_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__58983),
            .in2(N__58810),
            .in3(N__45568),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n142_adj_414 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17942 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_18_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_18_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_4_lut_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(N__52572),
            .in2(N__54625),
            .in3(N__45565),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n191 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17943 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_18_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_18_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_5_lut_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__52344),
            .in2(N__54386),
            .in3(N__45697),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n240 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17944 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_18_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_18_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_6_lut_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__50154),
            .in2(N__54080),
            .in3(N__45694),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n289 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17945 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_18_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_18_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_7_lut_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__52062),
            .in2(N__53819),
            .in3(N__45691),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n338 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17946 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17947 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_18_8_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_18_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_8_lut_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(N__49956),
            .in2(N__53585),
            .in3(N__45688),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n387 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17947 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17948 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_18_8_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_18_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_9_lut_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(N__47679),
            .in2(N__53427),
            .in3(N__45685),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n436 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17948 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17949 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_18_9_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_18_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_10_lut_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(N__47472),
            .in2(N__53075),
            .in3(N__45682),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n485 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17950 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_18_9_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_18_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_11_lut_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(N__49794),
            .in2(N__56090),
            .in3(N__45679),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n534 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17950 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17951 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_18_9_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_18_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_12_lut_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__45676),
            .in2(N__55915),
            .in3(N__45661),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n583 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17951 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17952 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_18_9_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_18_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_13_lut_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(N__45658),
            .in2(N__55615),
            .in3(N__45778),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n632 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17952 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17953 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_18_9_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_18_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_14_lut_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(N__55229),
            .in2(N__45775),
            .in3(N__45760),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n681 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17953 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17954 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_18_9_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_18_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_15_lut_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(N__55093),
            .in2(N__45757),
            .in3(N__45730),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n730 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17954 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17955 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_18_9_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_18_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_575_16_lut_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__45727),
            .in2(N__55005),
            .in3(N__45721),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n794_adj_413 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17955 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_LUT4_0_LC_18_9_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_LUT4_0_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_LUT4_0_LC_18_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_LUT4_0_LC_18_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45718),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n795_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_18_10_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_18_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__60839),
            .in2(N__67296),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n84_adj_389 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17882 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_18_10_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_18_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__58755),
            .in2(N__45715),
            .in3(N__45706),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n130_adj_453 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17882 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17883 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_18_10_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_18_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__50125),
            .in2(N__54680),
            .in3(N__45703),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n179_adj_452 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17883 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17884 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_18_10_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_18_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__50104),
            .in2(N__54480),
            .in3(N__45700),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n228_adj_450 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17884 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17885 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_18_10_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_18_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(N__50083),
            .in2(N__54156),
            .in3(N__45805),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n277_adj_448 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17885 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17886 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_18_10_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_18_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__50062),
            .in2(N__53937),
            .in3(N__45802),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n326_adj_443 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17886 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17887 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_18_10_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_18_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__50038),
            .in2(N__53636),
            .in3(N__45799),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n375_adj_438 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17887 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_18_10_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_18_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__50311),
            .in2(N__53373),
            .in3(N__45796),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n424_adj_435 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17888 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_18_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_18_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__50290),
            .in2(N__53088),
            .in3(N__45793),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n473_adj_431 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_18_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_18_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__50272),
            .in2(N__56149),
            .in3(N__45790),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n522_adj_430 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17890 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_18_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__50251),
            .in2(N__55916),
            .in3(N__45787),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n571 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17891 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_18_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_18_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__50230),
            .in2(N__55659),
            .in3(N__45784),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n620 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17892 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_18_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_18_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__50209),
            .in2(N__55306),
            .in3(N__45781),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n669 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17893 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_18_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_18_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__55122),
            .in2(N__50188),
            .in3(N__45871),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n718 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17894 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_18_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_18_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__54914),
            .in2(N__50434),
            .in3(N__45868),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n778 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17895 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_LUT4_0_LC_18_11_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_LUT4_0_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_LUT4_0_LC_18_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_LUT4_0_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45865),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n779_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_18_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_18_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__60903),
            .in2(N__67351),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n81_adj_457 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17867 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_18_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__45862),
            .in2(N__58870),
            .in3(N__45856),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n127_adj_479 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17867 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17868 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_18_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_18_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__45853),
            .in2(N__54771),
            .in3(N__45844),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n176_adj_478 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17868 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17869 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_18_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_18_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__45841),
            .in2(N__54481),
            .in3(N__45832),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n225_adj_477 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17869 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17870 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_18_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_18_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__45829),
            .in2(N__54207),
            .in3(N__45820),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n274_adj_476 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17870 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17871 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_18_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_18_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__45817),
            .in2(N__53970),
            .in3(N__45808),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n323_adj_475 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17871 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17872 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_18_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_18_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__53637),
            .in2(N__45985),
            .in3(N__45973),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n372_adj_473 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17872 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17873 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_18_12_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_18_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__45970),
            .in2(N__53408),
            .in3(N__45961),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n421_adj_465 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17873 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17874 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_18_13_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_18_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__45958),
            .in2(N__53189),
            .in3(N__45949),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n470_adj_463 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17875 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_18_13_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_18_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__45946),
            .in2(N__56150),
            .in3(N__45937),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n519_adj_461 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17875 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17876 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_18_13_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_18_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__45934),
            .in2(N__55918),
            .in3(N__45925),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n568_adj_460 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17876 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17877 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_18_13_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_18_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__45922),
            .in2(N__55698),
            .in3(N__45913),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n617_adj_459 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17877 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17878 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_18_13_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_18_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__45910),
            .in2(N__55341),
            .in3(N__45901),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n666 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17878 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17879 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_18_13_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_18_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__55125),
            .in2(N__45898),
            .in3(N__45883),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n715 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17879 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17880 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_18_13_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_18_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__45880),
            .in2(N__54945),
            .in3(N__46063),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n774 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17880 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_LUT4_0_LC_18_13_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_LUT4_0_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_LUT4_0_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_LUT4_0_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46060),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_18_14_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_18_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__60958),
            .in2(N__67396),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n78_adj_480 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17841 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_18_14_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_18_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__46057),
            .in2(N__58874),
            .in3(N__46051),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n124_adj_507 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17841 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17842 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_18_14_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_18_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__46048),
            .in2(N__54773),
            .in3(N__46039),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n173_adj_506 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17842 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17843 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_18_14_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_18_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__46036),
            .in2(N__54526),
            .in3(N__46027),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n222_adj_505 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17843 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17844 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_18_14_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_18_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__46024),
            .in2(N__54220),
            .in3(N__46015),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n271_adj_503 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17844 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17845 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_18_14_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_18_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__46012),
            .in2(N__53991),
            .in3(N__46003),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n320_adj_502 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17845 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17846 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_18_14_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_18_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__53650),
            .in2(N__46000),
            .in3(N__45988),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n369_adj_501 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17846 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17847 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_18_14_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_18_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__46171),
            .in2(N__53469),
            .in3(N__46162),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n418_adj_500 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17847 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17848 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_18_15_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_18_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__46159),
            .in2(N__53211),
            .in3(N__46150),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n467_adj_499 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17849 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_18_15_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_18_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__46147),
            .in2(N__56190),
            .in3(N__46138),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n516_adj_498 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17849 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17850 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_18_15_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_18_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__46135),
            .in2(N__55945),
            .in3(N__46126),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n565_adj_497 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17850 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17851 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_18_15_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_18_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__46123),
            .in2(N__55724),
            .in3(N__46114),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n614_adj_496 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17851 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17852 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_18_15_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_18_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__46111),
            .in2(N__55349),
            .in3(N__46102),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n663_adj_494 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17852 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17853 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_18_15_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_18_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__55150),
            .in2(N__46099),
            .in3(N__46084),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n712_adj_493 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17853 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17854 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_18_15_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_18_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__54959),
            .in2(N__46081),
            .in3(N__46069),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n770 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17854 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_LUT4_0_LC_18_15_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_LUT4_0_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_LUT4_0_LC_18_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_LUT4_0_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46066),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_adj_353_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_18_16_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_18_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__60959),
            .in2(N__67465),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n75 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17826 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_18_16_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_18_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__46255),
            .in2(N__58906),
            .in3(N__46249),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n121 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17826 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17827 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_18_16_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_18_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__46246),
            .in2(N__54802),
            .in3(N__46237),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n170 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17827 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17828 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_18_16_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_18_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__46234),
            .in2(N__54517),
            .in3(N__46225),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n219 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17828 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17829 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_18_16_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_18_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__46222),
            .in2(N__54249),
            .in3(N__46213),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n268_adj_437 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17829 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17830 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_18_16_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_18_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__46210),
            .in2(N__53992),
            .in3(N__46201),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n317_adj_428 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17830 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17831 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_18_16_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_18_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__46198),
            .in2(N__53707),
            .in3(N__46189),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n366_adj_426 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17831 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17832 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_18_16_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_18_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__53474),
            .in2(N__46186),
            .in3(N__46174),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n415 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17832 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17833 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_18_17_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__46345),
            .in2(N__53190),
            .in3(N__46336),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n464_adj_423 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17834 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_18_17_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__46333),
            .in2(N__56207),
            .in3(N__46324),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n513_adj_412 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17834 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17835 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_18_17_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__46321),
            .in2(N__55946),
            .in3(N__46312),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n562_adj_378 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17835 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17836 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_18_17_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__46309),
            .in2(N__55725),
            .in3(N__46300),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n611_adj_373 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17836 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17837 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_18_17_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__46297),
            .in2(N__55378),
            .in3(N__46288),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n660_adj_372 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17837 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17838 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_18_17_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__46285),
            .in2(N__55180),
            .in3(N__46276),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n709 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17838 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17839 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_18_17_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__54987),
            .in2(N__46273),
            .in3(N__46261),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n766 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17839 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_LUT4_0_LC_18_17_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_LUT4_0_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_LUT4_0_LC_18_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_LUT4_0_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46258),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_18_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__60967),
            .in2(N__67466),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n60 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_18_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__46423),
            .in2(N__58908),
            .in3(N__46417),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n106 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17751 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_18_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__46414),
            .in2(N__54804),
            .in3(N__46408),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n155_adj_369 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17752 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_18_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__54521),
            .in2(N__46405),
            .in3(N__46396),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n204_adj_361 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17753 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_18_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__46393),
            .in2(N__54251),
            .in3(N__46387),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n253 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17754 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_18_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__46384),
            .in2(N__54001),
            .in3(N__46378),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n302_adj_364 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17755 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_18_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__46375),
            .in2(N__53711),
            .in3(N__46369),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n351 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17756 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_18_18_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_18_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__53479),
            .in2(N__46366),
            .in3(N__46357),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n400_adj_511 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17757 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_18_19_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_18_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__46354),
            .in2(N__53215),
            .in3(N__46348),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n449_adj_492 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_18_19_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__46495),
            .in2(N__56205),
            .in3(N__46489),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n498_adj_469 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17759 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_18_19_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__46486),
            .in2(N__55966),
            .in3(N__46480),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n547_adj_454 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17760 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_18_19_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__46477),
            .in2(N__55736),
            .in3(N__46471),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n596_adj_434 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17761 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_18_19_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__46468),
            .in2(N__55363),
            .in3(N__46462),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n645_adj_429 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17762 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_18_19_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__55186),
            .in2(N__46459),
            .in3(N__46450),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n694_adj_427 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17763 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_18_19_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__54988),
            .in2(N__46447),
            .in3(N__46438),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n746 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17764 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_LUT4_0_LC_18_19_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_LUT4_0_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_LUT4_0_LC_18_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_LUT4_0_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46435),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_221_LC_18_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_221_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_221_LC_18_20_1 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_221_LC_18_20_1  (
            .in0(N__59351),
            .in1(N__59151),
            .in2(N__50655),
            .in3(N__46432),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_222_LC_18_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_222_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_222_LC_18_20_2 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_222_LC_18_20_2  (
            .in0(N__52929),
            .in1(N__52704),
            .in2(N__46426),
            .in3(N__52746),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19914_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_223_LC_18_20_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_223_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_223_LC_18_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_223_LC_18_20_3  (
            .in0(N__50976),
            .in1(N__50873),
            .in2(N__46576),
            .in3(N__50949),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_215_LC_18_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_215_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_215_LC_18_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_215_LC_18_20_4  (
            .in0(N__50948),
            .in1(N__46525),
            .in2(N__50877),
            .in3(N__50975),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_18_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_18_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i51_2_lut_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46572),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_18_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_18_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i55_2_lut_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46555),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_213_LC_18_21_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_213_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_213_LC_18_21_0 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_213_LC_18_21_0  (
            .in0(N__59350),
            .in1(N__59150),
            .in2(N__50654),
            .in3(N__46537),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n20086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_214_LC_18_21_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_214_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_214_LC_18_21_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1_4_lut_adj_214_LC_18_21_1  (
            .in0(N__52928),
            .in1(N__52703),
            .in2(N__46528),
            .in3(N__52745),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.n19890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_18_21_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_18_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i45_2_lut_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46519),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15877_4_lut_LC_18_21_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15877_4_lut_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15877_4_lut_LC_18_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i15877_4_lut_LC_18_21_4  (
            .in0(N__46683),
            .in1(N__46746),
            .in2(N__46717),
            .in3(N__46773),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20858_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15889_4_lut_LC_18_21_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15889_4_lut_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i15889_4_lut_LC_18_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i15889_4_lut_LC_18_21_5  (
            .in0(N__46620),
            .in1(N__46590),
            .in2(N__46498),
            .in3(N__46650),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20870 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_18_21_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_18_21_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i59_2_lut_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46789),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_2_lut_LC_18_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_2_lut_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_2_lut_LC_18_22_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_2_lut_LC_18_22_0  (
            .in0(N__56913),
            .in1(N__57384),
            .in2(N__64693),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20174 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15883 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_3_lut_LC_18_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_3_lut_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_3_lut_LC_18_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_3_lut_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__57333),
            .in2(N__46762),
            .in3(N__46735),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_2 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15883 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15884 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_4_lut_LC_18_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_4_lut_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_4_lut_LC_18_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_4_lut_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__57297),
            .in2(N__46732),
            .in3(N__46702),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_3 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15884 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15885 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_5_lut_LC_18_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_5_lut_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_5_lut_LC_18_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_5_lut_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__46699),
            .in2(N__57276),
            .in3(N__46672),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_4 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15885 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15886 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_6_lut_LC_18_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_6_lut_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_6_lut_LC_18_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_6_lut_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(N__57219),
            .in2(N__46669),
            .in3(N__46639),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_5 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15886 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15887 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_7_lut_LC_18_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_7_lut_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_7_lut_LC_18_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_7_lut_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(N__57195),
            .in2(N__46636),
            .in3(N__46609),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_6 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15887 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_8_lut_LC_18_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_8_lut_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_8_lut_LC_18_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_8_lut_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(N__57153),
            .in2(N__46606),
            .in3(N__46579),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_7 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15888 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_9_lut_LC_18_22_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_9_lut_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_9_lut_LC_18_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_9_lut_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(N__57114),
            .in2(N__46927),
            .in3(N__46912),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_8 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15889 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_10_lut_LC_18_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_10_lut_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_10_lut_LC_18_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_10_lut_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__57852),
            .in2(N__46909),
            .in3(N__46897),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_9 ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_11_lut_LC_18_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_11_lut_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_11_lut_LC_18_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_11_lut_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__57813),
            .in2(N__46894),
            .in3(N__46879),
            .lcout(\foc.preSatVoltage_10 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15891 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_12_lut_LC_18_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_12_lut_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_12_lut_LC_18_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_12_lut_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__57744),
            .in2(N__46876),
            .in3(N__46861),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_11 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15892 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_13_lut_LC_18_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_13_lut_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_13_lut_LC_18_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_13_lut_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__57684),
            .in2(N__46858),
            .in3(N__46843),
            .lcout(\foc.preSatVoltage_12 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15893 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_14_lut_LC_18_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_14_lut_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_14_lut_LC_18_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_14_lut_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__57600),
            .in2(N__46840),
            .in3(N__46825),
            .lcout(\foc.preSatVoltage_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15894 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_15_lut_LC_18_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_15_lut_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_15_lut_LC_18_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_15_lut_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__57525),
            .in2(N__46822),
            .in3(N__46807),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_14 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15895 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15896 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_16_lut_LC_18_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_16_lut_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_16_lut_LC_18_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_16_lut_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__46804),
            .in2(N__57463),
            .in3(N__46792),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15896 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_17_lut_LC_18_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_17_lut_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_17_lut_LC_18_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_17_lut_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__58278),
            .in2(N__47104),
            .in3(N__47089),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15897 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_18_lut_LC_18_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_18_lut_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_18_lut_LC_18_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_18_lut_LC_18_24_0  (
            .in0(_gnd_net_),
            .in1(N__47086),
            .in2(N__58213),
            .in3(N__47074),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_17 ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15899 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_19_lut_LC_18_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_19_lut_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_19_lut_LC_18_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_19_lut_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__58147),
            .in2(N__47071),
            .in3(N__47053),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15899 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_20_lut_LC_18_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_20_lut_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_20_lut_LC_18_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_20_lut_LC_18_24_2  (
            .in0(_gnd_net_),
            .in1(N__58080),
            .in2(N__47050),
            .in3(N__47032),
            .lcout(\foc.preSatVoltage_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15900 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_21_lut_LC_18_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_21_lut_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_21_lut_LC_18_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_21_lut_LC_18_24_3  (
            .in0(_gnd_net_),
            .in1(N__47029),
            .in2(N__58011),
            .in3(N__47014),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15901 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_22_lut_LC_18_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_22_lut_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_22_lut_LC_18_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_22_lut_LC_18_24_4  (
            .in0(_gnd_net_),
            .in1(N__57964),
            .in2(N__47011),
            .in3(N__46993),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15902 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_23_lut_LC_18_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_23_lut_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_23_lut_LC_18_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_23_lut_LC_18_24_5  (
            .in0(_gnd_net_),
            .in1(N__57909),
            .in2(N__46990),
            .in3(N__46972),
            .lcout(\foc.preSatVoltage_22 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15903 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_24_lut_LC_18_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_24_lut_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_24_lut_LC_18_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_24_lut_LC_18_24_6  (
            .in0(_gnd_net_),
            .in1(N__58512),
            .in2(N__46969),
            .in3(N__46951),
            .lcout(\foc.preSatVoltage_23 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15904 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_25_lut_LC_18_24_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_25_lut_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_25_lut_LC_18_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_25_lut_LC_18_24_7  (
            .in0(_gnd_net_),
            .in1(N__58433),
            .in2(N__46948),
            .in3(N__46930),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15905 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_26_lut_LC_18_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_26_lut_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_26_lut_LC_18_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_26_lut_LC_18_25_0  (
            .in0(_gnd_net_),
            .in1(N__58434),
            .in2(N__47233),
            .in3(N__47218),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_25 ),
            .ltout(),
            .carryin(bfn_18_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_27_lut_LC_18_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_27_lut_LC_18_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_27_lut_LC_18_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_27_lut_LC_18_25_1  (
            .in0(_gnd_net_),
            .in1(N__47215),
            .in2(N__58450),
            .in3(N__47203),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15907 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_28_lut_LC_18_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_28_lut_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_28_lut_LC_18_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_28_lut_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__58438),
            .in2(N__47200),
            .in3(N__47182),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15908 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_29_lut_LC_18_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_29_lut_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_29_lut_LC_18_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_29_lut_LC_18_25_3  (
            .in0(_gnd_net_),
            .in1(N__47179),
            .in2(N__58451),
            .in3(N__47164),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15909 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_30_lut_LC_18_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_30_lut_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_30_lut_LC_18_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_30_lut_LC_18_25_4  (
            .in0(_gnd_net_),
            .in1(N__58442),
            .in2(N__47161),
            .in3(N__47143),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15910 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15911 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_31_lut_LC_18_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_31_lut_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_31_lut_LC_18_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_31_lut_LC_18_25_5  (
            .in0(_gnd_net_),
            .in1(N__47140),
            .in2(N__58452),
            .in3(N__47125),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_30 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15911 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_32_lut_LC_18_25_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_32_lut_LC_18_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_32_lut_LC_18_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_548_32_lut_LC_18_25_6  (
            .in0(N__47122),
            .in1(N__58446),
            .in2(_gnd_net_),
            .in3(N__47107),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Voltage_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_18_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_18_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_18_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_18_26_0  (
            .in0(_gnd_net_),
            .in1(N__64921),
            .in2(N__64726),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18354 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_18_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_18_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_18_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_18_26_1  (
            .in0(_gnd_net_),
            .in1(N__64440),
            .in2(N__47326),
            .in3(N__47317),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n139 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18354 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18355 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_18_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_18_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_18_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__64132),
            .in2(N__47314),
            .in3(N__47305),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n188 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18355 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18356 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_18_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_18_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_18_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_18_26_3  (
            .in0(_gnd_net_),
            .in1(N__63862),
            .in2(N__47302),
            .in3(N__47293),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n237 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18356 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18357 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_18_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_18_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_18_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_18_26_4  (
            .in0(_gnd_net_),
            .in1(N__47290),
            .in2(N__63608),
            .in3(N__47284),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n286 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18357 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18358 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_18_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_18_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_18_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_18_26_5  (
            .in0(_gnd_net_),
            .in1(N__47281),
            .in2(N__63361),
            .in3(N__47275),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n335 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18358 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18359 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_18_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_18_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_18_26_6  (
            .in0(_gnd_net_),
            .in1(N__47272),
            .in2(N__62974),
            .in3(N__47266),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n384 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18359 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18360 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_18_26_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_18_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_18_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_18_26_7  (
            .in0(_gnd_net_),
            .in1(N__47263),
            .in2(N__66824),
            .in3(N__47257),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n433 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18360 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18361 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_18_27_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_18_27_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_18_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_18_27_0  (
            .in0(_gnd_net_),
            .in1(N__47254),
            .in2(N__66629),
            .in3(N__47245),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n482 ),
            .ltout(),
            .carryin(bfn_18_27_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18362 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_18_27_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_18_27_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_18_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_18_27_1  (
            .in0(_gnd_net_),
            .in1(N__47242),
            .in2(N__66327),
            .in3(N__47236),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n531 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18362 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18363 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_18_27_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_18_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_18_27_2  (
            .in0(_gnd_net_),
            .in1(N__47380),
            .in2(N__66090),
            .in3(N__47374),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n580 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18363 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18364 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_18_27_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_18_27_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_18_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_18_27_3  (
            .in0(_gnd_net_),
            .in1(N__47371),
            .in2(N__65807),
            .in3(N__47365),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n629 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18364 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18365 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_18_27_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_18_27_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_18_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_18_27_4  (
            .in0(_gnd_net_),
            .in1(N__47362),
            .in2(N__65580),
            .in3(N__47356),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n678 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18365 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18366 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_18_27_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_18_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_18_27_5  (
            .in0(_gnd_net_),
            .in1(N__65341),
            .in2(N__47353),
            .in3(N__47344),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n727 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18366 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18367 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_18_27_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_18_27_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_18_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_18_27_6  (
            .in0(_gnd_net_),
            .in1(N__47341),
            .in2(N__65188),
            .in3(N__47335),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n790 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18367 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_LUT4_0_LC_18_27_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_LUT4_0_LC_18_27_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_LUT4_0_LC_18_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_LUT4_0_LC_18_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47332),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n791_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_19_5_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_19_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_19_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_2_lut_LC_19_5_0  (
            .in0(_gnd_net_),
            .in1(N__53147),
            .in2(N__53464),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n75_adj_510 ),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_19_5_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_19_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_3_lut_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__53434),
            .in2(N__49441),
            .in3(N__47329),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n124 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17641 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_19_5_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_19_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_4_lut_LC_19_5_2  (
            .in0(_gnd_net_),
            .in1(N__49708),
            .in2(N__53465),
            .in3(N__47407),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n173 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17642 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17643 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_19_5_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_19_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_5_lut_LC_19_5_3  (
            .in0(_gnd_net_),
            .in1(N__53438),
            .in2(N__49690),
            .in3(N__47404),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n222 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17643 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17644 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_19_5_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_19_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_6_lut_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(N__49666),
            .in2(N__53466),
            .in3(N__47401),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n271 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17644 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17645 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_19_5_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_19_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_7_lut_LC_19_5_5  (
            .in0(_gnd_net_),
            .in1(N__49648),
            .in2(N__53468),
            .in3(N__47398),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n320 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17645 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17646 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_19_5_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_19_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_8_lut_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(N__49627),
            .in2(N__53467),
            .in3(N__47395),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n369 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17646 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17647 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_19_5_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_19_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_9_lut_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__53445),
            .in2(N__49606),
            .in3(N__47392),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n418 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17647 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17648 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_19_6_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_19_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_19_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_10_lut_LC_19_6_0  (
            .in0(_gnd_net_),
            .in1(N__53378),
            .in2(N__49585),
            .in3(N__47389),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n467 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17649 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_19_6_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_19_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_11_lut_LC_19_6_1  (
            .in0(_gnd_net_),
            .in1(N__49561),
            .in2(N__53428),
            .in3(N__47386),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n516 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17649 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_19_6_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_19_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_12_lut_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(N__53382),
            .in2(N__49837),
            .in3(N__47383),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n565 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17650 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_19_6_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_19_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_13_lut_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(N__49825),
            .in2(N__53429),
            .in3(N__47488),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n614 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17651 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_19_6_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_19_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_14_lut_LC_19_6_4  (
            .in0(_gnd_net_),
            .in1(N__53386),
            .in2(N__49816),
            .in3(N__47485),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n663 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17652 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_19_6_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_19_6_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_19_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_15_lut_LC_19_6_5  (
            .in0(_gnd_net_),
            .in1(N__49814),
            .in2(N__53430),
            .in3(N__47482),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n712 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17653 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_19_6_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_19_6_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_19_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_569_16_lut_LC_19_6_6  (
            .in0(_gnd_net_),
            .in1(N__49815),
            .in2(N__47479),
            .in3(N__47455),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n770_adj_381 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17654 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_LUT4_0_LC_19_6_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_LUT4_0_LC_19_6_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_LUT4_0_LC_19_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_LUT4_0_LC_19_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47452),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n771_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_19_7_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_19_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_19_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_2_lut_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(N__53377),
            .in2(N__53607),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n72_adj_508 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_19_7_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_19_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_3_lut_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__53559),
            .in2(N__47449),
            .in3(N__47437),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n121_adj_504 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17626 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_19_7_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_19_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_4_lut_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(N__47434),
            .in2(N__53608),
            .in3(N__47425),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n170_adj_490 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17627 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_19_7_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_19_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_5_lut_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__53563),
            .in2(N__47422),
            .in3(N__47410),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n219_adj_472 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17628 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_19_7_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_19_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_19_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_6_lut_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(N__47608),
            .in2(N__53609),
            .in3(N__47599),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n268 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17629 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_19_7_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_19_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_19_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_7_lut_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__53567),
            .in2(N__47596),
            .in3(N__47584),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n317 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17630 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_19_7_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_19_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_8_lut_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(N__53568),
            .in2(N__47581),
            .in3(N__47569),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n366 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17631 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_19_7_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_19_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_9_lut_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(N__47566),
            .in2(N__53610),
            .in3(N__47557),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n415_adj_449 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17632 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_19_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_19_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_19_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_10_lut_LC_19_8_0  (
            .in0(_gnd_net_),
            .in1(N__47554),
            .in2(N__53693),
            .in3(N__47545),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n464 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_19_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_19_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_19_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_11_lut_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__53657),
            .in2(N__47542),
            .in3(N__47530),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n513 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17634 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_19_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_19_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_19_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_12_lut_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(N__47527),
            .in2(N__53694),
            .in3(N__47518),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n562 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17635 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_19_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_19_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_19_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_13_lut_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__53661),
            .in2(N__47515),
            .in3(N__47503),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n611 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17636 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_19_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_19_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_14_lut_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(N__47500),
            .in2(N__53695),
            .in3(N__47491),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n660 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17637 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_19_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_19_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_19_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_15_lut_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__53665),
            .in2(N__47695),
            .in3(N__47683),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n709_adj_512 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17638 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_19_8_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_19_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_19_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_568_16_lut_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(N__47680),
            .in2(N__47668),
            .in3(N__47656),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n766_adj_385 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17639 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_LUT4_0_LC_19_8_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_LUT4_0_LC_19_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_LUT4_0_LC_19_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_LUT4_0_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47653),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n767_adj_382_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_19_9_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_19_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_LC_19_9_0  (
            .in0(_gnd_net_),
            .in1(N__60796),
            .in2(N__67404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_9_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17927 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_19_9_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_19_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_3_lut_LC_19_9_1  (
            .in0(_gnd_net_),
            .in1(N__47650),
            .in2(N__58845),
            .in3(N__47644),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n139_adj_419 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17927 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17928 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_19_9_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_19_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_4_lut_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(N__47641),
            .in2(N__54714),
            .in3(N__47635),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n188_adj_418 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17928 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_19_9_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_19_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_5_lut_LC_19_9_3  (
            .in0(_gnd_net_),
            .in1(N__54433),
            .in2(N__47632),
            .in3(N__47623),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n237_adj_417 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17929 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_19_9_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_19_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_6_lut_LC_19_9_4  (
            .in0(_gnd_net_),
            .in1(N__54175),
            .in2(N__47620),
            .in3(N__47611),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n286 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17930 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_19_9_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_19_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_7_lut_LC_19_9_5  (
            .in0(_gnd_net_),
            .in1(N__47785),
            .in2(N__53938),
            .in3(N__47779),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n335 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17931 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_19_9_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_19_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_19_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_8_lut_LC_19_9_6  (
            .in0(_gnd_net_),
            .in1(N__47776),
            .in2(N__53706),
            .in3(N__47770),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n384 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17932 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_19_9_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_19_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_19_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_9_lut_LC_19_9_7  (
            .in0(_gnd_net_),
            .in1(N__47767),
            .in2(N__53284),
            .in3(N__47761),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n433 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17933 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17934 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_19_10_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_19_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_10_lut_LC_19_10_0  (
            .in0(_gnd_net_),
            .in1(N__53089),
            .in2(N__47758),
            .in3(N__47746),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n482 ),
            .ltout(),
            .carryin(bfn_19_10_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_19_10_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_19_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_11_lut_LC_19_10_1  (
            .in0(_gnd_net_),
            .in1(N__47743),
            .in2(N__56160),
            .in3(N__47737),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n531 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17935 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_19_10_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_19_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_12_lut_LC_19_10_2  (
            .in0(_gnd_net_),
            .in1(N__47734),
            .in2(N__55917),
            .in3(N__47728),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n580 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17936 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_19_10_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_19_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_13_lut_LC_19_10_3  (
            .in0(_gnd_net_),
            .in1(N__47725),
            .in2(N__55697),
            .in3(N__47719),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n629 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17937 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_19_10_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_19_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_14_lut_LC_19_10_4  (
            .in0(_gnd_net_),
            .in1(N__47716),
            .in2(N__55356),
            .in3(N__47710),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n678 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17938 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_19_10_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_19_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_15_lut_LC_19_10_5  (
            .in0(_gnd_net_),
            .in1(N__55123),
            .in2(N__47707),
            .in3(N__47698),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n727 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17939 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_19_10_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_19_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_16_lut_LC_19_10_6  (
            .in0(_gnd_net_),
            .in1(N__54996),
            .in2(N__47860),
            .in3(N__47851),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n790_adj_415 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17940 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_LUT4_0_LC_19_10_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_LUT4_0_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_LUT4_0_LC_19_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_LUT4_0_LC_19_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47848),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n791_adj_416_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_11_0  (
            .in0(_gnd_net_),
            .in1(N__60828),
            .in2(N__67405),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n90_adj_420 ),
            .ltout(),
            .carryin(bfn_19_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_11_1  (
            .in0(_gnd_net_),
            .in1(N__58780),
            .in2(N__47845),
            .in3(N__47836),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n136 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17912 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_11_2  (
            .in0(_gnd_net_),
            .in1(N__47833),
            .in2(N__54772),
            .in3(N__47824),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n185 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17913 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_11_3  (
            .in0(_gnd_net_),
            .in1(N__47821),
            .in2(N__54501),
            .in3(N__47812),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n234 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17914 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17915 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_11_4  (
            .in0(_gnd_net_),
            .in1(N__47809),
            .in2(N__54256),
            .in3(N__47800),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n283_adj_514 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17915 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17916 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_11_5  (
            .in0(_gnd_net_),
            .in1(N__47797),
            .in2(N__53942),
            .in3(N__47788),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n332_adj_513 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17916 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17917 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_11_6  (
            .in0(_gnd_net_),
            .in1(N__47977),
            .in2(N__53715),
            .in3(N__47968),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n381 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17917 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17918 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_11_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_11_7  (
            .in0(_gnd_net_),
            .in1(N__47965),
            .in2(N__53409),
            .in3(N__47956),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n430 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17918 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17919 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_12_0  (
            .in0(_gnd_net_),
            .in1(N__47953),
            .in2(N__53201),
            .in3(N__47944),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n479 ),
            .ltout(),
            .carryin(bfn_19_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17920 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_12_1  (
            .in0(_gnd_net_),
            .in1(N__47941),
            .in2(N__56197),
            .in3(N__47932),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n528 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17920 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17921 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_12_2  (
            .in0(_gnd_net_),
            .in1(N__47929),
            .in2(N__55939),
            .in3(N__47920),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n577 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17921 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17922 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_12_3  (
            .in0(_gnd_net_),
            .in1(N__47917),
            .in2(N__55717),
            .in3(N__47908),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n626 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17922 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17923 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_12_4  (
            .in0(_gnd_net_),
            .in1(N__47905),
            .in2(N__55364),
            .in3(N__47896),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n675 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17923 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17924 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_12_5  (
            .in0(_gnd_net_),
            .in1(N__55124),
            .in2(N__47893),
            .in3(N__47878),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n724 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17924 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17925 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_12_6  (
            .in0(_gnd_net_),
            .in1(N__54940),
            .in2(N__47875),
            .in3(N__47863),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n786 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17925 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_LUT4_0_LC_19_12_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_LUT4_0_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_LUT4_0_LC_19_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_LUT4_0_LC_19_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48055),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n787_adj_421_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_19_13_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_19_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_19_13_0  (
            .in0(_gnd_net_),
            .in1(N__60857),
            .in2(N__67395),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n72 ),
            .ltout(),
            .carryin(bfn_19_13_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_19_13_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_19_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(N__58866),
            .in2(N__48052),
            .in3(N__48043),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n118 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17811 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_19_13_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_19_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_19_13_2  (
            .in0(_gnd_net_),
            .in1(N__48040),
            .in2(N__54774),
            .in3(N__48031),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n167 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17812 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_19_13_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_19_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_19_13_3  (
            .in0(_gnd_net_),
            .in1(N__48028),
            .in2(N__54525),
            .in3(N__48019),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n216 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17813 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_19_13_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_19_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_19_13_4  (
            .in0(_gnd_net_),
            .in1(N__48016),
            .in2(N__54255),
            .in3(N__48007),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n265 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17814 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_19_13_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_19_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(N__48004),
            .in2(N__53969),
            .in3(N__47995),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n314_adj_401 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17815 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_19_13_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_19_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(N__53705),
            .in2(N__47992),
            .in3(N__47980),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n363_adj_380 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17816 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17817 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_19_13_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_19_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_19_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_19_13_7  (
            .in0(_gnd_net_),
            .in1(N__48172),
            .in2(N__53410),
            .in3(N__48160),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n412 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17817 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17818 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_19_14_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_19_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_19_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_19_14_0  (
            .in0(_gnd_net_),
            .in1(N__53130),
            .in2(N__48157),
            .in3(N__48145),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n461 ),
            .ltout(),
            .carryin(bfn_19_14_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17819 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_19_14_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_19_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_19_14_1  (
            .in0(_gnd_net_),
            .in1(N__48142),
            .in2(N__56189),
            .in3(N__48130),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n510 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17819 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17820 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_19_14_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_19_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(N__48127),
            .in2(N__55956),
            .in3(N__48118),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n559_adj_358 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17820 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17821 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_19_14_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_19_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_19_14_3  (
            .in0(_gnd_net_),
            .in1(N__48115),
            .in2(N__55729),
            .in3(N__48106),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n608_adj_377 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17821 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17822 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_19_14_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_19_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_19_14_4  (
            .in0(_gnd_net_),
            .in1(N__55370),
            .in2(N__48103),
            .in3(N__48091),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n657_adj_360 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17822 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17823 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_19_14_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_19_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(N__48088),
            .in2(N__55166),
            .in3(N__48076),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n706_adj_371 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17823 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17824 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_19_14_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_19_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(N__54989),
            .in2(N__48073),
            .in3(N__48061),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n762 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17824 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_LUT4_0_LC_19_14_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_LUT4_0_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_LUT4_0_LC_19_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_LUT4_0_LC_19_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48058),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_19_15_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_19_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_19_15_0  (
            .in0(_gnd_net_),
            .in1(N__60858),
            .in2(N__67455),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n69 ),
            .ltout(),
            .carryin(bfn_19_15_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_19_15_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_19_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_19_15_1  (
            .in0(_gnd_net_),
            .in1(N__48328),
            .in2(N__58904),
            .in3(N__48313),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n115 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17796 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_19_15_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_19_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_19_15_2  (
            .in0(_gnd_net_),
            .in1(N__48310),
            .in2(N__54803),
            .in3(N__48292),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n164 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17797 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_19_15_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_19_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_19_15_3  (
            .in0(_gnd_net_),
            .in1(N__54508),
            .in2(N__48289),
            .in3(N__48268),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n213 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17798 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_19_15_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_19_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_19_15_4  (
            .in0(_gnd_net_),
            .in1(N__48265),
            .in2(N__54264),
            .in3(N__48247),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n262_adj_425 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17799 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_19_15_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_19_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_19_15_5  (
            .in0(_gnd_net_),
            .in1(N__48244),
            .in2(N__53986),
            .in3(N__48223),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n311_adj_422 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17800 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_19_15_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_19_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_19_15_6  (
            .in0(_gnd_net_),
            .in1(N__48220),
            .in2(N__53728),
            .in3(N__48199),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n360 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17801 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_19_15_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_19_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_19_15_7  (
            .in0(_gnd_net_),
            .in1(N__48196),
            .in2(N__53470),
            .in3(N__48175),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n409 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17802 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_19_16_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_19_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_19_16_0  (
            .in0(_gnd_net_),
            .in1(N__53206),
            .in2(N__48484),
            .in3(N__48463),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n458 ),
            .ltout(),
            .carryin(bfn_19_16_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_19_16_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_19_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_19_16_1  (
            .in0(_gnd_net_),
            .in1(N__48460),
            .in2(N__56206),
            .in3(N__48442),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n507 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17804 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_19_16_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_19_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_19_16_2  (
            .in0(_gnd_net_),
            .in1(N__48439),
            .in2(N__55965),
            .in3(N__48421),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n556_adj_370 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17805 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_19_16_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_19_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_19_16_3  (
            .in0(_gnd_net_),
            .in1(N__48418),
            .in2(N__55722),
            .in3(N__48400),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n605_adj_462 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17806 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_19_16_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_19_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(N__48397),
            .in2(N__55366),
            .in3(N__48376),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n654_adj_456 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17807 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_19_16_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_19_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(N__55151),
            .in2(N__48373),
            .in3(N__48349),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n703_adj_359 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17808 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_19_16_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_19_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_19_16_6  (
            .in0(_gnd_net_),
            .in1(N__54997),
            .in2(N__48346),
            .in3(N__48334),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n758 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17809 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_LUT4_0_LC_19_16_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_LUT4_0_LC_19_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_LUT4_0_LC_19_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_LUT4_0_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48331),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_adj_354_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_1_LC_19_17_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_1_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_1_LC_19_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_1_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(N__51093),
            .in2(N__51097),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17711 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_2_lut_LC_19_17_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_2_lut_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_2_lut_LC_19_17_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_2_lut_LC_19_17_1  (
            .in0(N__55486),
            .in1(_gnd_net_),
            .in2(N__51158),
            .in3(N__48610),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17711 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17712 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_3_lut_LC_19_17_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_3_lut_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_3_lut_LC_19_17_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_3_lut_LC_19_17_2  (
            .in0(N__55490),
            .in1(N__50896),
            .in2(N__54862),
            .in3(N__48607),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17712 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17713 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_4_lut_LC_19_17_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_4_lut_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_4_lut_LC_19_17_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_4_lut_LC_19_17_3  (
            .in0(N__55487),
            .in1(N__48604),
            .in2(N__54841),
            .in3(N__48595),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17713 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17714 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_5_lut_LC_19_17_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_5_lut_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_5_lut_LC_19_17_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_5_lut_LC_19_17_4  (
            .in0(N__55491),
            .in1(N__48592),
            .in2(N__48580),
            .in3(N__48565),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17714 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17715 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_6_lut_LC_19_17_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_6_lut_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_6_lut_LC_19_17_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_6_lut_LC_19_17_5  (
            .in0(N__55488),
            .in1(N__48562),
            .in2(N__48547),
            .in3(N__48532),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17715 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_7_lut_LC_19_17_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_7_lut_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_7_lut_LC_19_17_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_7_lut_LC_19_17_6  (
            .in0(N__55492),
            .in1(N__48529),
            .in2(N__48523),
            .in3(N__48508),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17716 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17717 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_8_lut_LC_19_17_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_8_lut_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_8_lut_LC_19_17_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_8_lut_LC_19_17_7  (
            .in0(N__55489),
            .in1(N__48505),
            .in2(N__48496),
            .in3(N__48487),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_22 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17717 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17718 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_9_lut_LC_19_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_9_lut_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_9_lut_LC_19_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_9_lut_LC_19_18_0  (
            .in0(N__55512),
            .in1(N__48808),
            .in2(N__48799),
            .in3(N__48790),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_23 ),
            .ltout(),
            .carryin(bfn_19_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17719 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_10_lut_LC_19_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_10_lut_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_10_lut_LC_19_18_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_10_lut_LC_19_18_1  (
            .in0(N__55493),
            .in1(N__48787),
            .in2(N__48778),
            .in3(N__48769),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17719 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17720 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_11_lut_LC_19_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_11_lut_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_11_lut_LC_19_18_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_11_lut_LC_19_18_2  (
            .in0(N__55509),
            .in1(N__48766),
            .in2(N__48754),
            .in3(N__48739),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17720 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_12_lut_LC_19_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_12_lut_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_12_lut_LC_19_18_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_12_lut_LC_19_18_3  (
            .in0(N__55494),
            .in1(N__48736),
            .in2(N__48721),
            .in3(N__48706),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17721 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17722 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_13_lut_LC_19_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_13_lut_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_13_lut_LC_19_18_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_13_lut_LC_19_18_4  (
            .in0(N__55510),
            .in1(N__50404),
            .in2(N__48703),
            .in3(N__48688),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17722 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_14_lut_LC_19_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_14_lut_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_14_lut_LC_19_18_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_14_lut_LC_19_18_5  (
            .in0(N__55495),
            .in1(N__48685),
            .in2(N__50386),
            .in3(N__48676),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17723 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17724 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_15_lut_LC_19_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_15_lut_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_15_lut_LC_19_18_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_15_lut_LC_19_18_6  (
            .in0(N__55511),
            .in1(N__48673),
            .in2(N__48661),
            .in3(N__48646),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17724 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17725 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_16_lut_LC_19_18_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_16_lut_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_16_lut_LC_19_18_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_16_lut_LC_19_18_7  (
            .in0(N__55496),
            .in1(N__48643),
            .in2(N__48628),
            .in3(N__48613),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_30 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17725 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17726 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_17_lut_LC_19_19_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_17_lut_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_17_lut_LC_19_19_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_4257_17_lut_LC_19_19_0  (
            .in0(N__48889),
            .in1(N__50734),
            .in2(N__55519),
            .in3(N__48874),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6663_2_lut_LC_19_19_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6663_2_lut_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6663_2_lut_LC_19_19_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i6663_2_lut_LC_19_19_1  (
            .in0(N__56677),
            .in1(_gnd_net_),
            .in2(N__48973),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n8356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6661_2_lut_LC_19_19_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6661_2_lut_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i6661_2_lut_LC_19_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i6661_2_lut_LC_19_19_6  (
            .in0(_gnd_net_),
            .in1(N__48969),
            .in2(_gnd_net_),
            .in3(N__56676),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i7_LC_19_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i7_LC_19_20_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i7_LC_19_20_0 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i7_LC_19_20_0  (
            .in0(N__56455),
            .in1(_gnd_net_),
            .in2(N__56365),
            .in3(N__62725),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.preSatVoltage_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i9_LC_19_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i9_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i9_LC_19_20_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i9_LC_19_20_1  (
            .in0(N__60358),
            .in1(N__56456),
            .in2(_gnd_net_),
            .in3(N__56352),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i15_LC_19_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i15_LC_19_20_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i15_LC_19_20_2 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i15_LC_19_20_2  (
            .in0(N__56454),
            .in1(_gnd_net_),
            .in2(N__56364),
            .in3(N__60229),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i14_LC_19_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i14_LC_19_20_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i14_LC_19_20_4 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i14_LC_19_20_4  (
            .in0(N__56345),
            .in1(_gnd_net_),
            .in2(N__56480),
            .in3(N__60196),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i11_LC_19_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i11_LC_19_20_5 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i11_LC_19_20_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i11_LC_19_20_5  (
            .in0(N__60289),
            .in1(N__56450),
            .in2(_gnd_net_),
            .in3(N__56344),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_LC_19_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_LC_19_20_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_LC_19_20_6  (
            .in0(N__48871),
            .in1(N__48856),
            .in2(N__48850),
            .in3(N__48823),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i10_LC_19_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i10_LC_19_20_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i10_LC_19_20_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i10_LC_19_20_7  (
            .in0(N__60412),
            .in1(N__56343),
            .in2(_gnd_net_),
            .in3(N__56449),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62105),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_1_LC_19_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_1_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_1_LC_19_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_1_LC_19_21_0  (
            .in0(_gnd_net_),
            .in1(N__48987),
            .in2(N__48991),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18144 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_2_lut_LC_19_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_2_lut_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_2_lut_LC_19_21_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_2_lut_LC_19_21_1  (
            .in0(N__56817),
            .in1(N__48952),
            .in2(_gnd_net_),
            .in3(N__48919),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18144 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18145 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_3_lut_LC_19_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_3_lut_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_3_lut_LC_19_21_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_3_lut_LC_19_21_2  (
            .in0(N__56821),
            .in1(N__48916),
            .in2(N__56647),
            .in3(N__48907),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18145 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18146 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_4_lut_LC_19_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_4_lut_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_4_lut_LC_19_21_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_4_lut_LC_19_21_3  (
            .in0(N__56818),
            .in1(N__49132),
            .in2(N__56626),
            .in3(N__48904),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18146 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18147 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_5_lut_LC_19_21_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_5_lut_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_5_lut_LC_19_21_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_5_lut_LC_19_21_4  (
            .in0(N__56822),
            .in1(N__51394),
            .in2(N__49234),
            .in3(N__48901),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18147 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18148 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_6_lut_LC_19_21_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_6_lut_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_6_lut_LC_19_21_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_6_lut_LC_19_21_5  (
            .in0(N__56819),
            .in1(N__51586),
            .in2(N__51376),
            .in3(N__48898),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18148 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_7_lut_LC_19_21_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_7_lut_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_7_lut_LC_19_21_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_7_lut_LC_19_21_6  (
            .in0(N__56823),
            .in1(N__60595),
            .in2(N__51568),
            .in3(N__48895),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18149 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18150 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_8_lut_LC_19_21_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_8_lut_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_8_lut_LC_19_21_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_8_lut_LC_19_21_7  (
            .in0(N__56820),
            .in1(N__62770),
            .in2(N__60574),
            .in3(N__48892),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_22 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18150 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18151 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_9_lut_LC_19_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_9_lut_LC_19_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_9_lut_LC_19_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_9_lut_LC_19_22_0  (
            .in0(N__56813),
            .in1(N__65029),
            .in2(N__62749),
            .in3(N__49099),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_23 ),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18152 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_10_lut_LC_19_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_10_lut_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_10_lut_LC_19_22_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_10_lut_LC_19_22_1  (
            .in0(N__56806),
            .in1(N__61006),
            .in2(N__66994),
            .in3(N__49096),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18152 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18153 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_11_lut_LC_19_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_11_lut_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_11_lut_LC_19_22_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_11_lut_LC_19_22_2  (
            .in0(N__56810),
            .in1(N__58534),
            .in2(N__60985),
            .in3(N__49093),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18153 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18154 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_12_lut_LC_19_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_12_lut_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_12_lut_LC_19_22_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_12_lut_LC_19_22_3  (
            .in0(N__56807),
            .in1(N__51811),
            .in2(N__58933),
            .in3(N__49090),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18154 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18155 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_13_lut_LC_19_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_13_lut_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_13_lut_LC_19_22_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_13_lut_LC_19_22_4  (
            .in0(N__56811),
            .in1(N__49474),
            .in2(N__51790),
            .in3(N__49087),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18155 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18156 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_14_lut_LC_19_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_14_lut_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_14_lut_LC_19_22_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_14_lut_LC_19_22_5  (
            .in0(N__56808),
            .in1(N__49267),
            .in2(N__49456),
            .in3(N__49084),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18156 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18157 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_15_lut_LC_19_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_15_lut_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_15_lut_LC_19_22_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_15_lut_LC_19_22_6  (
            .in0(N__56812),
            .in1(N__49081),
            .in2(N__49252),
            .in3(N__49069),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18157 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18158 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_16_lut_LC_19_22_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_16_lut_LC_19_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_16_lut_LC_19_22_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_16_lut_LC_19_22_7  (
            .in0(N__56809),
            .in1(N__49066),
            .in2(N__49051),
            .in3(N__49036),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_30 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18158 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18159 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_17_lut_LC_19_23_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_17_lut_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_17_lut_LC_19_23_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_4259_17_lut_LC_19_23_0  (
            .in0(N__56824),
            .in1(N__49033),
            .in2(N__49021),
            .in3(N__48994),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i17_LC_19_23_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i17_LC_19_23_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i17_LC_19_23_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i17_LC_19_23_1  (
            .in0(N__56493),
            .in1(N__56367),
            .in2(_gnd_net_),
            .in3(N__57785),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62117),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i18_LC_19_23_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i18_LC_19_23_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i18_LC_19_23_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i18_LC_19_23_3  (
            .in0(N__56494),
            .in1(N__56368),
            .in2(_gnd_net_),
            .in3(N__57716),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62117),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i16_LC_19_23_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i16_LC_19_23_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i16_LC_19_23_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i16_LC_19_23_7  (
            .in0(N__56492),
            .in1(N__56366),
            .in2(_gnd_net_),
            .in3(N__60259),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62117),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_19_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_19_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_2_lut_LC_19_24_0  (
            .in0(_gnd_net_),
            .in1(N__64862),
            .in2(N__64734),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n60 ),
            .ltout(),
            .carryin(bfn_19_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18189 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_19_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_19_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_3_lut_LC_19_24_1  (
            .in0(_gnd_net_),
            .in1(N__49120),
            .in2(N__64466),
            .in3(N__49114),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n106 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18189 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18190 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_19_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_19_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_4_lut_LC_19_24_2  (
            .in0(_gnd_net_),
            .in1(N__64111),
            .in2(N__51352),
            .in3(N__49111),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n155 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18190 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18191 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_19_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_19_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_5_lut_LC_19_24_3  (
            .in0(_gnd_net_),
            .in1(N__51340),
            .in2(N__63955),
            .in3(N__49108),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n204 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18191 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18192 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_19_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_19_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_6_lut_LC_19_24_4  (
            .in0(_gnd_net_),
            .in1(N__51331),
            .in2(N__63648),
            .in3(N__49105),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n253 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18192 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18193 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_19_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_19_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_7_lut_LC_19_24_5  (
            .in0(_gnd_net_),
            .in1(N__51322),
            .in2(N__63377),
            .in3(N__49102),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n302 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18193 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18194 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_19_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_19_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_8_lut_LC_19_24_6  (
            .in0(_gnd_net_),
            .in1(N__51313),
            .in2(N__63031),
            .in3(N__49156),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n351 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18194 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18195 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_19_24_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_19_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_19_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_9_lut_LC_19_24_7  (
            .in0(_gnd_net_),
            .in1(N__51304),
            .in2(N__66823),
            .in3(N__49153),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n400 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18195 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18196 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_19_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_19_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_10_lut_LC_19_25_0  (
            .in0(_gnd_net_),
            .in1(N__51295),
            .in2(N__66608),
            .in3(N__49150),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n449 ),
            .ltout(),
            .carryin(bfn_19_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18197 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_19_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_19_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_11_lut_LC_19_25_1  (
            .in0(_gnd_net_),
            .in1(N__51454),
            .in2(N__66294),
            .in3(N__49147),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n498 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18197 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18198 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_19_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_19_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_19_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_12_lut_LC_19_25_2  (
            .in0(_gnd_net_),
            .in1(N__51445),
            .in2(N__66036),
            .in3(N__49144),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n547 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18198 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18199 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_19_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_19_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_13_lut_LC_19_25_3  (
            .in0(_gnd_net_),
            .in1(N__51436),
            .in2(N__65776),
            .in3(N__49141),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n596 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18199 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18200 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_19_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_19_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_19_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_14_lut_LC_19_25_4  (
            .in0(_gnd_net_),
            .in1(N__51427),
            .in2(N__65546),
            .in3(N__49138),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n645 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18200 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18201 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_19_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_19_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_15_lut_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__65320),
            .in2(N__51418),
            .in3(N__49135),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n694 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18201 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18202 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_19_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_19_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_16_lut_LC_19_25_6  (
            .in0(_gnd_net_),
            .in1(N__65135),
            .in2(N__51406),
            .in3(N__49123),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n746 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18202 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_LUT4_0_LC_19_25_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_LUT4_0_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_LUT4_0_LC_19_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_LUT4_0_LC_19_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49237),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n747_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_574_2_lut_LC_19_26_0  (
            .in0(_gnd_net_),
            .in1(N__64863),
            .in2(N__64727),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n90 ),
            .ltout(),
            .carryin(bfn_19_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18339 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_3_lut_LC_19_26_1  (
            .in0(_gnd_net_),
            .in1(N__49222),
            .in2(N__64470),
            .in3(N__49216),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n136 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18339 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18340 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_4_lut_LC_19_26_2  (
            .in0(_gnd_net_),
            .in1(N__64182),
            .in2(N__49213),
            .in3(N__49204),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n185 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18340 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18341 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_5_lut_LC_19_26_3  (
            .in0(_gnd_net_),
            .in1(N__49201),
            .in2(N__63962),
            .in3(N__49195),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n234 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18341 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18342 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_6_lut_LC_19_26_4  (
            .in0(_gnd_net_),
            .in1(N__49192),
            .in2(N__63682),
            .in3(N__49186),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n283 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18342 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18343 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_7_lut_LC_19_26_5  (
            .in0(_gnd_net_),
            .in1(N__49183),
            .in2(N__63400),
            .in3(N__49177),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n332 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18343 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18344 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_8_lut_LC_19_26_6  (
            .in0(_gnd_net_),
            .in1(N__49174),
            .in2(N__63099),
            .in3(N__49168),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n381 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18344 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18345 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_26_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_9_lut_LC_19_26_7  (
            .in0(_gnd_net_),
            .in1(N__49165),
            .in2(N__66828),
            .in3(N__49159),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n430 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18345 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18346 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_27_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_27_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_10_lut_LC_19_27_0  (
            .in0(_gnd_net_),
            .in1(N__66612),
            .in2(N__49336),
            .in3(N__49327),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n479 ),
            .ltout(),
            .carryin(bfn_19_27_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18347 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_27_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_27_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_11_lut_LC_19_27_1  (
            .in0(_gnd_net_),
            .in1(N__49324),
            .in2(N__66343),
            .in3(N__49318),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n528 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18347 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18348 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_27_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_27_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_12_lut_LC_19_27_2  (
            .in0(_gnd_net_),
            .in1(N__66040),
            .in2(N__49315),
            .in3(N__49306),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n577 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18348 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18349 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_27_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_27_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_13_lut_LC_19_27_3  (
            .in0(_gnd_net_),
            .in1(N__49303),
            .in2(N__65809),
            .in3(N__49297),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n626 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18349 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18350 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_27_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_27_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_14_lut_LC_19_27_4  (
            .in0(_gnd_net_),
            .in1(N__49294),
            .in2(N__65581),
            .in3(N__49288),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n675 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18350 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18351 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_27_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_27_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_15_lut_LC_19_27_5  (
            .in0(_gnd_net_),
            .in1(N__49285),
            .in2(N__65386),
            .in3(N__49279),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n724 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18351 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18352 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_27_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_27_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_16_lut_LC_19_27_6  (
            .in0(_gnd_net_),
            .in1(N__65171),
            .in2(N__49276),
            .in3(N__49258),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n786 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18352 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_LUT4_0_LC_19_27_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_LUT4_0_LC_19_27_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_LUT4_0_LC_19_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_LUT4_0_LC_19_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49255),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n787_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_19_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_19_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_19_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_19_28_0  (
            .in0(_gnd_net_),
            .in1(N__64747),
            .in2(N__64955),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n87 ),
            .ltout(),
            .carryin(bfn_19_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18324 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_19_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_19_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_19_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_19_28_1  (
            .in0(_gnd_net_),
            .in1(N__64471),
            .in2(N__49432),
            .in3(N__49423),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n133 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18324 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18325 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_19_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_19_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_19_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_19_28_2  (
            .in0(_gnd_net_),
            .in1(N__49420),
            .in2(N__64231),
            .in3(N__49411),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n182 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18325 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18326 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_19_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_19_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_19_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_19_28_3  (
            .in0(_gnd_net_),
            .in1(N__63975),
            .in2(N__49408),
            .in3(N__49396),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n231 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18326 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18327 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_19_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_19_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_19_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_19_28_4  (
            .in0(_gnd_net_),
            .in1(N__49393),
            .in2(N__63688),
            .in3(N__49384),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n280 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18327 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18328 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_19_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_19_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__49381),
            .in2(N__63389),
            .in3(N__49372),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n329 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18328 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18329 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_19_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_19_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_19_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_19_28_6  (
            .in0(_gnd_net_),
            .in1(N__49369),
            .in2(N__63127),
            .in3(N__49360),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n378 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18329 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18330 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_19_28_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_19_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_19_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_19_28_7  (
            .in0(_gnd_net_),
            .in1(N__49357),
            .in2(N__66880),
            .in3(N__49348),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n427 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18330 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18331 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_19_29_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_19_29_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_19_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_19_29_0  (
            .in0(_gnd_net_),
            .in1(N__49345),
            .in2(N__66630),
            .in3(N__49552),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n476 ),
            .ltout(),
            .carryin(bfn_19_29_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18332 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_19_29_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_19_29_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_19_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_19_29_1  (
            .in0(_gnd_net_),
            .in1(N__49549),
            .in2(N__66344),
            .in3(N__49540),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n525 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18332 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18333 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_19_29_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_19_29_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_19_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_19_29_2  (
            .in0(_gnd_net_),
            .in1(N__49537),
            .in2(N__66092),
            .in3(N__49528),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n574 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18333 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18334 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_19_29_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_19_29_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_19_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_19_29_3  (
            .in0(_gnd_net_),
            .in1(N__49525),
            .in2(N__65845),
            .in3(N__49516),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n623 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18334 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18335 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_19_29_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_19_29_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_19_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_19_29_4  (
            .in0(_gnd_net_),
            .in1(N__49513),
            .in2(N__65582),
            .in3(N__49504),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n672 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18335 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18336 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_19_29_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_19_29_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_19_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_19_29_5  (
            .in0(_gnd_net_),
            .in1(N__65374),
            .in2(N__49501),
            .in3(N__49486),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n721 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18336 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18337 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_19_29_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_19_29_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_19_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_19_29_6  (
            .in0(_gnd_net_),
            .in1(N__49483),
            .in2(N__65169),
            .in3(N__49462),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n782 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18337 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_LUT4_0_LC_19_29_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_LUT4_0_LC_19_29_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_LUT4_0_LC_19_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_LUT4_0_LC_19_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49459),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n783_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_20_5_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_20_5_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_20_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_2_lut_LC_20_5_0  (
            .in0(_gnd_net_),
            .in1(N__56121),
            .in2(N__53197),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n78 ),
            .ltout(),
            .carryin(bfn_20_5_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18122 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_20_5_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_20_5_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_20_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_3_lut_LC_20_5_1  (
            .in0(_gnd_net_),
            .in1(N__53161),
            .in2(N__49720),
            .in3(N__49702),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n127 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18122 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18123 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_20_5_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_20_5_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_20_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_4_lut_LC_20_5_2  (
            .in0(_gnd_net_),
            .in1(N__49699),
            .in2(N__53198),
            .in3(N__49681),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n176 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18123 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18124 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_20_5_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_20_5_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_20_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_5_lut_LC_20_5_3  (
            .in0(_gnd_net_),
            .in1(N__53165),
            .in2(N__49678),
            .in3(N__49660),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n225 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18124 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18125 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_20_5_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_20_5_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_20_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_6_lut_LC_20_5_4  (
            .in0(_gnd_net_),
            .in1(N__49657),
            .in2(N__53199),
            .in3(N__49642),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n274 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18125 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18126 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_20_5_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_20_5_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_20_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_7_lut_LC_20_5_5  (
            .in0(_gnd_net_),
            .in1(N__53169),
            .in2(N__49639),
            .in3(N__49621),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n323 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18126 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18127 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_20_5_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_20_5_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_20_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_8_lut_LC_20_5_6  (
            .in0(_gnd_net_),
            .in1(N__53170),
            .in2(N__49618),
            .in3(N__49597),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n372 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18127 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18128 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_20_5_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_20_5_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_20_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_9_lut_LC_20_5_7  (
            .in0(_gnd_net_),
            .in1(N__49594),
            .in2(N__53200),
            .in3(N__49576),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n421 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18128 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18129 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_20_6_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_20_6_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_20_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_10_lut_LC_20_6_0  (
            .in0(_gnd_net_),
            .in1(N__49573),
            .in2(N__53194),
            .in3(N__49555),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n470 ),
            .ltout(),
            .carryin(bfn_20_6_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18130 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_20_6_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_20_6_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_20_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_11_lut_LC_20_6_1  (
            .in0(_gnd_net_),
            .in1(N__49846),
            .in2(N__53196),
            .in3(N__49828),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n519 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18130 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18131 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_20_6_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_20_6_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_20_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_12_lut_LC_20_6_2  (
            .in0(_gnd_net_),
            .in1(N__49763),
            .in2(N__53195),
            .in3(N__49819),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n568 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18131 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18132 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_20_6_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_20_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_13_lut_LC_20_6_3  (
            .in0(_gnd_net_),
            .in1(N__53154),
            .in2(N__49770),
            .in3(N__49798),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n617 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18132 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n18133 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_20_6_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_20_6_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_20_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_570_14_lut_LC_20_6_4  (
            .in0(_gnd_net_),
            .in1(N__49795),
            .in2(N__49771),
            .in3(N__49747),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n774_adj_374 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n18133 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_LUT4_0_LC_20_6_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_LUT4_0_LC_20_6_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_LUT4_0_LC_20_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_LUT4_0_LC_20_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49744),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n775_adj_357_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_20_7_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_20_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_2_lut_LC_20_7_0  (
            .in0(_gnd_net_),
            .in1(N__53611),
            .in2(N__53881),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n69_adj_489 ),
            .ltout(),
            .carryin(bfn_20_7_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_20_7_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_20_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_3_lut_LC_20_7_1  (
            .in0(_gnd_net_),
            .in1(N__49741),
            .in2(N__53884),
            .in3(N__49735),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n118_adj_487 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17611 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17612 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_20_7_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_20_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_4_lut_LC_20_7_2  (
            .in0(_gnd_net_),
            .in1(N__53832),
            .in2(N__49732),
            .in3(N__49723),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n167_adj_486 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17612 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17613 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_20_7_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_20_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_5_lut_LC_20_7_3  (
            .in0(_gnd_net_),
            .in1(N__49930),
            .in2(N__53885),
            .in3(N__49924),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n216_adj_485 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17613 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17614 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_20_7_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_20_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_6_lut_LC_20_7_4  (
            .in0(_gnd_net_),
            .in1(N__49921),
            .in2(N__53882),
            .in3(N__49915),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n265_adj_471 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17614 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17615 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_20_7_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_20_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_7_lut_LC_20_7_5  (
            .in0(_gnd_net_),
            .in1(N__49912),
            .in2(N__53886),
            .in3(N__49906),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n314 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17615 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17616 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_20_7_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_20_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_8_lut_LC_20_7_6  (
            .in0(_gnd_net_),
            .in1(N__49903),
            .in2(N__53883),
            .in3(N__49897),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n363 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17616 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17617 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_20_7_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_20_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_9_lut_LC_20_7_7  (
            .in0(_gnd_net_),
            .in1(N__49894),
            .in2(N__53887),
            .in3(N__49888),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n412_adj_482 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17617 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17618 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_20_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_20_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_10_lut_LC_20_8_0  (
            .in0(_gnd_net_),
            .in1(N__49885),
            .in2(N__53939),
            .in3(N__49879),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n461_adj_470 ),
            .ltout(),
            .carryin(bfn_20_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_20_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_20_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_11_lut_LC_20_8_1  (
            .in0(_gnd_net_),
            .in1(N__53903),
            .in2(N__49876),
            .in3(N__49867),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n510_adj_458 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17619 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_20_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_20_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_12_lut_LC_20_8_2  (
            .in0(_gnd_net_),
            .in1(N__49864),
            .in2(N__53940),
            .in3(N__49858),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n559 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17620 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_20_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_20_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_13_lut_LC_20_8_3  (
            .in0(_gnd_net_),
            .in1(N__53907),
            .in2(N__49855),
            .in3(N__49996),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n608 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17621 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_20_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_20_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_14_lut_LC_20_8_4  (
            .in0(_gnd_net_),
            .in1(N__49993),
            .in2(N__53941),
            .in3(N__49987),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n657 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17622 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_20_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_20_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_15_lut_LC_20_8_5  (
            .in0(_gnd_net_),
            .in1(N__53911),
            .in2(N__49984),
            .in3(N__49975),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n706 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17623 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_20_8_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_20_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_20_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_567_16_lut_LC_20_8_6  (
            .in0(_gnd_net_),
            .in1(N__49972),
            .in2(N__49966),
            .in3(N__49945),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n762_adj_402 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17624 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_LUT4_0_LC_20_8_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_LUT4_0_LC_20_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_LUT4_0_LC_20_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_LUT4_0_LC_20_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49942),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n763_adj_386_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_20_9_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_20_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_2_lut_LC_20_9_0  (
            .in0(_gnd_net_),
            .in1(N__54176),
            .in2(N__54497),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n63 ),
            .ltout(),
            .carryin(bfn_20_9_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_20_9_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_20_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_3_lut_LC_20_9_1  (
            .in0(_gnd_net_),
            .in1(N__51772),
            .in2(N__54499),
            .in3(N__49939),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n112_adj_442 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17581 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_20_9_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_20_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_4_lut_LC_20_9_2  (
            .in0(_gnd_net_),
            .in1(N__54445),
            .in2(N__51754),
            .in3(N__49936),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n161_adj_395 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17582 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_20_9_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_20_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_5_lut_LC_20_9_3  (
            .in0(_gnd_net_),
            .in1(N__51997),
            .in2(N__54500),
            .in3(N__49933),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n210_adj_393 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17583 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_20_9_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_20_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_6_lut_LC_20_9_4  (
            .in0(_gnd_net_),
            .in1(N__54449),
            .in2(N__51979),
            .in3(N__50023),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n259_adj_391 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17584 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_20_9_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_20_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_7_lut_LC_20_9_5  (
            .in0(_gnd_net_),
            .in1(N__54437),
            .in2(N__51958),
            .in3(N__50020),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n308 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17585 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_20_9_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_20_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_8_lut_LC_20_9_6  (
            .in0(_gnd_net_),
            .in1(N__51937),
            .in2(N__54498),
            .in3(N__50017),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n357 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17586 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_20_9_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_20_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_9_lut_LC_20_9_7  (
            .in0(_gnd_net_),
            .in1(N__54441),
            .in2(N__51919),
            .in3(N__50014),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n406 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17587 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_20_10_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_20_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_10_lut_LC_20_10_0  (
            .in0(_gnd_net_),
            .in1(N__51898),
            .in2(N__54509),
            .in3(N__50011),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n455 ),
            .ltout(),
            .carryin(bfn_20_10_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_20_10_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_20_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_11_lut_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__51880),
            .in2(N__54510),
            .in3(N__50008),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n504_adj_467 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17589 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_20_10_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_20_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_12_lut_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__54469),
            .in2(N__52174),
            .in3(N__50005),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n553_adj_446 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17590 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_20_10_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_20_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_13_lut_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(N__52153),
            .in2(N__54511),
            .in3(N__50002),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n602_adj_355 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17591 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_20_10_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_20_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_14_lut_LC_20_10_4  (
            .in0(_gnd_net_),
            .in1(N__54473),
            .in2(N__52132),
            .in3(N__49999),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n651 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17592 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_20_10_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_20_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_15_lut_LC_20_10_5  (
            .in0(_gnd_net_),
            .in1(N__52111),
            .in2(N__54512),
            .in3(N__50161),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n700 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17593 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_20_10_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_20_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_565_16_lut_LC_20_10_6  (
            .in0(_gnd_net_),
            .in1(N__50158),
            .in2(N__52087),
            .in3(N__50137),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n754_adj_405 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17594 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_LUT4_0_LC_20_10_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_LUT4_0_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_LUT4_0_LC_20_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_LUT4_0_LC_20_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50134),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n755_adj_404_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_20_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_20_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_573_2_lut_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(N__60829),
            .in2(N__67409),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n87 ),
            .ltout(),
            .carryin(bfn_20_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_20_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_20_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_3_lut_LC_20_11_1  (
            .in0(_gnd_net_),
            .in1(N__50131),
            .in2(N__58899),
            .in3(N__50113),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n133_adj_388 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17897 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_20_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_20_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_4_lut_LC_20_11_2  (
            .in0(_gnd_net_),
            .in1(N__50110),
            .in2(N__54805),
            .in3(N__50092),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n182_adj_451 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17898 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17899 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_20_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_20_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_5_lut_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(N__50089),
            .in2(N__54534),
            .in3(N__50071),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n231_adj_387 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17899 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_20_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_20_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_6_lut_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__50068),
            .in2(N__54257),
            .in3(N__50050),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n280_adj_379 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17900 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_20_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_20_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_7_lut_LC_20_11_5  (
            .in0(_gnd_net_),
            .in1(N__53915),
            .in2(N__50047),
            .in3(N__50026),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n329_adj_439 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17901 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_20_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_20_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_8_lut_LC_20_11_6  (
            .in0(_gnd_net_),
            .in1(N__50317),
            .in2(N__53724),
            .in3(N__50299),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n378_adj_436 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17902 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_20_11_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_20_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_9_lut_LC_20_11_7  (
            .in0(_gnd_net_),
            .in1(N__50296),
            .in2(N__53369),
            .in3(N__50281),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n427_adj_432 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17903 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_20_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_20_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_10_lut_LC_20_12_0  (
            .in0(_gnd_net_),
            .in1(N__50278),
            .in2(N__53202),
            .in3(N__50260),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n476 ),
            .ltout(),
            .carryin(bfn_20_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_20_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_20_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_11_lut_LC_20_12_1  (
            .in0(_gnd_net_),
            .in1(N__50257),
            .in2(N__56214),
            .in3(N__50239),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n525 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17905 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_20_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_20_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_12_lut_LC_20_12_2  (
            .in0(_gnd_net_),
            .in1(N__50236),
            .in2(N__55940),
            .in3(N__50218),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n574 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17906 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_20_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_20_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_13_lut_LC_20_12_3  (
            .in0(_gnd_net_),
            .in1(N__50215),
            .in2(N__55718),
            .in3(N__50197),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n623 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17907 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_20_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_20_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_14_lut_LC_20_12_4  (
            .in0(_gnd_net_),
            .in1(N__50194),
            .in2(N__55365),
            .in3(N__50173),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n672 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17908 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_20_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_20_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_15_lut_LC_20_12_5  (
            .in0(_gnd_net_),
            .in1(N__55155),
            .in2(N__50170),
            .in3(N__50416),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n721 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17909 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_20_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_20_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_572_16_lut_LC_20_12_6  (
            .in0(_gnd_net_),
            .in1(N__54941),
            .in2(N__50413),
            .in3(N__50392),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n782 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17910 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_LUT4_0_LC_20_12_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_LUT4_0_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_LUT4_0_LC_20_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_LUT4_0_LC_20_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50389),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n783_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12703_3_lut_LC_20_13_5.C_ON=1'b0;
    defparam i12703_3_lut_LC_20_13_5.SEQ_MODE=4'b0000;
    defparam i12703_3_lut_LC_20_13_5.LUT_INIT=16'b0100010001100110;
    LogicCell40 i12703_3_lut_LC_20_13_5 (
            .in0(_gnd_net_),
            .in1(N__55001),
            .in2(_gnd_net_),
            .in3(N__50371),
            .lcout(n794_adj_2420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_20_13_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_20_13_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_i542_2_lut_LC_20_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51139),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_1_LC_20_14_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_1_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_1_LC_20_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_1_LC_20_14_0  (
            .in0(_gnd_net_),
            .in1(N__61200),
            .in2(N__61204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_14_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17505 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_2_lut_LC_20_14_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_2_lut_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_2_lut_LC_20_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_2_lut_LC_20_14_1  (
            .in0(_gnd_net_),
            .in1(N__51149),
            .in2(_gnd_net_),
            .in3(N__50326),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17505 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17506 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_3_lut_LC_20_14_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_3_lut_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_3_lut_LC_20_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_3_lut_LC_20_14_2  (
            .in0(_gnd_net_),
            .in1(N__58966),
            .in2(N__61177),
            .in3(N__50323),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17506 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17507 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_4_lut_LC_20_14_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_4_lut_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_4_lut_LC_20_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_4_lut_LC_20_14_3  (
            .in0(_gnd_net_),
            .in1(N__58948),
            .in2(N__52546),
            .in3(N__50320),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17507 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17508 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_5_lut_LC_20_14_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_5_lut_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_5_lut_LC_20_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_5_lut_LC_20_14_4  (
            .in0(_gnd_net_),
            .in1(N__52324),
            .in2(N__52528),
            .in3(N__50620),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17508 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17509 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_6_lut_LC_20_14_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_6_lut_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_6_lut_LC_20_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_6_lut_LC_20_14_5  (
            .in0(_gnd_net_),
            .in1(N__50617),
            .in2(N__52306),
            .in3(N__50608),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_19 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17509 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17510 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_7_lut_LC_20_14_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_7_lut_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_7_lut_LC_20_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_7_lut_LC_20_14_6  (
            .in0(_gnd_net_),
            .in1(N__52042),
            .in2(N__50605),
            .in3(N__50593),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17510 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17511 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_8_lut_LC_20_14_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_8_lut_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_8_lut_LC_20_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_8_lut_LC_20_14_7  (
            .in0(_gnd_net_),
            .in1(N__50590),
            .in2(N__52024),
            .in3(N__50581),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17511 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17512 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_9_lut_LC_20_15_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_9_lut_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_9_lut_LC_20_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_9_lut_LC_20_15_0  (
            .in0(_gnd_net_),
            .in1(N__50578),
            .in2(N__50566),
            .in3(N__50554),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_22 ),
            .ltout(),
            .carryin(bfn_20_15_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17513 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_10_lut_LC_20_15_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_10_lut_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_10_lut_LC_20_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_10_lut_LC_20_15_1  (
            .in0(_gnd_net_),
            .in1(N__50551),
            .in2(N__50536),
            .in3(N__50521),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_23 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17513 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17514 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_11_lut_LC_20_15_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_11_lut_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_11_lut_LC_20_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_11_lut_LC_20_15_2  (
            .in0(_gnd_net_),
            .in1(N__50518),
            .in2(N__50506),
            .in3(N__50491),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17514 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17515 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_12_lut_LC_20_15_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_12_lut_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_12_lut_LC_20_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_12_lut_LC_20_15_3  (
            .in0(_gnd_net_),
            .in1(N__50488),
            .in2(N__50470),
            .in3(N__50455),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17515 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17516 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_13_lut_LC_20_15_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_13_lut_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_13_lut_LC_20_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_13_lut_LC_20_15_4  (
            .in0(_gnd_net_),
            .in1(N__50452),
            .in2(N__50851),
            .in3(N__50830),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17516 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17517 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_14_lut_LC_20_15_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_14_lut_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_14_lut_LC_20_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_14_lut_LC_20_15_5  (
            .in0(_gnd_net_),
            .in1(N__50827),
            .in2(N__50812),
            .in3(N__50797),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17517 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_15_lut_LC_20_15_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_15_lut_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_15_lut_LC_20_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_15_lut_LC_20_15_6  (
            .in0(_gnd_net_),
            .in1(N__50794),
            .in2(N__50782),
            .in3(N__50764),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17518 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17519 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_16_lut_LC_20_15_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_16_lut_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_16_lut_LC_20_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_16_lut_LC_20_15_7  (
            .in0(_gnd_net_),
            .in1(N__50761),
            .in2(N__50752),
            .in3(N__50737),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17519 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17520 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_17_lut_LC_20_16_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_17_lut_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_17_lut_LC_20_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_3099_17_lut_LC_20_16_0  (
            .in0(_gnd_net_),
            .in1(N__50730),
            .in2(_gnd_net_),
            .in3(N__50716),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_269_LC_20_16_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_269_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_269_LC_20_16_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_269_LC_20_16_1  (
            .in0(N__50671),
            .in1(N__50664),
            .in2(N__50713),
            .in3(N__50626),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13205_2_lut_3_lut_LC_20_16_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13205_2_lut_3_lut_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13205_2_lut_3_lut_LC_20_16_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13205_2_lut_3_lut_LC_20_16_2  (
            .in0(N__59418),
            .in1(N__59295),
            .in2(_gnd_net_),
            .in3(N__51022),
            .lcout(\foc.qVoltage_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13212_2_lut_3_lut_LC_20_16_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13212_2_lut_3_lut_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13212_2_lut_3_lut_LC_20_16_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13212_2_lut_3_lut_LC_20_16_4  (
            .in0(N__59419),
            .in1(N__50712),
            .in2(_gnd_net_),
            .in3(N__59296),
            .lcout(\foc.qVoltage_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13215_2_lut_3_lut_LC_20_16_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13215_2_lut_3_lut_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13215_2_lut_3_lut_LC_20_16_6 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13215_2_lut_3_lut_LC_20_16_6  (
            .in0(N__50665),
            .in1(_gnd_net_),
            .in2(N__59440),
            .in3(N__59297),
            .lcout(\foc.qVoltage_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13206_2_lut_3_lut_LC_20_17_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13206_2_lut_3_lut_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13206_2_lut_3_lut_LC_20_17_0 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13206_2_lut_3_lut_LC_20_17_0  (
            .in0(N__51055),
            .in1(_gnd_net_),
            .in2(N__59315),
            .in3(N__59426),
            .lcout(),
            .ltout(\foc.qVoltage_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_266_LC_20_17_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_266_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_266_LC_20_17_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_266_LC_20_17_1  (
            .in0(N__51061),
            .in1(N__51054),
            .in2(N__51025),
            .in3(N__51021),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13209_2_lut_3_lut_LC_20_17_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13209_2_lut_3_lut_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13209_2_lut_3_lut_LC_20_17_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13209_2_lut_3_lut_LC_20_17_2  (
            .in0(N__59304),
            .in1(N__51208),
            .in2(_gnd_net_),
            .in3(N__59427),
            .lcout(\foc.qVoltage_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i27_3_lut_LC_20_17_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i27_3_lut_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i27_3_lut_LC_20_17_4 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i27_3_lut_LC_20_17_4  (
            .in0(N__59299),
            .in1(N__50983),
            .in2(_gnd_net_),
            .in3(N__59424),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_260_LC_20_17_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_260_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_260_LC_20_17_5 .LUT_INIT=16'b1010111011100100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_260_LC_20_17_5  (
            .in0(N__59425),
            .in1(N__59300),
            .in2(N__50959),
            .in3(N__52842),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13210_2_lut_3_lut_LC_20_17_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13210_2_lut_3_lut_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13210_2_lut_3_lut_LC_20_17_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13210_2_lut_3_lut_LC_20_17_6  (
            .in0(N__59305),
            .in1(N__50932),
            .in2(_gnd_net_),
            .in3(N__59428),
            .lcout(),
            .ltout(\foc.qVoltage_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i18_2_lut_LC_20_17_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i18_2_lut_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i18_2_lut_LC_20_17_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i18_2_lut_LC_20_17_7  (
            .in0(N__50931),
            .in1(_gnd_net_),
            .in2(N__50899),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6572_2_lut_LC_20_18_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6572_2_lut_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6572_2_lut_LC_20_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i6572_2_lut_LC_20_18_1  (
            .in0(N__55033),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51160),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n8265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_261_LC_20_18_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_261_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_261_LC_20_18_3 .LUT_INIT=16'b1011101001110010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_261_LC_20_18_3  (
            .in0(N__59442),
            .in1(N__50890),
            .in2(N__59326),
            .in3(N__50881),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20586_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_265_LC_20_18_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_265_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_265_LC_20_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_265_LC_20_18_4  (
            .in0(N__51235),
            .in1(N__51229),
            .in2(N__51223),
            .in3(N__51220),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_270_LC_20_18_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_270_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_270_LC_20_18_5 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_270_LC_20_18_5  (
            .in0(N__51214),
            .in1(N__51204),
            .in2(N__51169),
            .in3(N__51166),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6570_2_lut_LC_20_18_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6570_2_lut_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i6570_2_lut_LC_20_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i6570_2_lut_LC_20_18_7  (
            .in0(N__55032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51159),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n738_adj_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i20_LC_20_19_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i20_LC_20_19_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i20_LC_20_19_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i20_LC_20_19_2  (
            .in0(N__56463),
            .in1(N__56342),
            .in2(_gnd_net_),
            .in3(N__57561),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62106),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_20_19_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_20_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.paramCurrentControlP_15__I_0_i37_2_lut_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51078),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i27_LC_20_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i27_LC_20_20_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i27_LC_20_20_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i27_LC_20_20_0  (
            .in0(N__56441),
            .in1(N__56308),
            .in2(_gnd_net_),
            .in3(N__57987),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62108),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i24_LC_20_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i24_LC_20_20_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i24_LC_20_20_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i24_LC_20_20_1  (
            .in0(N__56306),
            .in1(N__56440),
            .in2(_gnd_net_),
            .in3(N__58170),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62108),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i29_LC_20_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i29_LC_20_20_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i29_LC_20_20_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i29_LC_20_20_2  (
            .in0(N__56442),
            .in1(N__56309),
            .in2(_gnd_net_),
            .in3(N__57887),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62108),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_289_LC_20_20_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_289_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_289_LC_20_20_3 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_289_LC_20_20_3  (
            .in0(N__57562),
            .in1(N__51274),
            .in2(N__57424),
            .in3(N__57492),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_290_LC_20_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_290_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_290_LC_20_20_4 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_290_LC_20_20_4  (
            .in0(N__58171),
            .in1(N__58240),
            .in2(N__51265),
            .in3(N__58111),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i790_4_lut_LC_20_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i790_4_lut_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i790_4_lut_LC_20_20_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i790_4_lut_LC_20_20_5  (
            .in0(N__57988),
            .in1(N__57940),
            .in2(N__51262),
            .in3(N__58042),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_293_LC_20_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_293_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_293_LC_20_20_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_293_LC_20_20_6  (
            .in0(N__58487),
            .in1(N__57888),
            .in2(N__51259),
            .in3(N__58369),
            .lcout(Saturate_out1_31__N_266_adj_2417),
            .ltout(Saturate_out1_31__N_266_adj_2417_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i26_LC_20_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i26_LC_20_20_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i26_LC_20_20_7 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i26_LC_20_20_7  (
            .in0(N__56307),
            .in1(_gnd_net_),
            .in2(N__51256),
            .in3(N__58041),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62108),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i21_LC_20_21_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i21_LC_20_21_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i21_LC_20_21_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i21_LC_20_21_0  (
            .in0(N__56458),
            .in1(N__56298),
            .in2(_gnd_net_),
            .in3(N__57493),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i19_LC_20_21_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i19_LC_20_21_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i19_LC_20_21_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i19_LC_20_21_1  (
            .in0(N__57640),
            .in1(N__56297),
            .in2(_gnd_net_),
            .in3(N__56457),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i2_LC_20_21_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i2_LC_20_21_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i2_LC_20_21_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i2_LC_20_21_2  (
            .in0(N__56460),
            .in1(N__60076),
            .in2(_gnd_net_),
            .in3(N__56300),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i62_4_lut_LC_20_21_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i62_4_lut_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i62_4_lut_LC_20_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.equal_13244_i62_4_lut_LC_20_21_3  (
            .in0(N__51253),
            .in1(N__59122),
            .in2(N__52957),
            .in3(N__51244),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Not_Equal_relop1_N_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_283_LC_20_21_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_283_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_283_LC_20_21_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_283_LC_20_21_4  (
            .in0(N__58368),
            .in1(N__58489),
            .in2(N__57889),
            .in3(N__56608),
            .lcout(Saturate_out1_31__N_267_adj_2418),
            .ltout(Saturate_out1_31__N_267_adj_2418_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i6_LC_20_21_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i6_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i6_LC_20_21_5 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i6_LC_20_21_5  (
            .in0(N__62671),
            .in1(_gnd_net_),
            .in2(N__51286),
            .in3(N__56462),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i30_LC_20_21_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i30_LC_20_21_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i30_LC_20_21_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i30_LC_20_21_6  (
            .in0(N__56461),
            .in1(N__56301),
            .in2(_gnd_net_),
            .in3(N__58488),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i23_LC_20_21_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i23_LC_20_21_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i23_LC_20_21_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i23_LC_20_21_7  (
            .in0(N__56299),
            .in1(N__58239),
            .in2(_gnd_net_),
            .in3(N__56459),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62113),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i12_LC_20_22_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i12_LC_20_22_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i12_LC_20_22_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i12_LC_20_22_0  (
            .in0(N__56481),
            .in1(N__56302),
            .in2(_gnd_net_),
            .in3(N__60327),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62118),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i4_LC_20_22_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i4_LC_20_22_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i4_LC_20_22_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i4_LC_20_22_1  (
            .in0(N__56304),
            .in1(N__60112),
            .in2(_gnd_net_),
            .in3(N__56483),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62118),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i772_4_lut_LC_20_22_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i772_4_lut_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i772_4_lut_LC_20_22_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i772_4_lut_LC_20_22_2  (
            .in0(N__62647),
            .in1(N__60411),
            .in2(N__60354),
            .in3(N__60382),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n22_adj_762_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_286_LC_20_22_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_286_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_286_LC_20_22_3 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_286_LC_20_22_3  (
            .in0(N__60328),
            .in1(N__60310),
            .in2(N__51283),
            .in3(N__60285),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20694_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_287_LC_20_22_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_287_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_287_LC_20_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_287_LC_20_22_4  (
            .in0(N__60222),
            .in1(N__60189),
            .in2(N__51280),
            .in3(N__60258),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_288_LC_20_22_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_288_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_288_LC_20_22_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_288_LC_20_22_5  (
            .in0(N__57786),
            .in1(N__57639),
            .in2(N__51277),
            .in3(N__57717),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i8_LC_20_22_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i8_LC_20_22_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i8_LC_20_22_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i8_LC_20_22_6  (
            .in0(N__56484),
            .in1(N__56305),
            .in2(_gnd_net_),
            .in3(N__60381),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62118),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i13_LC_20_22_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i13_LC_20_22_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i13_LC_20_22_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i13_LC_20_22_7  (
            .in0(N__56303),
            .in1(N__60309),
            .in2(_gnd_net_),
            .in3(N__56482),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62118),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_20_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_20_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_2_lut_LC_20_23_0  (
            .in0(_gnd_net_),
            .in1(N__64712),
            .in2(N__64887),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n63 ),
            .ltout(),
            .carryin(bfn_20_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18204 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_20_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_20_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_3_lut_LC_20_23_1  (
            .in0(_gnd_net_),
            .in1(N__64454),
            .in2(N__51361),
            .in3(N__51343),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n109 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18204 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18205 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_20_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_20_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_20_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_4_lut_LC_20_23_2  (
            .in0(_gnd_net_),
            .in1(N__51544),
            .in2(N__64178),
            .in3(N__51334),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n158 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18205 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18206 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_20_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_20_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_5_lut_LC_20_23_3  (
            .in0(_gnd_net_),
            .in1(N__51532),
            .in2(N__63888),
            .in3(N__51325),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n207 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18206 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18207 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_20_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_20_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_6_lut_LC_20_23_4  (
            .in0(_gnd_net_),
            .in1(N__51520),
            .in2(N__63631),
            .in3(N__51316),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n256 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18207 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18208 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_20_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_20_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_7_lut_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(N__51508),
            .in2(N__63378),
            .in3(N__51307),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n305 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18208 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18209 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_20_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_20_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_8_lut_LC_20_23_6  (
            .in0(_gnd_net_),
            .in1(N__62938),
            .in2(N__51496),
            .in3(N__51298),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n354 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18209 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18210 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_20_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_20_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_9_lut_LC_20_23_7  (
            .in0(_gnd_net_),
            .in1(N__66760),
            .in2(N__51481),
            .in3(N__51457),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n403 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18210 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18211 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_20_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_20_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_10_lut_LC_20_24_0  (
            .in0(_gnd_net_),
            .in1(N__51466),
            .in2(N__66599),
            .in3(N__51448),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n452 ),
            .ltout(),
            .carryin(bfn_20_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_20_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_20_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_11_lut_LC_20_24_1  (
            .in0(_gnd_net_),
            .in1(N__51670),
            .in2(N__66286),
            .in3(N__51439),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n501 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18212 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18213 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_20_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_20_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_12_lut_LC_20_24_2  (
            .in0(_gnd_net_),
            .in1(N__51658),
            .in2(N__66091),
            .in3(N__51430),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n550 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18213 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18214 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_20_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_20_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_13_lut_LC_20_24_3  (
            .in0(_gnd_net_),
            .in1(N__51646),
            .in2(N__65830),
            .in3(N__51421),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n599 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18214 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18215 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_20_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_20_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_14_lut_LC_20_24_4  (
            .in0(_gnd_net_),
            .in1(N__65595),
            .in2(N__51634),
            .in3(N__51409),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n648 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18215 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_20_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_20_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_15_lut_LC_20_24_5  (
            .in0(_gnd_net_),
            .in1(N__65348),
            .in2(N__51619),
            .in3(N__51397),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n697 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18216 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18217 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_20_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_20_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_564_16_lut_LC_20_24_6  (
            .in0(_gnd_net_),
            .in1(N__65139),
            .in2(N__51601),
            .in3(N__51382),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n750 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18217 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_LUT4_0_LC_20_24_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_LUT4_0_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_LUT4_0_LC_20_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_LUT4_0_LC_20_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51379),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n751_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_20_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_20_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_2_lut_LC_20_25_0  (
            .in0(_gnd_net_),
            .in1(N__64713),
            .in2(N__64900),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n66 ),
            .ltout(),
            .carryin(bfn_20_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18219 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_20_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_20_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_20_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_3_lut_LC_20_25_1  (
            .in0(_gnd_net_),
            .in1(N__64478),
            .in2(N__51553),
            .in3(N__51535),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n112 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18219 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18220 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_20_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_20_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_4_lut_LC_20_25_2  (
            .in0(_gnd_net_),
            .in1(N__60544),
            .in2(N__64230),
            .in3(N__51523),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n161 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18220 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18221 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_20_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_20_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_5_lut_LC_20_25_3  (
            .in0(_gnd_net_),
            .in1(N__60532),
            .in2(N__63963),
            .in3(N__51511),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n210 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18221 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18222 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_20_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_20_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_6_lut_LC_20_25_4  (
            .in0(_gnd_net_),
            .in1(N__60520),
            .in2(N__63647),
            .in3(N__51499),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n259 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18222 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18223 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_20_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_20_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_7_lut_LC_20_25_5  (
            .in0(_gnd_net_),
            .in1(N__60508),
            .in2(N__63382),
            .in3(N__51484),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n308 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18223 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18224 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_20_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_20_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_20_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_8_lut_LC_20_25_6  (
            .in0(_gnd_net_),
            .in1(N__63093),
            .in2(N__60496),
            .in3(N__51469),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n357 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18224 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18225 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_20_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_20_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_9_lut_LC_20_25_7  (
            .in0(_gnd_net_),
            .in1(N__66782),
            .in2(N__60481),
            .in3(N__51460),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n406 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18225 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18226 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_20_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_20_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_10_lut_LC_20_26_0  (
            .in0(_gnd_net_),
            .in1(N__60466),
            .in2(N__66600),
            .in3(N__51661),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n455 ),
            .ltout(),
            .carryin(bfn_20_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18227 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_20_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_20_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_20_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_11_lut_LC_20_26_1  (
            .in0(_gnd_net_),
            .in1(N__60673),
            .in2(N__66348),
            .in3(N__51649),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n504 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18227 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18228 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_20_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_20_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_12_lut_LC_20_26_2  (
            .in0(_gnd_net_),
            .in1(N__60661),
            .in2(N__66070),
            .in3(N__51637),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n553 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18228 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18229 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_20_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_20_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_20_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_13_lut_LC_20_26_3  (
            .in0(_gnd_net_),
            .in1(N__60649),
            .in2(N__65839),
            .in3(N__51622),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n602 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18229 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18230 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_20_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_20_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_20_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_14_lut_LC_20_26_4  (
            .in0(_gnd_net_),
            .in1(N__60637),
            .in2(N__65600),
            .in3(N__51604),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n651 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18230 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18231 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_20_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_20_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_20_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_15_lut_LC_20_26_5  (
            .in0(_gnd_net_),
            .in1(N__65352),
            .in2(N__60625),
            .in3(N__51589),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n700 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18231 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18232 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_20_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_20_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_20_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_565_16_lut_LC_20_26_6  (
            .in0(_gnd_net_),
            .in1(N__65170),
            .in2(N__60610),
            .in3(N__51574),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n754 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18232 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_LUT4_0_LC_20_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_LUT4_0_LC_20_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_LUT4_0_LC_20_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_LUT4_0_LC_20_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51571),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n755_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_20_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_20_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_20_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_572_2_lut_LC_20_28_0  (
            .in0(_gnd_net_),
            .in1(N__64888),
            .in2(N__64748),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n84 ),
            .ltout(),
            .carryin(bfn_20_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18309 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_20_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_20_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_20_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_3_lut_LC_20_28_1  (
            .in0(_gnd_net_),
            .in1(N__51742),
            .in2(N__64488),
            .in3(N__51736),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n130 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18309 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18310 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_20_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_20_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_20_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_4_lut_LC_20_28_2  (
            .in0(_gnd_net_),
            .in1(N__51733),
            .in2(N__64232),
            .in3(N__51727),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n179 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18310 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18311 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_20_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_20_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_20_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_5_lut_LC_20_28_3  (
            .in0(_gnd_net_),
            .in1(N__51724),
            .in2(N__63982),
            .in3(N__51718),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n228 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18311 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18312 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_20_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_20_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_20_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_6_lut_LC_20_28_4  (
            .in0(_gnd_net_),
            .in1(N__51715),
            .in2(N__63655),
            .in3(N__51709),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n277 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18312 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18313 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_20_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_20_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_20_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_7_lut_LC_20_28_5  (
            .in0(_gnd_net_),
            .in1(N__51706),
            .in2(N__63385),
            .in3(N__51700),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n326_adj_588 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18313 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18314 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_20_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_20_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_20_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_8_lut_LC_20_28_6  (
            .in0(_gnd_net_),
            .in1(N__51697),
            .in2(N__63095),
            .in3(N__51691),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n375_adj_587 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18314 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18315 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_20_28_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_20_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_20_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_9_lut_LC_20_28_7  (
            .in0(_gnd_net_),
            .in1(N__51688),
            .in2(N__66921),
            .in3(N__51682),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n424_adj_586 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18315 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18316 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_20_29_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_20_29_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_20_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_10_lut_LC_20_29_0  (
            .in0(_gnd_net_),
            .in1(N__51679),
            .in2(N__66625),
            .in3(N__51673),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n473_adj_585 ),
            .ltout(),
            .carryin(bfn_20_29_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18317 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_20_29_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_20_29_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_20_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_11_lut_LC_20_29_1  (
            .in0(_gnd_net_),
            .in1(N__51868),
            .in2(N__66346),
            .in3(N__51862),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n522_adj_584 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18317 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18318 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_20_29_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_20_29_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_20_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_12_lut_LC_20_29_2  (
            .in0(_gnd_net_),
            .in1(N__51859),
            .in2(N__66093),
            .in3(N__51853),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n571 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18318 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18319 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_20_29_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_20_29_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_20_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_13_lut_LC_20_29_3  (
            .in0(_gnd_net_),
            .in1(N__51850),
            .in2(N__65831),
            .in3(N__51844),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n620 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18319 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18320 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_20_29_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_20_29_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_20_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_14_lut_LC_20_29_4  (
            .in0(_gnd_net_),
            .in1(N__51841),
            .in2(N__65601),
            .in3(N__51835),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n669 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18320 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18321 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_20_29_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_20_29_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_20_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_15_lut_LC_20_29_5  (
            .in0(_gnd_net_),
            .in1(N__65361),
            .in2(N__51832),
            .in3(N__51823),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n718 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18321 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18322 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_20_29_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_20_29_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_20_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_16_lut_LC_20_29_6  (
            .in0(_gnd_net_),
            .in1(N__65192),
            .in2(N__51820),
            .in3(N__51796),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n778 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18322 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_LUT4_0_LC_20_29_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_LUT4_0_LC_20_29_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_LUT4_0_LC_20_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_LUT4_0_LC_20_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51793),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n779_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_21_7_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_21_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_2_lut_LC_21_7_0  (
            .in0(_gnd_net_),
            .in1(N__53888),
            .in2(N__54135),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n66 ),
            .ltout(),
            .carryin(bfn_21_7_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_21_7_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_21_7_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_21_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_3_lut_LC_21_7_1  (
            .in0(_gnd_net_),
            .in1(N__54084),
            .in2(N__51763),
            .in3(N__52009),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n115_adj_488 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17596 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_21_7_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_21_7_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_21_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_4_lut_LC_21_7_2  (
            .in0(_gnd_net_),
            .in1(N__54138),
            .in2(N__52006),
            .in3(N__51988),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n164_adj_466 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17597 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_21_7_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_21_7_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_21_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_5_lut_LC_21_7_3  (
            .in0(_gnd_net_),
            .in1(N__51985),
            .in2(N__54193),
            .in3(N__51967),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n213_adj_445 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17598 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17599 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_21_7_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_21_7_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_21_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_6_lut_LC_21_7_4  (
            .in0(_gnd_net_),
            .in1(N__51964),
            .in2(N__54136),
            .in3(N__51946),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n262 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17599 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_21_7_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_21_7_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_21_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_7_lut_LC_21_7_5  (
            .in0(_gnd_net_),
            .in1(N__51943),
            .in2(N__54194),
            .in3(N__51928),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n311 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17600 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17601 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_21_7_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_21_7_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_21_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_8_lut_LC_21_7_6  (
            .in0(_gnd_net_),
            .in1(N__51925),
            .in2(N__54137),
            .in3(N__51907),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n360_adj_484 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17601 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_21_7_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_21_7_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_21_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_9_lut_LC_21_7_7  (
            .in0(_gnd_net_),
            .in1(N__51904),
            .in2(N__54195),
            .in3(N__51889),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n409_adj_483 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17602 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_21_8_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_21_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_10_lut_LC_21_8_0  (
            .in0(_gnd_net_),
            .in1(N__51886),
            .in2(N__54252),
            .in3(N__51871),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n458_adj_468 ),
            .ltout(),
            .carryin(bfn_21_8_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17604 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_21_8_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_21_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_11_lut_LC_21_8_1  (
            .in0(_gnd_net_),
            .in1(N__54224),
            .in2(N__52183),
            .in3(N__52162),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n507_adj_447 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17604 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17605 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_21_8_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_21_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_12_lut_LC_21_8_2  (
            .in0(_gnd_net_),
            .in1(N__52159),
            .in2(N__54253),
            .in3(N__52144),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n556 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17605 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_21_8_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_21_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_13_lut_LC_21_8_3  (
            .in0(_gnd_net_),
            .in1(N__54228),
            .in2(N__52141),
            .in3(N__52120),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n605 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17606 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_21_8_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_21_8_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_21_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_14_lut_LC_21_8_4  (
            .in0(_gnd_net_),
            .in1(N__52117),
            .in2(N__54254),
            .in3(N__52099),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n654 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17607 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_21_8_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_21_8_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_21_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_15_lut_LC_21_8_5  (
            .in0(_gnd_net_),
            .in1(N__54232),
            .in2(N__52096),
            .in3(N__52072),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n703 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17608 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17609 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_21_8_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_21_8_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_21_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_566_16_lut_LC_21_8_6  (
            .in0(_gnd_net_),
            .in1(N__52069),
            .in2(N__52051),
            .in3(N__52030),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n758_adj_403 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17609 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_LUT4_0_LC_21_8_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_LUT4_0_LC_21_8_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_LUT4_0_LC_21_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_LUT4_0_LC_21_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52027),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n759_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_21_9_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_21_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_2_lut_LC_21_9_0  (
            .in0(_gnd_net_),
            .in1(N__54450),
            .in2(N__54796),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n60_adj_495 ),
            .ltout(),
            .carryin(bfn_21_9_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17566 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_21_9_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_21_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_3_lut_LC_21_9_1  (
            .in0(_gnd_net_),
            .in1(N__54750),
            .in2(N__52276),
            .in3(N__52267),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n109 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17566 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17567 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_21_9_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_21_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_4_lut_LC_21_9_2  (
            .in0(_gnd_net_),
            .in1(N__52264),
            .in2(N__54797),
            .in3(N__52258),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n158 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17567 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_21_9_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_21_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_5_lut_LC_21_9_3  (
            .in0(_gnd_net_),
            .in1(N__52255),
            .in2(N__54800),
            .in3(N__52249),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n207_adj_394 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17568 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_21_9_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_21_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_6_lut_LC_21_9_4  (
            .in0(_gnd_net_),
            .in1(N__52246),
            .in2(N__54798),
            .in3(N__52240),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n256_adj_392 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17569 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_21_9_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_21_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_7_lut_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(N__54757),
            .in2(N__52237),
            .in3(N__52228),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n305_adj_390 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17570 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_21_9_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_21_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_8_lut_LC_21_9_6  (
            .in0(_gnd_net_),
            .in1(N__52225),
            .in2(N__54799),
            .in3(N__52219),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n354 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17571 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_21_9_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_21_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_9_lut_LC_21_9_7  (
            .in0(_gnd_net_),
            .in1(N__54761),
            .in2(N__52216),
            .in3(N__52207),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n403 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17572 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_21_10_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_21_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_10_lut_LC_21_10_0  (
            .in0(_gnd_net_),
            .in1(N__52204),
            .in2(N__54768),
            .in3(N__52198),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n452 ),
            .ltout(),
            .carryin(bfn_21_10_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_21_10_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_21_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_11_lut_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(N__54705),
            .in2(N__52195),
            .in3(N__52186),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n501_adj_481 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17574 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_21_10_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_21_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_12_lut_LC_21_10_2  (
            .in0(_gnd_net_),
            .in1(N__52393),
            .in2(N__54769),
            .in3(N__52387),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n550_adj_441 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17575 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_21_10_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_21_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_13_lut_LC_21_10_3  (
            .in0(_gnd_net_),
            .in1(N__54709),
            .in2(N__52384),
            .in3(N__52375),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n599_adj_376 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17576 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_21_10_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_21_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_14_lut_LC_21_10_4  (
            .in0(_gnd_net_),
            .in1(N__52372),
            .in2(N__54770),
            .in3(N__52366),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n648 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17577 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_21_10_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_21_10_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_21_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_15_lut_LC_21_10_5  (
            .in0(_gnd_net_),
            .in1(N__54713),
            .in2(N__52363),
            .in3(N__52354),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n697_adj_444 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17578 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_21_10_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_21_10_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_21_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_564_16_lut_LC_21_10_6  (
            .in0(_gnd_net_),
            .in1(N__52351),
            .in2(N__52333),
            .in3(N__52312),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n750_adj_407 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17579 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_LUT4_0_LC_21_10_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_LUT4_0_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_LUT4_0_LC_21_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_LUT4_0_LC_21_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52309),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n751_adj_406_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_21_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_21_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_2_lut_LC_21_11_0  (
            .in0(_gnd_net_),
            .in1(N__54801),
            .in2(N__58900),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n57_adj_491 ),
            .ltout(),
            .carryin(bfn_21_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17551 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_21_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_21_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_3_lut_LC_21_11_1  (
            .in0(_gnd_net_),
            .in1(N__58852),
            .in2(N__52291),
            .in3(N__52279),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n106_adj_509 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17551 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17552 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_21_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_21_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_4_lut_LC_21_11_2  (
            .in0(_gnd_net_),
            .in1(N__52510),
            .in2(N__58901),
            .in3(N__52501),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n155 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17552 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_21_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_21_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_5_lut_LC_21_11_3  (
            .in0(_gnd_net_),
            .in1(N__58856),
            .in2(N__52498),
            .in3(N__52486),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n204 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17553 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_21_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_21_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_6_lut_LC_21_11_4  (
            .in0(_gnd_net_),
            .in1(N__52483),
            .in2(N__58902),
            .in3(N__52474),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n253_adj_464 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17554 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_21_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_21_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_7_lut_LC_21_11_5  (
            .in0(_gnd_net_),
            .in1(N__58860),
            .in2(N__52471),
            .in3(N__52459),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n302 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17555 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_21_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_21_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_8_lut_LC_21_11_6  (
            .in0(_gnd_net_),
            .in1(N__52456),
            .in2(N__58903),
            .in3(N__52447),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n351_adj_396 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17556 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_21_11_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_21_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_9_lut_LC_21_11_7  (
            .in0(_gnd_net_),
            .in1(N__58864),
            .in2(N__52444),
            .in3(N__52432),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n400 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17557 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_21_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_21_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_10_lut_LC_21_12_0  (
            .in0(_gnd_net_),
            .in1(N__52429),
            .in2(N__58909),
            .in3(N__52420),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n449 ),
            .ltout(),
            .carryin(bfn_21_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_21_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_21_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_11_lut_LC_21_12_1  (
            .in0(_gnd_net_),
            .in1(N__58887),
            .in2(N__52417),
            .in3(N__52405),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n498 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17559 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_21_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_21_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_12_lut_LC_21_12_2  (
            .in0(_gnd_net_),
            .in1(N__52402),
            .in2(N__58910),
            .in3(N__52624),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n547 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17560 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17561 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_21_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_21_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_13_lut_LC_21_12_3  (
            .in0(_gnd_net_),
            .in1(N__58891),
            .in2(N__52621),
            .in3(N__52609),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n596 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17561 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17562 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_21_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_21_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_14_lut_LC_21_12_4  (
            .in0(_gnd_net_),
            .in1(N__52606),
            .in2(N__58911),
            .in3(N__52597),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n645 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17562 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17563 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_21_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_21_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_15_lut_LC_21_12_5  (
            .in0(_gnd_net_),
            .in1(N__58895),
            .in2(N__52594),
            .in3(N__52582),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n694 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17563 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17564 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_21_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_21_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_563_16_lut_LC_21_12_6  (
            .in0(_gnd_net_),
            .in1(N__52579),
            .in2(N__52558),
            .in3(N__52534),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n746_adj_409 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17564 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_LUT4_0_LC_21_12_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_LUT4_0_LC_21_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_LUT4_0_LC_21_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_LUT4_0_LC_21_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52531),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n747_adj_408_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13161_2_lut_3_lut_LC_21_13_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13161_2_lut_3_lut_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13161_2_lut_3_lut_LC_21_13_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13161_2_lut_3_lut_LC_21_13_6  (
            .in0(N__61389),
            .in1(N__67618),
            .in2(_gnd_net_),
            .in3(N__61454),
            .lcout(),
            .ltout(\foc.dVoltage_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_119_LC_21_13_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_119_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_119_LC_21_13_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_119_LC_21_13_7  (
            .in0(N__67617),
            .in1(N__67978),
            .in2(N__52513),
            .in3(N__59071),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13174_2_lut_3_lut_LC_21_14_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13174_2_lut_3_lut_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13174_2_lut_3_lut_LC_21_14_0 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13174_2_lut_3_lut_LC_21_14_0  (
            .in0(N__68608),
            .in1(_gnd_net_),
            .in2(N__61479),
            .in3(N__61377),
            .lcout(\foc.dVoltage_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13168_2_lut_3_lut_LC_21_14_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13168_2_lut_3_lut_LC_21_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13168_2_lut_3_lut_LC_21_14_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13168_2_lut_3_lut_LC_21_14_1  (
            .in0(N__61375),
            .in1(N__67899),
            .in2(_gnd_net_),
            .in3(N__61462),
            .lcout(\foc.dVoltage_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13169_2_lut_3_lut_LC_21_14_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13169_2_lut_3_lut_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13169_2_lut_3_lut_LC_21_14_2 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13169_2_lut_3_lut_LC_21_14_2  (
            .in0(N__68944),
            .in1(_gnd_net_),
            .in2(N__61478),
            .in3(N__61376),
            .lcout(\foc.dVoltage_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_118_LC_21_14_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_118_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_118_LC_21_14_3 .LUT_INIT=16'b1100111011100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_118_LC_21_14_3  (
            .in0(N__61374),
            .in1(N__61461),
            .in2(N__68557),
            .in3(N__69208),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_121_LC_21_14_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_121_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_121_LC_21_14_4 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_121_LC_21_14_4  (
            .in0(N__68607),
            .in1(N__59104),
            .in2(N__52678),
            .in3(N__52675),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_124_LC_21_14_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_124_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_124_LC_21_14_5 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_124_LC_21_14_5  (
            .in0(N__59080),
            .in1(N__68943),
            .in2(N__52669),
            .in3(N__52666),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_127_LC_21_14_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_127_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_127_LC_21_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_127_LC_21_14_6  (
            .in0(N__59218),
            .in1(N__61501),
            .in2(N__52660),
            .in3(N__59203),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19727_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i62_4_lut_LC_21_14_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i62_4_lut_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i62_4_lut_LC_21_14_7 .LUT_INIT=16'b0000110000001101;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i62_4_lut_LC_21_14_7  (
            .in0(N__61373),
            .in1(N__61306),
            .in2(N__52657),
            .in3(N__61460),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Not_Equal_relop1_N_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13207_2_lut_3_lut_LC_21_15_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13207_2_lut_3_lut_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13207_2_lut_3_lut_LC_21_15_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13207_2_lut_3_lut_LC_21_15_4  (
            .in0(N__52651),
            .in1(N__59298),
            .in2(_gnd_net_),
            .in3(N__59423),
            .lcout(),
            .ltout(\foc.qVoltage_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_LC_21_15_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_LC_21_15_5 .LUT_INIT=16'b1010111111111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_3_lut_LC_21_15_5  (
            .in0(N__52909),
            .in1(_gnd_net_),
            .in2(N__52654),
            .in3(N__52650),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_267_LC_21_15_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_267_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_267_LC_21_15_6 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_267_LC_21_15_6  (
            .in0(N__52684),
            .in1(N__52726),
            .in2(N__52960),
            .in3(N__59161),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_262_LC_21_16_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_262_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_262_LC_21_16_1 .LUT_INIT=16'b1111101001001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_262_LC_21_16_1  (
            .in0(N__52874),
            .in1(N__59292),
            .in2(N__52942),
            .in3(N__59415),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1223_rep_3_4_lut_LC_21_16_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1223_rep_3_4_lut_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1223_rep_3_4_lut_LC_21_16_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i1223_rep_3_4_lut_LC_21_16_2  (
            .in0(N__52903),
            .in1(N__52875),
            .in2(N__52857),
            .in3(N__52824),
            .lcout(\foc.Out_31__N_333 ),
            .ltout(\foc.Out_31__N_333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13211_2_lut_3_lut_LC_21_16_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13211_2_lut_3_lut_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13211_2_lut_3_lut_LC_21_16_3 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13211_2_lut_3_lut_LC_21_16_3  (
            .in0(N__52795),
            .in1(_gnd_net_),
            .in2(N__52891),
            .in3(N__59416),
            .lcout(\foc.qVoltage_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i12830_4_lut_LC_21_16_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i12830_4_lut_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i12830_4_lut_LC_21_16_4 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i12830_4_lut_LC_21_16_4  (
            .in0(N__52888),
            .in1(N__52876),
            .in2(N__52858),
            .in3(N__52825),
            .lcout(\foc.Out_31__N_332 ),
            .ltout(\foc.Out_31__N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13216_2_lut_3_lut_LC_21_16_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13216_2_lut_3_lut_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13216_2_lut_3_lut_LC_21_16_5 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13216_2_lut_3_lut_LC_21_16_5  (
            .in0(N__52756),
            .in1(_gnd_net_),
            .in2(N__52804),
            .in3(N__59293),
            .lcout(),
            .ltout(\foc.qVoltage_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_264_LC_21_16_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_264_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_264_LC_21_16_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_264_LC_21_16_6  (
            .in0(N__52801),
            .in1(N__52794),
            .in2(N__52759),
            .in3(N__52755),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13217_2_lut_3_lut_LC_21_16_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13217_2_lut_3_lut_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13217_2_lut_3_lut_LC_21_16_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13217_2_lut_3_lut_LC_21_16_7  (
            .in0(N__52722),
            .in1(N__59294),
            .in2(_gnd_net_),
            .in3(N__59417),
            .lcout(\foc.qVoltage_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_17_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_17_0  (
            .in0(_gnd_net_),
            .in1(N__60902),
            .in2(N__67467),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n57 ),
            .ltout(),
            .carryin(bfn_21_17_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_17_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_17_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_17_1  (
            .in0(N__55444),
            .in1(N__54826),
            .in2(N__58915),
            .in3(N__54820),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_4 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17736 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_17_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_17_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_17_2  (
            .in0(N__55448),
            .in1(N__54817),
            .in2(N__54568),
            .in3(N__54553),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_5 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17737 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_17_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_17_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_17_3  (
            .in0(N__55445),
            .in1(N__54550),
            .in2(N__54538),
            .in3(N__54286),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_6 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17738 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_17_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_17_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_17_4  (
            .in0(N__55449),
            .in1(N__54283),
            .in2(N__54271),
            .in3(N__54016),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_7 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17739 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_17_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_17_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_17_5  (
            .in0(N__55446),
            .in1(N__54013),
            .in2(N__53999),
            .in3(N__53743),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_8 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17740 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_17_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_17_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_17_6  (
            .in0(N__55450),
            .in1(N__53740),
            .in2(N__53723),
            .in3(N__53494),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_9 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17741 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_17_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_17_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_17_7  (
            .in0(N__55447),
            .in1(N__53491),
            .in2(N__53478),
            .in3(N__53227),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_10 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17742 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_18_0  (
            .in0(N__55451),
            .in1(N__53224),
            .in2(N__53136),
            .in3(N__52963),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_11 ),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_18_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_18_1  (
            .in0(N__55454),
            .in1(N__56227),
            .in2(N__56215),
            .in3(N__55981),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_12 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17744 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_18_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_18_2  (
            .in0(N__55452),
            .in1(N__55978),
            .in2(N__55964),
            .in3(N__55753),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17745 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_18_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_18_3  (
            .in0(N__55455),
            .in1(N__55750),
            .in2(N__55737),
            .in3(N__55522),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_14 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17746 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_18_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_18_4  (
            .in0(N__55453),
            .in1(N__55390),
            .in2(N__55377),
            .in3(N__55189),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Switch_out1_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17747 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__55179),
            .in2(N__55048),
            .in3(N__55024),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n691 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17748 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_18_6  (
            .in0(_gnd_net_),
            .in1(N__55021),
            .in2(N__55009),
            .in3(N__54847),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n742 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17749 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_LUT4_0_LC_21_18_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_LUT4_0_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_LUT4_0_LC_21_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_LUT4_0_LC_21_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54844),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i5_LC_21_19_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i5_LC_21_19_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i5_LC_21_19_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i5_LC_21_19_3  (
            .in0(N__56478),
            .in1(N__56363),
            .in2(_gnd_net_),
            .in3(N__62697),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62109),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i1_LC_21_19_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i1_LC_21_19_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i1_LC_21_19_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i1_LC_21_19_4  (
            .in0(N__56361),
            .in1(N__56476),
            .in2(_gnd_net_),
            .in3(N__60151),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62109),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i3_LC_21_19_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i3_LC_21_19_5 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i3_LC_21_19_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i3_LC_21_19_5  (
            .in0(N__56477),
            .in1(N__56362),
            .in2(_gnd_net_),
            .in3(N__60097),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62109),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i22_LC_21_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i22_LC_21_20_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i22_LC_21_20_0 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i22_LC_21_20_0  (
            .in0(N__56330),
            .in1(_gnd_net_),
            .in2(N__56479),
            .in3(N__57419),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62114),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i0_LC_21_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i0_LC_21_20_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i0_LC_21_20_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i0_LC_21_20_1  (
            .in0(N__60127),
            .in1(N__56329),
            .in2(_gnd_net_),
            .in3(N__56443),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62114),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i28_LC_21_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i28_LC_21_20_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i28_LC_21_20_2 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i28_LC_21_20_2  (
            .in0(N__56448),
            .in1(_gnd_net_),
            .in2(N__56360),
            .in3(N__57938),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62114),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i25_LC_21_20_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i25_LC_21_20_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i25_LC_21_20_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_i25_LC_21_20_3  (
            .in0(N__58109),
            .in1(N__56447),
            .in2(_gnd_net_),
            .in3(N__56331),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.currentControlITerm_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62114),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_280_LC_21_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_280_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_280_LC_21_20_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_280_LC_21_20_4  (
            .in0(N__57635),
            .in1(N__57787),
            .in2(N__57718),
            .in3(N__60163),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_281_LC_21_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_281_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_281_LC_21_20_5 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_281_LC_21_20_5  (
            .in0(N__57420),
            .in1(N__57491),
            .in2(N__56233),
            .in3(N__57551),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20654_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_282_LC_21_20_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_282_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_282_LC_21_20_6 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_282_LC_21_20_6  (
            .in0(N__58169),
            .in1(N__58110),
            .in2(N__56230),
            .in3(N__58238),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20640_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i14382_4_lut_LC_21_20_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i14382_4_lut_LC_21_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i14382_4_lut_LC_21_20_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i14382_4_lut_LC_21_20_7  (
            .in0(N__58040),
            .in1(N__57939),
            .in2(N__56611),
            .in3(N__57986),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_563_2_lut_LC_21_21_0  (
            .in0(_gnd_net_),
            .in1(N__64632),
            .in2(N__64844),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n57 ),
            .ltout(),
            .carryin(bfn_21_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18174 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_21_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_3_lut_LC_21_21_1  (
            .in0(N__56778),
            .in1(N__56602),
            .in2(N__64489),
            .in3(N__56596),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_4 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18174 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18175 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_21_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_4_lut_LC_21_21_2  (
            .in0(N__56782),
            .in1(N__64101),
            .in2(N__56593),
            .in3(N__56575),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_5 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18175 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18176 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_21_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_5_lut_LC_21_21_3  (
            .in0(N__56779),
            .in1(N__56572),
            .in2(N__63936),
            .in3(N__56560),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_6 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18176 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18177 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_21_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_21_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_6_lut_LC_21_21_4  (
            .in0(N__56783),
            .in1(N__56557),
            .in2(N__63609),
            .in3(N__56545),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_7 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18177 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18178 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_21_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_21_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_7_lut_LC_21_21_5  (
            .in0(N__56780),
            .in1(N__56542),
            .in2(N__63399),
            .in3(N__56530),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_8 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18178 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18179 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_21_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_21_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_8_lut_LC_21_21_6  (
            .in0(N__56784),
            .in1(N__56527),
            .in2(N__63065),
            .in3(N__56512),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_9 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18179 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18180 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_21_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_21_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_9_lut_LC_21_21_7  (
            .in0(N__56781),
            .in1(N__56509),
            .in2(N__66875),
            .in3(N__56497),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_10 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18180 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18181 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_10_lut_LC_21_22_0  (
            .in0(N__56801),
            .in1(N__56884),
            .in2(N__66521),
            .in3(N__56872),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_11 ),
            .ltout(),
            .carryin(bfn_21_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18182 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_22_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_11_lut_LC_21_22_1  (
            .in0(N__56804),
            .in1(N__56869),
            .in2(N__66261),
            .in3(N__56857),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_12 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18182 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18183 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_22_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_12_lut_LC_21_22_2  (
            .in0(N__56802),
            .in1(N__56854),
            .in2(N__66012),
            .in3(N__56842),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18183 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18184 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_22_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_13_lut_LC_21_22_3  (
            .in0(N__56805),
            .in1(N__56839),
            .in2(N__65791),
            .in3(N__56827),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_14 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18184 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18185 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_22_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_14_lut_LC_21_22_4  (
            .in0(N__56803),
            .in1(N__56707),
            .in2(N__65570),
            .in3(N__56695),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Switch_out1_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18185 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18186 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_15_lut_LC_21_22_5  (
            .in0(_gnd_net_),
            .in1(N__65342),
            .in2(N__56692),
            .in3(N__56662),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n691 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18186 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18187 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_562_16_lut_LC_21_22_6  (
            .in0(_gnd_net_),
            .in1(N__56659),
            .in2(N__65178),
            .in3(N__56632),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n742 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18187 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_LUT4_0_LC_21_22_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_LUT4_0_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_LUT4_0_LC_21_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_LUT4_0_LC_21_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56629),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n743_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_2_lut_LC_21_23_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_2_lut_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_2_lut_LC_21_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_2_lut_LC_21_23_0  (
            .in0(_gnd_net_),
            .in1(N__57082),
            .in2(N__57073),
            .in3(_gnd_net_),
            .lcout(Add_add_temp_4_adj_2416),
            .ltout(),
            .carryin(bfn_21_23_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_3_lut_LC_21_23_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_3_lut_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_3_lut_LC_21_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_3_lut_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(N__57061),
            .in2(N__57052),
            .in3(N__57040),
            .lcout(Add_add_temp_5_adj_2415),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15913 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_4_lut_LC_21_23_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_4_lut_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_4_lut_LC_21_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_4_lut_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(N__57037),
            .in2(N__57028),
            .in3(N__57013),
            .lcout(Add_add_temp_6_adj_2414),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15914 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15915 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_5_lut_LC_21_23_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_5_lut_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_5_lut_LC_21_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_5_lut_LC_21_23_3  (
            .in0(_gnd_net_),
            .in1(N__57010),
            .in2(N__57001),
            .in3(N__56989),
            .lcout(Add_add_temp_7_adj_2413),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15915 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15916 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_6_lut_LC_21_23_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_6_lut_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_6_lut_LC_21_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_6_lut_LC_21_23_4  (
            .in0(_gnd_net_),
            .in1(N__56986),
            .in2(N__56980),
            .in3(N__56968),
            .lcout(Add_add_temp_8_adj_2412),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15916 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15917 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_7_lut_LC_21_23_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_7_lut_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_7_lut_LC_21_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_7_lut_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(N__56965),
            .in2(N__56956),
            .in3(N__56944),
            .lcout(Add_add_temp_9_adj_2411),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15917 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15918 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_8_lut_LC_21_23_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_8_lut_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_8_lut_LC_21_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_8_lut_LC_21_23_6  (
            .in0(_gnd_net_),
            .in1(N__56941),
            .in2(N__56932),
            .in3(N__56920),
            .lcout(Add_add_temp_10_adj_2410),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15918 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15919 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_9_lut_LC_21_23_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_9_lut_LC_21_23_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_9_lut_LC_21_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_9_lut_LC_21_23_7  (
            .in0(_gnd_net_),
            .in1(N__56917),
            .in2(N__56896),
            .in3(N__56887),
            .lcout(Add_add_temp_11_adj_2409),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15919 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15920 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_10_lut_LC_21_24_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_10_lut_LC_21_24_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_10_lut_LC_21_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_10_lut_LC_21_24_0  (
            .in0(_gnd_net_),
            .in1(N__57385),
            .in2(N__57367),
            .in3(N__57352),
            .lcout(Add_add_temp_12_adj_2408),
            .ltout(),
            .carryin(bfn_21_24_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15921 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_11_lut_LC_21_24_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_11_lut_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_11_lut_LC_21_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_11_lut_LC_21_24_1  (
            .in0(_gnd_net_),
            .in1(N__57349),
            .in2(N__57340),
            .in3(N__57316),
            .lcout(Add_add_temp_13_adj_2407),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15921 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15922 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_12_lut_LC_21_24_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_12_lut_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_12_lut_LC_21_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_12_lut_LC_21_24_2  (
            .in0(_gnd_net_),
            .in1(N__57313),
            .in2(N__57304),
            .in3(N__57280),
            .lcout(Add_add_temp_14_adj_2406),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15922 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15923 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_13_lut_LC_21_24_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_13_lut_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_13_lut_LC_21_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_13_lut_LC_21_24_3  (
            .in0(_gnd_net_),
            .in1(N__57277),
            .in2(N__57253),
            .in3(N__57238),
            .lcout(Add_add_temp_15_adj_2405),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15923 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15924 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_14_lut_LC_21_24_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_14_lut_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_14_lut_LC_21_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_14_lut_LC_21_24_4  (
            .in0(_gnd_net_),
            .in1(N__57235),
            .in2(N__57223),
            .in3(N__57202),
            .lcout(Add_add_temp_16_adj_2404),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15924 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15925 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_15_lut_LC_21_24_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_15_lut_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_15_lut_LC_21_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_15_lut_LC_21_24_5  (
            .in0(_gnd_net_),
            .in1(N__57199),
            .in2(N__57178),
            .in3(N__57163),
            .lcout(Add_add_temp_17_adj_2403),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15925 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15926 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_16_lut_LC_21_24_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_16_lut_LC_21_24_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_16_lut_LC_21_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_16_lut_LC_21_24_6  (
            .in0(_gnd_net_),
            .in1(N__57160),
            .in2(N__57136),
            .in3(N__57121),
            .lcout(Add_add_temp_18_adj_2402),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15926 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15927 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_17_lut_LC_21_24_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_17_lut_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_17_lut_LC_21_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_17_lut_LC_21_24_7  (
            .in0(_gnd_net_),
            .in1(N__57118),
            .in2(N__57097),
            .in3(N__57862),
            .lcout(Add_add_temp_19_adj_2401),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15927 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15928 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_18_lut_LC_21_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_18_lut_LC_21_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_18_lut_LC_21_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_18_lut_LC_21_25_0  (
            .in0(_gnd_net_),
            .in1(N__57859),
            .in2(N__57841),
            .in3(N__57823),
            .lcout(Add_add_temp_20_adj_2400),
            .ltout(),
            .carryin(bfn_21_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_19_lut_LC_21_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_19_lut_LC_21_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_19_lut_LC_21_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_19_lut_LC_21_25_1  (
            .in0(_gnd_net_),
            .in1(N__57820),
            .in2(N__57802),
            .in3(N__57754),
            .lcout(Add_add_temp_21_adj_2399),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15929 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_20_lut_LC_21_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_20_lut_LC_21_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_20_lut_LC_21_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_20_lut_LC_21_25_2  (
            .in0(_gnd_net_),
            .in1(N__57751),
            .in2(N__57733),
            .in3(N__57688),
            .lcout(Add_add_temp_22_adj_2398),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15930 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_21_lut_LC_21_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_21_lut_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_21_lut_LC_21_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_21_lut_LC_21_25_3  (
            .in0(_gnd_net_),
            .in1(N__57685),
            .in2(N__57658),
            .in3(N__57604),
            .lcout(Add_add_temp_23_adj_2397),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15931 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_22_lut_LC_21_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_22_lut_LC_21_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_22_lut_LC_21_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_22_lut_LC_21_25_4  (
            .in0(_gnd_net_),
            .in1(N__57601),
            .in2(N__57577),
            .in3(N__57532),
            .lcout(Add_add_temp_24_adj_2396),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15932 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_23_lut_LC_21_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_23_lut_LC_21_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_23_lut_LC_21_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_23_lut_LC_21_25_5  (
            .in0(_gnd_net_),
            .in1(N__57529),
            .in2(N__57508),
            .in3(N__57466),
            .lcout(Add_add_temp_25_adj_2395),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15933 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15934 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_24_lut_LC_21_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_24_lut_LC_21_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_24_lut_LC_21_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_24_lut_LC_21_25_6  (
            .in0(_gnd_net_),
            .in1(N__57456),
            .in2(N__57439),
            .in3(N__57388),
            .lcout(Add_add_temp_26_adj_2394),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15934 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_25_lut_LC_21_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_25_lut_LC_21_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_25_lut_LC_21_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_25_lut_LC_21_25_7  (
            .in0(_gnd_net_),
            .in1(N__58279),
            .in2(N__58255),
            .in3(N__58216),
            .lcout(Add_add_temp_27_adj_2393),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15935 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_26_lut_LC_21_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_26_lut_LC_21_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_26_lut_LC_21_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_26_lut_LC_21_26_0  (
            .in0(_gnd_net_),
            .in1(N__58212),
            .in2(N__58186),
            .in3(N__58150),
            .lcout(Add_add_temp_28_adj_2392),
            .ltout(),
            .carryin(bfn_21_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_27_lut_LC_21_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_27_lut_LC_21_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_27_lut_LC_21_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_27_lut_LC_21_26_1  (
            .in0(_gnd_net_),
            .in1(N__58140),
            .in2(N__58126),
            .in3(N__58084),
            .lcout(Add_add_temp_29_adj_2391),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15937 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_28_lut_LC_21_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_28_lut_LC_21_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_28_lut_LC_21_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_28_lut_LC_21_26_2  (
            .in0(_gnd_net_),
            .in1(N__58081),
            .in2(N__58057),
            .in3(N__58018),
            .lcout(Add_add_temp_30_adj_2390),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15938 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_29_lut_LC_21_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_29_lut_LC_21_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_29_lut_LC_21_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_29_lut_LC_21_26_3  (
            .in0(_gnd_net_),
            .in1(N__58015),
            .in2(N__58403),
            .in3(N__57967),
            .lcout(Add_add_temp_31_adj_2389),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15939 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_30_lut_LC_21_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_30_lut_LC_21_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_30_lut_LC_21_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_30_lut_LC_21_26_4  (
            .in0(_gnd_net_),
            .in1(N__58395),
            .in2(N__57963),
            .in3(N__57916),
            .lcout(Add_add_temp_32_adj_2388),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15940 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15941 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_31_lut_LC_21_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_31_lut_LC_21_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_31_lut_LC_21_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_31_lut_LC_21_26_5  (
            .in0(_gnd_net_),
            .in1(N__57913),
            .in2(N__58404),
            .in3(N__57865),
            .lcout(Add_add_temp_33_adj_2387),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15941 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_32_lut_LC_21_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_32_lut_LC_21_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_32_lut_LC_21_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_32_lut_LC_21_26_6  (
            .in0(_gnd_net_),
            .in1(N__58399),
            .in2(N__58519),
            .in3(N__58459),
            .lcout(Add_add_temp_34_adj_2386),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15942 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_33_lut_LC_21_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_33_lut_LC_21_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_33_lut_LC_21_26_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.add_560_33_lut_LC_21_26_7  (
            .in0(N__58456),
            .in1(_gnd_net_),
            .in2(N__58405),
            .in3(N__58372),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.Saturate_out1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_21_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_21_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_21_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_571_2_lut_LC_21_28_0  (
            .in0(_gnd_net_),
            .in1(N__64899),
            .in2(N__64749),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n81 ),
            .ltout(),
            .carryin(bfn_21_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18294 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_21_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_21_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_21_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_3_lut_LC_21_28_1  (
            .in0(_gnd_net_),
            .in1(N__58339),
            .in2(N__64497),
            .in3(N__58333),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n127 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18294 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18295 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_21_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_21_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_21_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_4_lut_LC_21_28_2  (
            .in0(_gnd_net_),
            .in1(N__58330),
            .in2(N__64236),
            .in3(N__58324),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n176 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18295 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18296 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_21_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_21_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_21_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_5_lut_LC_21_28_3  (
            .in0(_gnd_net_),
            .in1(N__58321),
            .in2(N__63981),
            .in3(N__58315),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n225 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18296 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18297 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_21_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_21_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_21_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_6_lut_LC_21_28_4  (
            .in0(_gnd_net_),
            .in1(N__63630),
            .in2(N__58312),
            .in3(N__58303),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n274 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18297 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18298 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_21_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_21_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_21_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_7_lut_LC_21_28_5  (
            .in0(_gnd_net_),
            .in1(N__58300),
            .in2(N__63401),
            .in3(N__58294),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n323 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18298 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18299 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_21_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_21_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_21_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_8_lut_LC_21_28_6  (
            .in0(_gnd_net_),
            .in1(N__63094),
            .in2(N__58291),
            .in3(N__58282),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n372_adj_596 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18299 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18300 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_21_28_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_21_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_21_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_9_lut_LC_21_28_7  (
            .in0(_gnd_net_),
            .in1(N__66884),
            .in2(N__58615),
            .in3(N__58606),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n421_adj_595 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18300 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18301 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_21_29_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_21_29_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_21_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_10_lut_LC_21_29_0  (
            .in0(_gnd_net_),
            .in1(N__66638),
            .in2(N__58603),
            .in3(N__58594),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n470_adj_594 ),
            .ltout(),
            .carryin(bfn_21_29_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18302 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_21_29_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_21_29_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_21_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_11_lut_LC_21_29_1  (
            .in0(_gnd_net_),
            .in1(N__58591),
            .in2(N__66347),
            .in3(N__58585),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n519_adj_593 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18302 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18303 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_21_29_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_21_29_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_21_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_12_lut_LC_21_29_2  (
            .in0(_gnd_net_),
            .in1(N__58582),
            .in2(N__66094),
            .in3(N__58576),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n568_adj_592 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18303 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18304 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_21_29_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_21_29_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_21_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_13_lut_LC_21_29_3  (
            .in0(_gnd_net_),
            .in1(N__58573),
            .in2(N__65832),
            .in3(N__58567),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n617_adj_591 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18304 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18305 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_21_29_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_21_29_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_21_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_14_lut_LC_21_29_4  (
            .in0(_gnd_net_),
            .in1(N__58564),
            .in2(N__65602),
            .in3(N__58558),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n666 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18305 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18306 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_21_29_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_21_29_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_21_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_15_lut_LC_21_29_5  (
            .in0(_gnd_net_),
            .in1(N__65387),
            .in2(N__58555),
            .in3(N__58546),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n715 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18306 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18307 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_21_29_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_21_29_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_21_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_16_lut_LC_21_29_6  (
            .in0(_gnd_net_),
            .in1(N__65203),
            .in2(N__58543),
            .in3(N__58522),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n774_adj_589 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18307 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_LUT4_0_LC_21_29_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_LUT4_0_LC_21_29_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_LUT4_0_LC_21_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_LUT4_0_LC_21_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58936),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n775_adj_590_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_22_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_22_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_2_lut_LC_22_11_0  (
            .in0(_gnd_net_),
            .in1(N__58865),
            .in2(N__60951),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n54 ),
            .ltout(),
            .carryin(bfn_22_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17536 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_22_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_22_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_3_lut_LC_22_11_1  (
            .in0(_gnd_net_),
            .in1(N__60914),
            .in2(N__58687),
            .in3(N__58678),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n103 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17536 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17537 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_22_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_22_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_4_lut_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(N__58675),
            .in2(N__60952),
            .in3(N__58669),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n152 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17537 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17538 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_22_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_22_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_5_lut_LC_22_11_3  (
            .in0(_gnd_net_),
            .in1(N__60918),
            .in2(N__58666),
            .in3(N__58657),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n201 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17538 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17539 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_22_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_22_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_6_lut_LC_22_11_4  (
            .in0(_gnd_net_),
            .in1(N__58654),
            .in2(N__60953),
            .in3(N__58648),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n250 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17539 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17540 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_22_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_22_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_7_lut_LC_22_11_5  (
            .in0(_gnd_net_),
            .in1(N__60922),
            .in2(N__58645),
            .in3(N__58636),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n299 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17540 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17541 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_22_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_22_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_8_lut_LC_22_11_6  (
            .in0(_gnd_net_),
            .in1(N__58633),
            .in2(N__60954),
            .in3(N__58627),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n348 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17541 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17542 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_22_11_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_22_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_9_lut_LC_22_11_7  (
            .in0(_gnd_net_),
            .in1(N__60926),
            .in2(N__58624),
            .in3(N__59065),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n397 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17542 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17543 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_22_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_22_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_10_lut_LC_22_12_0  (
            .in0(_gnd_net_),
            .in1(N__59062),
            .in2(N__60955),
            .in3(N__59056),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n446 ),
            .ltout(),
            .carryin(bfn_22_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17544 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_22_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_22_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_11_lut_LC_22_12_1  (
            .in0(_gnd_net_),
            .in1(N__60930),
            .in2(N__59053),
            .in3(N__59044),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n495 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17544 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17545 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_22_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_22_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_12_lut_LC_22_12_2  (
            .in0(_gnd_net_),
            .in1(N__59041),
            .in2(N__60956),
            .in3(N__59035),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n544 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17545 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17546 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_22_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_22_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_13_lut_LC_22_12_3  (
            .in0(_gnd_net_),
            .in1(N__60934),
            .in2(N__59032),
            .in3(N__59023),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n593 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17546 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17547 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_22_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_22_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_14_lut_LC_22_12_4  (
            .in0(_gnd_net_),
            .in1(N__59020),
            .in2(N__60957),
            .in3(N__59014),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n642 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17547 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17548 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_22_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_22_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_15_lut_LC_22_12_5  (
            .in0(_gnd_net_),
            .in1(N__60938),
            .in2(N__59011),
            .in3(N__59002),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n691_adj_440 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17548 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_22_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_22_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_562_16_lut_LC_22_12_6  (
            .in0(_gnd_net_),
            .in1(N__58999),
            .in2(N__58993),
            .in3(N__58954),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n742_adj_411 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17549 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_LUT4_0_LC_22_12_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_LUT4_0_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_LUT4_0_LC_22_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_LUT4_0_LC_22_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58951),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n743_adj_410_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_117_LC_22_13_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_117_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_117_LC_22_13_0 .LUT_INIT=16'b1111010010101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_117_LC_22_13_0  (
            .in0(N__69156),
            .in1(N__61378),
            .in2(N__61475),
            .in3(N__69108),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_LC_22_13_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_LC_22_13_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_LC_22_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__59107),
            .in3(N__61156),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13171_2_lut_3_lut_LC_22_13_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13171_2_lut_3_lut_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13171_2_lut_3_lut_LC_22_13_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13171_2_lut_3_lut_LC_22_13_2  (
            .in0(N__61450),
            .in1(N__61381),
            .in2(_gnd_net_),
            .in3(N__68800),
            .lcout(\foc.dVoltage_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13164_2_lut_3_lut_LC_22_13_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13164_2_lut_3_lut_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13164_2_lut_3_lut_LC_22_13_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13164_2_lut_3_lut_LC_22_13_3  (
            .in0(N__61379),
            .in1(N__61449),
            .in2(_gnd_net_),
            .in3(N__68188),
            .lcout(),
            .ltout(\foc.dVoltage_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i15_2_lut_LC_22_13_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i15_2_lut_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i15_2_lut_LC_22_13_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.equal_13243_i15_2_lut_LC_22_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__59098),
            .in3(N__68187),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_120_LC_22_13_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_120_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_120_LC_22_13_5 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_120_LC_22_13_5  (
            .in0(N__68799),
            .in1(N__59095),
            .in2(N__59089),
            .in3(N__59086),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12820_4_lut_LC_22_13_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12820_4_lut_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12820_4_lut_LC_22_13_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12820_4_lut_LC_22_13_6  (
            .in0(N__69157),
            .in1(N__69109),
            .in2(N__69010),
            .in3(N__61162),
            .lcout(\foc.Out_31__N_332_adj_2312 ),
            .ltout(\foc.Out_31__N_332_adj_2312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13167_2_lut_3_lut_LC_22_13_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13167_2_lut_3_lut_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13167_2_lut_3_lut_LC_22_13_7 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13167_2_lut_3_lut_LC_22_13_7  (
            .in0(N__61380),
            .in1(_gnd_net_),
            .in2(N__59074),
            .in3(N__67977),
            .lcout(\foc.dVoltage_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1212_rep_6_4_lut_LC_22_14_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1212_rep_6_4_lut_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1212_rep_6_4_lut_LC_22_14_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1212_rep_6_4_lut_LC_22_14_0  (
            .in0(N__61294),
            .in1(N__61312),
            .in2(N__69006),
            .in3(N__69107),
            .lcout(\foc.Out_31__N_333_adj_2310 ),
            .ltout(\foc.Out_31__N_333_adj_2310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13173_2_lut_3_lut_LC_22_14_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13173_2_lut_3_lut_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13173_2_lut_3_lut_LC_22_14_1 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13173_2_lut_3_lut_LC_22_14_1  (
            .in0(_gnd_net_),
            .in1(N__68659),
            .in2(N__59230),
            .in3(N__61459),
            .lcout(\foc.dVoltage_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13162_2_lut_3_lut_LC_22_14_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13162_2_lut_3_lut_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13162_2_lut_3_lut_LC_22_14_2 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13162_2_lut_3_lut_LC_22_14_2  (
            .in0(N__67555),
            .in1(N__61477),
            .in2(_gnd_net_),
            .in3(N__61371),
            .lcout(),
            .ltout(\foc.dVoltage_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_126_LC_22_14_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_126_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_126_LC_22_14_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_126_LC_22_14_3  (
            .in0(N__59227),
            .in1(N__68658),
            .in2(N__59221),
            .in3(N__67554),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13170_2_lut_3_lut_LC_22_14_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13170_2_lut_3_lut_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13170_2_lut_3_lut_LC_22_14_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13170_2_lut_3_lut_LC_22_14_4  (
            .in0(N__61458),
            .in1(N__68872),
            .in2(_gnd_net_),
            .in3(N__61372),
            .lcout(),
            .ltout(\foc.dVoltage_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_123_LC_22_14_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_123_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_123_LC_22_14_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_123_LC_22_14_5  (
            .in0(N__68871),
            .in1(N__67898),
            .in2(N__59212),
            .in3(N__59209),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13204_2_lut_3_lut_LC_22_14_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13204_2_lut_3_lut_LC_22_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13204_2_lut_3_lut_LC_22_14_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13204_2_lut_3_lut_LC_22_14_6  (
            .in0(N__59197),
            .in1(N__59325),
            .in2(_gnd_net_),
            .in3(N__59443),
            .lcout(),
            .ltout(\foc.qVoltage_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_263_LC_22_14_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_263_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_263_LC_22_14_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_263_LC_22_14_7  (
            .in0(N__59359),
            .in1(N__59196),
            .in2(N__59164),
            .in3(N__59239),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.equal_13244_i21_2_lut_3_lut_LC_22_15_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.equal_13244_i21_2_lut_3_lut_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.equal_13244_i21_2_lut_3_lut_LC_22_15_3 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.equal_13244_i21_2_lut_3_lut_LC_22_15_3  (
            .in0(N__59429),
            .in1(N__59155),
            .in2(_gnd_net_),
            .in3(N__59306),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_268_LC_22_15_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_268_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_268_LC_22_15_4 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_268_LC_22_15_4  (
            .in0(N__59449),
            .in1(N__59481),
            .in2(N__59131),
            .in3(N__59128),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13208_2_lut_3_lut_LC_22_15_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13208_2_lut_3_lut_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13208_2_lut_3_lut_LC_22_15_5 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13208_2_lut_3_lut_LC_22_15_5  (
            .in0(N__59482),
            .in1(_gnd_net_),
            .in2(N__59441),
            .in3(N__59307),
            .lcout(\foc.qVoltage_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13214_2_lut_3_lut_LC_22_15_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13214_2_lut_3_lut_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13214_2_lut_3_lut_LC_22_15_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.u_Saturate_Output.i13214_2_lut_3_lut_LC_22_15_7  (
            .in0(N__59433),
            .in1(N__59358),
            .in2(_gnd_net_),
            .in3(N__59308),
            .lcout(\foc.qVoltage_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i30_LC_22_16_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i30_LC_22_16_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i30_LC_22_16_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i30_LC_22_16_1  (
            .in0(N__61974),
            .in1(N__61629),
            .in2(_gnd_net_),
            .in3(N__61910),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62110),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i0_LC_22_16_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i0_LC_22_16_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i0_LC_22_16_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i0_LC_22_16_2  (
            .in0(N__61907),
            .in1(N__61971),
            .in2(_gnd_net_),
            .in3(N__62551),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62110),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i27_LC_22_16_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i27_LC_22_16_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i27_LC_22_16_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i27_LC_22_16_3  (
            .in0(N__61972),
            .in1(N__61908),
            .in2(_gnd_net_),
            .in3(N__61712),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62110),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i29_LC_22_16_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i29_LC_22_16_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i29_LC_22_16_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i29_LC_22_16_7  (
            .in0(N__61973),
            .in1(N__61909),
            .in2(_gnd_net_),
            .in3(N__61597),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62110),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i6_LC_22_17_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i6_LC_22_17_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i6_LC_22_17_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i6_LC_22_17_0  (
            .in0(N__61906),
            .in1(N__61970),
            .in2(_gnd_net_),
            .in3(N__62416),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13327_4_lut_LC_22_17_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13327_4_lut_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13327_4_lut_LC_22_17_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i13327_4_lut_LC_22_17_1  (
            .in0(N__59614),
            .in1(N__61685),
            .in2(N__61716),
            .in3(N__61655),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_139_LC_22_17_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_139_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_139_LC_22_17_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_139_LC_22_17_2  (
            .in0(N__61592),
            .in1(N__62142),
            .in2(N__59233),
            .in3(N__61622),
            .lcout(Saturate_out1_31__N_267),
            .ltout(Saturate_out1_31__N_267_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i18_LC_22_17_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i18_LC_22_17_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i18_LC_22_17_3 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i18_LC_22_17_3  (
            .in0(N__62175),
            .in1(_gnd_net_),
            .in2(N__59491),
            .in3(N__61901),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i1_LC_22_17_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i1_LC_22_17_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i1_LC_22_17_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i1_LC_22_17_4  (
            .in0(N__61902),
            .in1(N__62569),
            .in2(_gnd_net_),
            .in3(N__61966),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i3_LC_22_17_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i3_LC_22_17_5 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i3_LC_22_17_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i3_LC_22_17_5  (
            .in0(N__61969),
            .in1(N__61905),
            .in2(_gnd_net_),
            .in3(N__62518),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i2_LC_22_17_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i2_LC_22_17_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i2_LC_22_17_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i2_LC_22_17_6  (
            .in0(N__61904),
            .in1(N__61968),
            .in2(_gnd_net_),
            .in3(N__62490),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i20_LC_22_17_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i20_LC_22_17_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i20_LC_22_17_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i20_LC_22_17_7  (
            .in0(N__61967),
            .in1(N__61903),
            .in2(_gnd_net_),
            .in3(N__59791),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62104),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i24_LC_22_18_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i24_LC_22_18_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i24_LC_22_18_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i24_LC_22_18_0  (
            .in0(N__61911),
            .in1(N__61985),
            .in2(_gnd_net_),
            .in3(N__60005),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62111),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i25_LC_22_18_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i25_LC_22_18_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i25_LC_22_18_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i25_LC_22_18_1  (
            .in0(N__61986),
            .in1(N__61912),
            .in2(_gnd_net_),
            .in3(N__59972),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62111),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_143_LC_22_18_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_143_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_143_LC_22_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_143_LC_22_18_2  (
            .in0(N__62307),
            .in1(N__62250),
            .in2(N__62284),
            .in3(N__61789),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19842_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_144_LC_22_18_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_144_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_144_LC_22_18_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_144_LC_22_18_3  (
            .in0(N__62226),
            .in1(N__62202),
            .in2(N__59488),
            .in3(N__62176),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20666_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_145_LC_22_18_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_145_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_145_LC_22_18_4 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_145_LC_22_18_4  (
            .in0(N__61551),
            .in1(N__62060),
            .in2(N__59485),
            .in3(N__59787),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_146_LC_22_18_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_146_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_146_LC_22_18_5 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_146_LC_22_18_5  (
            .in0(N__60007),
            .in1(N__59974),
            .in2(N__59620),
            .in3(N__61530),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_137_LC_22_18_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_137_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_137_LC_22_18_6 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_137_LC_22_18_6  (
            .in0(N__61550),
            .in1(N__62152),
            .in2(N__62064),
            .in3(N__59786),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20648_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_138_LC_22_18_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_138_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_138_LC_22_18_7 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_138_LC_22_18_7  (
            .in0(N__60006),
            .in1(N__59973),
            .in2(N__59617),
            .in3(N__61529),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_2_lut_LC_22_19_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_2_lut_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_2_lut_LC_22_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_2_lut_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(N__59608),
            .in2(N__59599),
            .in3(_gnd_net_),
            .lcout(Add_add_temp_4),
            .ltout(),
            .carryin(bfn_22_19_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_3_lut_LC_22_19_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_3_lut_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_3_lut_LC_22_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_3_lut_LC_22_19_1  (
            .in0(_gnd_net_),
            .in1(N__59587),
            .in2(N__59578),
            .in3(N__59563),
            .lcout(Add_add_temp_5),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15973 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_4_lut_LC_22_19_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_4_lut_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_4_lut_LC_22_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_4_lut_LC_22_19_2  (
            .in0(_gnd_net_),
            .in1(N__59560),
            .in2(N__59551),
            .in3(N__59539),
            .lcout(Add_add_temp_6),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15974 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_5_lut_LC_22_19_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_5_lut_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_5_lut_LC_22_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_5_lut_LC_22_19_3  (
            .in0(_gnd_net_),
            .in1(N__59536),
            .in2(N__59527),
            .in3(N__59512),
            .lcout(Add_add_temp_7),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15975 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_6_lut_LC_22_19_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_6_lut_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_6_lut_LC_22_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_6_lut_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__61561),
            .in2(N__59509),
            .in3(N__59494),
            .lcout(Add_add_temp_8),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15976 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15977 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_7_lut_LC_22_19_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_7_lut_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_7_lut_LC_22_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_7_lut_LC_22_19_5  (
            .in0(_gnd_net_),
            .in1(N__62035),
            .in2(N__59749),
            .in3(N__59737),
            .lcout(Add_add_temp_9),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15977 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_8_lut_LC_22_19_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_8_lut_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_8_lut_LC_22_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_8_lut_LC_22_19_6  (
            .in0(_gnd_net_),
            .in1(N__59734),
            .in2(N__59725),
            .in3(N__59710),
            .lcout(Add_add_temp_10),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15978 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15979 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_9_lut_LC_22_19_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_9_lut_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_9_lut_LC_22_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_9_lut_LC_22_19_7  (
            .in0(_gnd_net_),
            .in1(N__59707),
            .in2(N__67510),
            .in3(N__59701),
            .lcout(Add_add_temp_11),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15979 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15980 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_10_lut_LC_22_20_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_10_lut_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_10_lut_LC_22_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_10_lut_LC_22_20_0  (
            .in0(_gnd_net_),
            .in1(N__67492),
            .in2(N__59698),
            .in3(N__59686),
            .lcout(Add_add_temp_12),
            .ltout(),
            .carryin(bfn_22_20_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15981 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_11_lut_LC_22_20_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_11_lut_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_11_lut_LC_22_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_11_lut_LC_22_20_1  (
            .in0(_gnd_net_),
            .in1(N__67210),
            .in2(N__59683),
            .in3(N__59671),
            .lcout(Add_add_temp_13),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15981 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15982 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_12_lut_LC_22_20_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_12_lut_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_12_lut_LC_22_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_12_lut_LC_22_20_2  (
            .in0(_gnd_net_),
            .in1(N__67168),
            .in2(N__59668),
            .in3(N__59656),
            .lcout(Add_add_temp_14),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15982 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15983 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_13_lut_LC_22_20_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_13_lut_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_13_lut_LC_22_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_13_lut_LC_22_20_3  (
            .in0(_gnd_net_),
            .in1(N__59653),
            .in2(N__67126),
            .in3(N__59644),
            .lcout(Add_add_temp_15),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15983 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15984 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_14_lut_LC_22_20_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_14_lut_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_14_lut_LC_22_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_14_lut_LC_22_20_4  (
            .in0(_gnd_net_),
            .in1(N__67081),
            .in2(N__59641),
            .in3(N__59623),
            .lcout(Add_add_temp_16),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15984 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15985 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_15_lut_LC_22_20_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_15_lut_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_15_lut_LC_22_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_15_lut_LC_22_20_5  (
            .in0(_gnd_net_),
            .in1(N__67042),
            .in2(N__59923),
            .in3(N__59908),
            .lcout(Add_add_temp_17),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15985 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15986 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_16_lut_LC_22_20_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_16_lut_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_16_lut_LC_22_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_16_lut_LC_22_20_6  (
            .in0(_gnd_net_),
            .in1(N__67843),
            .in2(N__59905),
            .in3(N__59890),
            .lcout(Add_add_temp_18),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15986 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15987 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_17_lut_LC_22_20_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_17_lut_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_17_lut_LC_22_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_17_lut_LC_22_20_7  (
            .in0(_gnd_net_),
            .in1(N__59887),
            .in2(N__67816),
            .in3(N__59875),
            .lcout(Add_add_temp_19),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15987 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15988 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_18_lut_LC_22_21_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_18_lut_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_18_lut_LC_22_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_18_lut_LC_22_21_0  (
            .in0(_gnd_net_),
            .in1(N__67765),
            .in2(N__59872),
            .in3(N__59857),
            .lcout(Add_add_temp_20),
            .ltout(),
            .carryin(bfn_22_21_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15989 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_19_lut_LC_22_21_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_19_lut_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_19_lut_LC_22_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_19_lut_LC_22_21_1  (
            .in0(_gnd_net_),
            .in1(N__67702),
            .in2(N__59854),
            .in3(N__59839),
            .lcout(Add_add_temp_21),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15989 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15990 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_20_lut_LC_22_21_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_20_lut_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_20_lut_LC_22_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_20_lut_LC_22_21_2  (
            .in0(_gnd_net_),
            .in1(N__67651),
            .in2(N__59836),
            .in3(N__59821),
            .lcout(Add_add_temp_22),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15990 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15991 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_21_lut_LC_22_21_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_21_lut_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_21_lut_LC_22_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_21_lut_LC_22_21_3  (
            .in0(_gnd_net_),
            .in1(N__59818),
            .in2(N__67588),
            .in3(N__59806),
            .lcout(Add_add_temp_23),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15991 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15992 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_22_lut_LC_22_21_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_22_lut_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_22_lut_LC_22_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_22_lut_LC_22_21_4  (
            .in0(_gnd_net_),
            .in1(N__59803),
            .in2(N__68500),
            .in3(N__59770),
            .lcout(Add_add_temp_24),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15992 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15993 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_23_lut_LC_22_21_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_23_lut_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_23_lut_LC_22_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_23_lut_LC_22_21_5  (
            .in0(_gnd_net_),
            .in1(N__68218),
            .in2(N__59767),
            .in3(N__59752),
            .lcout(Add_add_temp_25),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15993 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15994 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_24_lut_LC_22_21_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_24_lut_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_24_lut_LC_22_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_24_lut_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__60055),
            .in2(N__68143),
            .in3(N__60043),
            .lcout(Add_add_temp_26),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15994 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15995 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_25_lut_LC_22_21_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_25_lut_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_25_lut_LC_22_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_25_lut_LC_22_21_7  (
            .in0(_gnd_net_),
            .in1(N__68080),
            .in2(N__60040),
            .in3(N__60025),
            .lcout(Add_add_temp_27),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15995 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15996 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_26_lut_LC_22_22_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_26_lut_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_26_lut_LC_22_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_26_lut_LC_22_22_0  (
            .in0(_gnd_net_),
            .in1(N__68017),
            .in2(N__60022),
            .in3(N__59992),
            .lcout(Add_add_temp_28),
            .ltout(),
            .carryin(bfn_22_22_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15997 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_27_lut_LC_22_22_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_27_lut_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_27_lut_LC_22_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_27_lut_LC_22_22_1  (
            .in0(_gnd_net_),
            .in1(N__67933),
            .in2(N__59989),
            .in3(N__59956),
            .lcout(Add_add_temp_29),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15997 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15998 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_28_lut_LC_22_22_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_28_lut_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_28_lut_LC_22_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_28_lut_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(N__68965),
            .in2(N__59953),
            .in3(N__59935),
            .lcout(Add_add_temp_30),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15998 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15999 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_29_lut_LC_22_22_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_29_lut_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_29_lut_LC_22_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_29_lut_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(N__68910),
            .in2(N__60447),
            .in3(N__59932),
            .lcout(Add_add_temp_31),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15999 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n16000 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_30_lut_LC_22_22_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_30_lut_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_30_lut_LC_22_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_30_lut_LC_22_22_4  (
            .in0(_gnd_net_),
            .in1(N__60441),
            .in2(N__68839),
            .in3(N__59929),
            .lcout(Add_add_temp_32),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n16000 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n16001 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_31_lut_LC_22_22_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_31_lut_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_31_lut_LC_22_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_31_lut_LC_22_22_5  (
            .in0(_gnd_net_),
            .in1(N__60443),
            .in2(N__68770),
            .in3(N__59926),
            .lcout(Add_add_temp_33),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n16001 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n16002 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_32_lut_LC_22_22_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_32_lut_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_32_lut_LC_22_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_32_lut_LC_22_22_6  (
            .in0(_gnd_net_),
            .in1(N__68698),
            .in2(N__60448),
            .in3(N__60451),
            .lcout(Add_add_temp_34),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n16002 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n16003 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_33_lut_LC_22_22_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_33_lut_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_33_lut_LC_22_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_559_33_lut_LC_22_22_7  (
            .in0(N__60442),
            .in1(N__69045),
            .in2(_gnd_net_),
            .in3(N__60415),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Saturate_out1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i13263_4_lut_LC_22_23_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i13263_4_lut_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i13263_4_lut_LC_22_23_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i13263_4_lut_LC_22_23_0  (
            .in0(N__60556),
            .in1(N__60398),
            .in2(N__60375),
            .in3(N__60341),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n15200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_278_LC_22_23_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_278_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_278_LC_22_23_1 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_278_LC_22_23_1  (
            .in0(N__60321),
            .in1(N__60303),
            .in2(N__60292),
            .in3(N__60270),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20680_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_279_LC_22_23_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_279_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_279_LC_22_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_279_LC_22_23_2  (
            .in0(N__60251),
            .in1(N__60215),
            .in2(N__60199),
            .in3(N__60174),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_284_LC_22_23_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_284_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_284_LC_22_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_284_LC_22_23_3  (
            .in0(N__60111),
            .in1(N__60093),
            .in2(N__60147),
            .in3(N__60069),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_2_lut_LC_22_23_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_2_lut_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_2_lut_LC_22_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_2_lut_LC_22_23_4  (
            .in0(_gnd_net_),
            .in1(N__60140),
            .in2(_gnd_net_),
            .in3(N__60123),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20722_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_276_LC_22_23_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_276_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_276_LC_22_23_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_276_LC_22_23_5  (
            .in0(N__60110),
            .in1(N__60092),
            .in2(N__60079),
            .in3(N__60068),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n19761_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_277_LC_22_23_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_277_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_277_LC_22_23_6 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_277_LC_22_23_6  (
            .in0(N__62660),
            .in1(N__62687),
            .in2(N__60559),
            .in3(N__62714),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_22_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_22_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_22_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_2_lut_LC_22_25_0  (
            .in0(_gnd_net_),
            .in1(N__64914),
            .in2(N__64753),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n69 ),
            .ltout(),
            .carryin(bfn_22_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18234 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_22_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_22_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_22_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_3_lut_LC_22_25_1  (
            .in0(_gnd_net_),
            .in1(N__60550),
            .in2(N__64450),
            .in3(N__60535),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n115 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18234 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18235 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_22_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_22_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_22_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_4_lut_LC_22_25_2  (
            .in0(_gnd_net_),
            .in1(N__62629),
            .in2(N__64220),
            .in3(N__60523),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n164 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18235 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18236 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_22_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_22_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_22_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_5_lut_LC_22_25_3  (
            .in0(_gnd_net_),
            .in1(N__62620),
            .in2(N__63967),
            .in3(N__60511),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n213 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18236 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18237 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_22_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_22_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_22_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_6_lut_LC_22_25_4  (
            .in0(_gnd_net_),
            .in1(N__62611),
            .in2(N__63668),
            .in3(N__60499),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n262 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18237 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18238 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_22_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_22_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_22_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_7_lut_LC_22_25_5  (
            .in0(_gnd_net_),
            .in1(N__62602),
            .in2(N__63383),
            .in3(N__60484),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n311 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18238 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18239 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_22_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_22_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_22_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_8_lut_LC_22_25_6  (
            .in0(_gnd_net_),
            .in1(N__62593),
            .in2(N__63109),
            .in3(N__60469),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n360 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18239 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18240 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_22_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_22_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_22_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_9_lut_LC_22_25_7  (
            .in0(_gnd_net_),
            .in1(N__62584),
            .in2(N__66829),
            .in3(N__60454),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n409 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18240 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18241 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_22_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_22_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_22_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_10_lut_LC_22_26_0  (
            .in0(_gnd_net_),
            .in1(N__62575),
            .in2(N__66631),
            .in3(N__60664),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n458 ),
            .ltout(),
            .carryin(bfn_22_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18242 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_22_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_22_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_22_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_11_lut_LC_22_26_1  (
            .in0(_gnd_net_),
            .in1(N__62830),
            .in2(N__66349),
            .in3(N__60652),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n507 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18242 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18243 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_22_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_22_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_22_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_12_lut_LC_22_26_2  (
            .in0(_gnd_net_),
            .in1(N__62821),
            .in2(N__66086),
            .in3(N__60640),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n556 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18243 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_22_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_22_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_22_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_13_lut_LC_22_26_3  (
            .in0(_gnd_net_),
            .in1(N__62812),
            .in2(N__65828),
            .in3(N__60628),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n605 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18244 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_22_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_22_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_22_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_14_lut_LC_22_26_4  (
            .in0(_gnd_net_),
            .in1(N__62803),
            .in2(N__65596),
            .in3(N__60613),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n654 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18245 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_22_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_22_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_22_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_15_lut_LC_22_26_5  (
            .in0(_gnd_net_),
            .in1(N__65384),
            .in2(N__62794),
            .in3(N__60598),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n703 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18246 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_22_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_22_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_22_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_566_16_lut_LC_22_26_6  (
            .in0(_gnd_net_),
            .in1(N__65194),
            .in2(N__62782),
            .in3(N__60580),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n758 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18247 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_LUT4_0_LC_22_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_LUT4_0_LC_22_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_LUT4_0_LC_22_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_LUT4_0_LC_22_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60577),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n759_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_22_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_22_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_22_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_570_2_lut_LC_22_28_0  (
            .in0(_gnd_net_),
            .in1(N__64960),
            .in2(N__64758),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n78 ),
            .ltout(),
            .carryin(bfn_22_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18279 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_22_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_22_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_22_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_3_lut_LC_22_28_1  (
            .in0(_gnd_net_),
            .in1(N__60748),
            .in2(N__64496),
            .in3(N__60742),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n124 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18279 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18280 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_22_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_22_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_22_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_4_lut_LC_22_28_2  (
            .in0(_gnd_net_),
            .in1(N__60739),
            .in2(N__64243),
            .in3(N__60733),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n173 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18280 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18281 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_22_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_22_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_22_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_5_lut_LC_22_28_3  (
            .in0(_gnd_net_),
            .in1(N__60730),
            .in2(N__63979),
            .in3(N__60724),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n222 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18281 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18282 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_22_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_22_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_22_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_6_lut_LC_22_28_4  (
            .in0(_gnd_net_),
            .in1(N__60721),
            .in2(N__63669),
            .in3(N__60715),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n271 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18282 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18283 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_22_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_22_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_22_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_7_lut_LC_22_28_5  (
            .in0(_gnd_net_),
            .in1(N__60712),
            .in2(N__63405),
            .in3(N__60706),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n320 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18283 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18284 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_22_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_22_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_22_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_8_lut_LC_22_28_6  (
            .in0(_gnd_net_),
            .in1(N__60703),
            .in2(N__63131),
            .in3(N__60697),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n369 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18284 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18285 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_22_28_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_22_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_22_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_9_lut_LC_22_28_7  (
            .in0(_gnd_net_),
            .in1(N__66922),
            .in2(N__60694),
            .in3(N__60685),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n418 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18285 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18286 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_22_29_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_22_29_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_22_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_10_lut_LC_22_29_0  (
            .in0(_gnd_net_),
            .in1(N__60682),
            .in2(N__66640),
            .in3(N__60676),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n467 ),
            .ltout(),
            .carryin(bfn_22_29_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18287 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_22_29_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_22_29_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_22_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_11_lut_LC_22_29_1  (
            .in0(_gnd_net_),
            .in1(N__61063),
            .in2(N__66361),
            .in3(N__61057),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n516 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18287 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18288 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_22_29_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_22_29_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_22_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_12_lut_LC_22_29_2  (
            .in0(_gnd_net_),
            .in1(N__61054),
            .in2(N__66098),
            .in3(N__61048),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n565 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18288 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18289 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_22_29_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_22_29_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_22_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_13_lut_LC_22_29_3  (
            .in0(_gnd_net_),
            .in1(N__61045),
            .in2(N__65844),
            .in3(N__61039),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n614 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18289 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18290 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_22_29_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_22_29_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_22_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_14_lut_LC_22_29_4  (
            .in0(_gnd_net_),
            .in1(N__61036),
            .in2(N__65611),
            .in3(N__61030),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n663 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18290 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18291 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_22_29_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_22_29_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_22_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_15_lut_LC_22_29_5  (
            .in0(_gnd_net_),
            .in1(N__65388),
            .in2(N__61027),
            .in3(N__61018),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n712 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18291 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18292 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_22_29_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_22_29_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_22_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_16_lut_LC_22_29_6  (
            .in0(_gnd_net_),
            .in1(N__65201),
            .in2(N__61015),
            .in3(N__60991),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n770 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18292 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_LUT4_0_LC_22_29_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_LUT4_0_LC_22_29_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_LUT4_0_LC_22_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_LUT4_0_LC_22_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60988),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n771_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_23_11_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_23_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_2_lut_LC_23_11_0  (
            .in0(_gnd_net_),
            .in1(N__60939),
            .in2(N__67456),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_1 ),
            .ltout(),
            .carryin(bfn_23_11_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17521 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_23_11_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_23_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_3_lut_LC_23_11_1  (
            .in0(_gnd_net_),
            .in1(N__67413),
            .in2(N__61150),
            .in3(N__61141),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_2 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17521 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17522 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_23_11_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_23_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_4_lut_LC_23_11_2  (
            .in0(_gnd_net_),
            .in1(N__61138),
            .in2(N__67457),
            .in3(N__61132),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_3 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17522 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17523 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_23_11_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_23_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_5_lut_LC_23_11_3  (
            .in0(_gnd_net_),
            .in1(N__67417),
            .in2(N__61129),
            .in3(N__61120),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_4 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17523 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17524 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_23_11_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_23_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_6_lut_LC_23_11_4  (
            .in0(_gnd_net_),
            .in1(N__61117),
            .in2(N__67458),
            .in3(N__61111),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_5 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17524 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17525 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_23_11_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_23_11_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_23_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_7_lut_LC_23_11_5  (
            .in0(_gnd_net_),
            .in1(N__67421),
            .in2(N__61108),
            .in3(N__61099),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_6 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17525 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17526 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_23_11_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_23_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_8_lut_LC_23_11_6  (
            .in0(_gnd_net_),
            .in1(N__61096),
            .in2(N__67459),
            .in3(N__61090),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_7 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17526 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17527 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_23_11_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_23_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_9_lut_LC_23_11_7  (
            .in0(_gnd_net_),
            .in1(N__67425),
            .in2(N__61087),
            .in3(N__61078),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_8 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17527 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17528 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_23_12_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_23_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_10_lut_LC_23_12_0  (
            .in0(_gnd_net_),
            .in1(N__67426),
            .in2(N__61075),
            .in3(N__61066),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_9 ),
            .ltout(),
            .carryin(bfn_23_12_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17529 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_23_12_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_23_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_11_lut_LC_23_12_1  (
            .in0(_gnd_net_),
            .in1(N__61288),
            .in2(N__67460),
            .in3(N__61282),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_10 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17529 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17530 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_23_12_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_23_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_12_lut_LC_23_12_2  (
            .in0(_gnd_net_),
            .in1(N__61279),
            .in2(N__67463),
            .in3(N__61273),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_11 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17530 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17531 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_23_12_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_23_12_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_23_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_13_lut_LC_23_12_3  (
            .in0(_gnd_net_),
            .in1(N__61270),
            .in2(N__67461),
            .in3(N__61264),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_12 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17531 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17532 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_23_12_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_23_12_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_23_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_14_lut_LC_23_12_4  (
            .in0(_gnd_net_),
            .in1(N__61261),
            .in2(N__67464),
            .in3(N__61255),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17532 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17533 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_23_12_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_23_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_15_lut_LC_23_12_5  (
            .in0(_gnd_net_),
            .in1(N__61252),
            .in2(N__67462),
            .in3(N__61246),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Proportional_Gain_mul_temp_14 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17533 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n17534 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_23_12_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_23_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.paramCurrentControlP_15__I_0_add_561_16_lut_LC_23_12_6  (
            .in0(_gnd_net_),
            .in1(N__61243),
            .in2(N__61213),
            .in3(N__61183),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n738 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n17534 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_LUT4_0_LC_23_12_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_LUT4_0_LC_23_12_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_LUT4_0_LC_23_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_LUT4_0_LC_23_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61180),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n739_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_20_LC_23_13_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_20_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_20_LC_23_13_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_20_LC_23_13_0  (
            .in0(N__69253),
            .in1(N__69204),
            .in2(N__69298),
            .in3(N__66976),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19932 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_LC_23_13_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_LC_23_13_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_LC_23_13_7 .LUT_INIT=16'b1111001011001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_LC_23_13_7  (
            .in0(N__61388),
            .in1(N__69294),
            .in2(N__61476),
            .in3(N__69252),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13172_2_lut_3_lut_LC_23_14_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13172_2_lut_3_lut_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13172_2_lut_3_lut_LC_23_14_0 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13172_2_lut_3_lut_LC_23_14_0  (
            .in0(N__68728),
            .in1(_gnd_net_),
            .in2(N__61480),
            .in3(N__61387),
            .lcout(),
            .ltout(\foc.dVoltage_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_122_LC_23_14_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_122_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_122_LC_23_14_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_122_LC_23_14_1  (
            .in0(N__68106),
            .in1(N__68727),
            .in2(N__61507),
            .in3(N__61486),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_125_LC_23_14_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_125_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_125_LC_23_14_2 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_125_LC_23_14_2  (
            .in0(N__61492),
            .in1(N__68049),
            .in2(N__61504),
            .in3(N__61318),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.equal_13243_i14_2_lut_3_lut_3_lut_LC_23_14_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.equal_13243_i14_2_lut_3_lut_3_lut_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.equal_13243_i14_2_lut_3_lut_3_lut_LC_23_14_3 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.equal_13243_i14_2_lut_3_lut_3_lut_LC_23_14_3  (
            .in0(N__61382),
            .in1(N__68464),
            .in2(_gnd_net_),
            .in3(N__61469),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13165_2_lut_3_lut_LC_23_14_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13165_2_lut_3_lut_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13165_2_lut_3_lut_LC_23_14_5 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13165_2_lut_3_lut_LC_23_14_5  (
            .in0(N__68107),
            .in1(_gnd_net_),
            .in2(N__61390),
            .in3(N__61470),
            .lcout(\foc.dVoltage_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13166_2_lut_3_lut_LC_23_14_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13166_2_lut_3_lut_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13166_2_lut_3_lut_LC_23_14_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13166_2_lut_3_lut_LC_23_14_6  (
            .in0(N__61471),
            .in1(N__68050),
            .in2(_gnd_net_),
            .in3(N__61386),
            .lcout(\foc.dVoltage_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_53_LC_23_15_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_53_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_53_LC_23_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_53_LC_23_15_0  (
            .in0(N__66949),
            .in1(N__68550),
            .in2(N__69155),
            .in3(N__68601),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_LC_23_15_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_LC_23_15_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_3_lut_LC_23_15_3  (
            .in0(N__67678),
            .in1(N__67732),
            .in2(_gnd_net_),
            .in3(N__67783),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_3_lut_LC_23_15_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_3_lut_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_3_lut_LC_23_15_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_3_lut_LC_23_15_5  (
            .in0(N__69203),
            .in1(N__69251),
            .in2(_gnd_net_),
            .in3(N__69293),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1202_3_lut_LC_23_16_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1202_3_lut_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1202_3_lut_LC_23_16_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1202_3_lut_LC_23_16_0  (
            .in0(N__67673),
            .in1(N__67728),
            .in2(_gnd_net_),
            .in3(N__67779),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_11_LC_23_16_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_11_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_11_LC_23_16_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_11_LC_23_16_1  (
            .in0(N__67610),
            .in1(N__68459),
            .in2(N__61510),
            .in3(N__67548),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i10_LC_23_16_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i10_LC_23_16_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i10_LC_23_16_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i10_LC_23_16_2  (
            .in0(N__62395),
            .in1(N__62017),
            .in2(_gnd_net_),
            .in3(N__61888),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62115),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i11_LC_23_16_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i11_LC_23_16_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i11_LC_23_16_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i11_LC_23_16_3  (
            .in0(N__62018),
            .in1(N__61891),
            .in2(_gnd_net_),
            .in3(N__61738),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62115),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i8_LC_23_16_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i8_LC_23_16_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i8_LC_23_16_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i8_LC_23_16_4  (
            .in0(N__62347),
            .in1(N__61890),
            .in2(_gnd_net_),
            .in3(N__62021),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62115),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i13_LC_23_16_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i13_LC_23_16_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i13_LC_23_16_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i13_LC_23_16_6  (
            .in0(N__61783),
            .in1(N__62019),
            .in2(_gnd_net_),
            .in3(N__61889),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62115),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i7_LC_23_16_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i7_LC_23_16_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i7_LC_23_16_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i7_LC_23_16_7  (
            .in0(N__62020),
            .in1(N__61892),
            .in2(_gnd_net_),
            .in3(N__62443),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62115),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i26_LC_23_17_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i26_LC_23_17_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i26_LC_23_17_0 .LUT_INIT=16'b1100111011001110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i26_LC_23_17_0  (
            .in0(N__61656),
            .in1(N__61886),
            .in2(N__62015),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i28_LC_23_17_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i28_LC_23_17_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i28_LC_23_17_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i28_LC_23_17_1  (
            .in0(N__61686),
            .in1(N__61885),
            .in2(_gnd_net_),
            .in3(N__61981),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i9_LC_23_17_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i9_LC_23_17_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i9_LC_23_17_2 .LUT_INIT=16'b1100111011001110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i9_LC_23_17_2  (
            .in0(N__62371),
            .in1(N__61887),
            .in2(N__62016),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i17_LC_23_17_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i17_LC_23_17_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i17_LC_23_17_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i17_LC_23_17_3  (
            .in0(N__62230),
            .in1(N__61884),
            .in2(_gnd_net_),
            .in3(N__61977),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i747_4_lut_LC_23_17_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i747_4_lut_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i747_4_lut_LC_23_17_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i747_4_lut_LC_23_17_4  (
            .in0(N__61717),
            .in1(N__61687),
            .in2(N__61660),
            .in3(N__61636),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_147_LC_23_17_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_147_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_147_LC_23_17_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_147_LC_23_17_5  (
            .in0(N__62143),
            .in1(N__61630),
            .in2(N__61600),
            .in3(N__61596),
            .lcout(Saturate_out1_31__N_266),
            .ltout(Saturate_out1_31__N_266_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i12_LC_23_17_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i12_LC_23_17_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i12_LC_23_17_6 .LUT_INIT=16'b0000111000001110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i12_LC_23_17_6  (
            .in0(N__61975),
            .in1(N__61762),
            .in2(N__61564),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i15_LC_23_17_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i15_LC_23_17_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i15_LC_23_17_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i15_LC_23_17_7  (
            .in0(N__62254),
            .in1(N__61883),
            .in2(_gnd_net_),
            .in3(N__61976),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62107),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i16_LC_23_18_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i16_LC_23_18_0 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i16_LC_23_18_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i16_LC_23_18_0  (
            .in0(N__61894),
            .in1(N__62023),
            .in2(_gnd_net_),
            .in3(N__62311),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i4_LC_23_18_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i4_LC_23_18_1 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i4_LC_23_18_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i4_LC_23_18_1  (
            .in0(N__62028),
            .in1(N__61899),
            .in2(_gnd_net_),
            .in3(N__62535),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i22_LC_23_18_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i22_LC_23_18_2 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i22_LC_23_18_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i22_LC_23_18_2  (
            .in0(N__61897),
            .in1(N__62026),
            .in2(_gnd_net_),
            .in3(N__61555),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i23_LC_23_18_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i23_LC_23_18_3 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i23_LC_23_18_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i23_LC_23_18_3  (
            .in0(N__62027),
            .in1(N__61898),
            .in2(_gnd_net_),
            .in3(N__61531),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i21_LC_23_18_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i21_LC_23_18_4 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i21_LC_23_18_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i21_LC_23_18_4  (
            .in0(N__61896),
            .in1(N__62025),
            .in2(_gnd_net_),
            .in3(N__62065),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i14_LC_23_18_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i14_LC_23_18_5 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i14_LC_23_18_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i14_LC_23_18_5  (
            .in0(N__62022),
            .in1(N__61893),
            .in2(_gnd_net_),
            .in3(N__62283),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i5_LC_23_18_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i5_LC_23_18_6 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i5_LC_23_18_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i5_LC_23_18_6  (
            .in0(N__61900),
            .in1(N__62029),
            .in2(_gnd_net_),
            .in3(N__62460),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i19_LC_23_18_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i19_LC_23_18_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i19_LC_23_18_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i19_LC_23_18_7  (
            .in0(N__62024),
            .in1(N__61895),
            .in2(_gnd_net_),
            .in3(N__62203),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62116),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_140_LC_23_19_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_140_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_140_LC_23_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_140_LC_23_19_0  (
            .in0(N__62483),
            .in1(N__62565),
            .in2(N__62517),
            .in3(N__62534),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_141_LC_23_19_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_141_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_141_LC_23_19_1 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_141_LC_23_19_1  (
            .in0(N__62459),
            .in1(N__62435),
            .in2(N__61798),
            .in3(N__62411),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i729_4_lut_LC_23_19_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i729_4_lut_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i729_4_lut_LC_23_19_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i729_4_lut_LC_23_19_2  (
            .in0(N__62367),
            .in1(N__62388),
            .in2(N__61795),
            .in3(N__62340),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n22_adj_519_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_142_LC_23_19_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_142_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_142_LC_23_19_3 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_142_LC_23_19_3  (
            .in0(N__61754),
            .in1(N__61776),
            .in2(N__61792),
            .in3(N__61731),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_133_LC_23_19_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_133_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_133_LC_23_19_5 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_133_LC_23_19_5  (
            .in0(N__62323),
            .in1(N__61775),
            .in2(N__61758),
            .in3(N__61730),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_130_LC_23_19_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_130_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_130_LC_23_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_2_lut_adj_130_LC_23_19_6  (
            .in0(_gnd_net_),
            .in1(N__62564),
            .in2(_gnd_net_),
            .in3(N__62547),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_131_LC_23_20_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_131_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_131_LC_23_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_131_LC_23_20_0  (
            .in0(N__62536),
            .in1(N__62516),
            .in2(N__62494),
            .in3(N__62467),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_132_LC_23_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_132_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_132_LC_23_20_1 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_132_LC_23_20_1  (
            .in0(N__62461),
            .in1(N__62436),
            .in2(N__62419),
            .in3(N__62415),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13268_4_lut_LC_23_20_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13268_4_lut_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i13268_4_lut_LC_23_20_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i13268_4_lut_LC_23_20_2  (
            .in0(N__62387),
            .in1(N__62366),
            .in2(N__62350),
            .in3(N__62339),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_134_LC_23_20_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_134_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_134_LC_23_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_134_LC_23_20_4  (
            .in0(N__62317),
            .in1(N__62300),
            .in2(N__62279),
            .in3(N__62243),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.n19746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_136_LC_23_20_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_136_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_136_LC_23_20_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.i1_4_lut_adj_136_LC_23_20_5  (
            .in0(N__62214),
            .in1(N__62190),
            .in2(N__62179),
            .in3(N__62165),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i31_LC_23_21_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i31_LC_23_21_7 .SEQ_MODE=4'b1000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i31_LC_23_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_i31_LC_23_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62130),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.currentControlITerm_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62119),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_285_LC_23_23_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_285_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_285_LC_23_23_2 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.i1_4_lut_adj_285_LC_23_23_2  (
            .in0(N__62731),
            .in1(N__62721),
            .in2(N__62698),
            .in3(N__62667),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n20718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_23_25_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_23_25_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_23_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_2_lut_LC_23_25_0  (
            .in0(_gnd_net_),
            .in1(N__64910),
            .in2(N__64754),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n72 ),
            .ltout(),
            .carryin(bfn_23_25_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_23_25_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_23_25_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_23_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_3_lut_LC_23_25_1  (
            .in0(_gnd_net_),
            .in1(N__62635),
            .in2(N__64451),
            .in3(N__62623),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n118 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18249 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18250 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_23_25_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_23_25_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_23_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_4_lut_LC_23_25_2  (
            .in0(_gnd_net_),
            .in1(N__64261),
            .in2(N__64241),
            .in3(N__62614),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n167 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18250 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_23_25_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_23_25_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_23_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_5_lut_LC_23_25_3  (
            .in0(_gnd_net_),
            .in1(N__64000),
            .in2(N__63980),
            .in3(N__62605),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n216 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18251 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_23_25_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_23_25_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_23_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_6_lut_LC_23_25_4  (
            .in0(_gnd_net_),
            .in1(N__63706),
            .in2(N__63686),
            .in3(N__62596),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n265 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18252 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_23_25_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_23_25_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_23_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_7_lut_LC_23_25_5  (
            .in0(_gnd_net_),
            .in1(N__63424),
            .in2(N__63384),
            .in3(N__62587),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n314 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18253 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_23_25_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_23_25_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_23_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_8_lut_LC_23_25_6  (
            .in0(_gnd_net_),
            .in1(N__63148),
            .in2(N__63136),
            .in3(N__62578),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n363 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18254 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_23_25_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_23_25_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_23_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_9_lut_LC_23_25_7  (
            .in0(_gnd_net_),
            .in1(N__62845),
            .in2(N__66830),
            .in3(N__62833),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n412 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18255 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18256 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_23_26_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_23_26_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_23_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_10_lut_LC_23_26_0  (
            .in0(_gnd_net_),
            .in1(N__66649),
            .in2(N__66639),
            .in3(N__62824),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n461 ),
            .ltout(),
            .carryin(bfn_23_26_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18257 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_23_26_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_23_26_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_23_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_11_lut_LC_23_26_1  (
            .in0(_gnd_net_),
            .in1(N__66379),
            .in2(N__66359),
            .in3(N__62815),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n510 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18257 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18258 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_23_26_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_23_26_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_23_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_12_lut_LC_23_26_2  (
            .in0(_gnd_net_),
            .in1(N__66118),
            .in2(N__66099),
            .in3(N__62806),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n559 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18258 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18259 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_23_26_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_23_26_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_23_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_13_lut_LC_23_26_3  (
            .in0(_gnd_net_),
            .in1(N__65863),
            .in2(N__65829),
            .in3(N__62797),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n608 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18259 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_23_26_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_23_26_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_23_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_14_lut_LC_23_26_4  (
            .in0(_gnd_net_),
            .in1(N__65629),
            .in2(N__65609),
            .in3(N__62785),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n657 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18260 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18261 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_23_26_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_23_26_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_23_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_15_lut_LC_23_26_5  (
            .in0(_gnd_net_),
            .in1(N__65385),
            .in2(N__65404),
            .in3(N__62773),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n706 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18261 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18262 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_23_26_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_23_26_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_23_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_567_16_lut_LC_23_26_6  (
            .in0(_gnd_net_),
            .in1(N__65202),
            .in2(N__65218),
            .in3(N__62755),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n762 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18262 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_LUT4_0_LC_23_26_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_LUT4_0_LC_23_26_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_LUT4_0_LC_23_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_LUT4_0_LC_23_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62752),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n763_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_23_27_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_23_27_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_23_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_569_2_lut_LC_23_27_0  (
            .in0(_gnd_net_),
            .in1(N__64956),
            .in2(N__64759),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n75 ),
            .ltout(),
            .carryin(bfn_23_27_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18264 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_23_27_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_23_27_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_23_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_3_lut_LC_23_27_1  (
            .in0(_gnd_net_),
            .in1(N__64507),
            .in2(N__64501),
            .in3(N__64252),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n121 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18264 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18265 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_23_27_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_23_27_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_23_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_4_lut_LC_23_27_2  (
            .in0(_gnd_net_),
            .in1(N__64249),
            .in2(N__64242),
            .in3(N__63991),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n170 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18265 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18266 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_23_27_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_23_27_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_23_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_5_lut_LC_23_27_3  (
            .in0(_gnd_net_),
            .in1(N__63988),
            .in2(N__63974),
            .in3(N__63697),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n219 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18266 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_23_27_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_23_27_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_23_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_6_lut_LC_23_27_4  (
            .in0(_gnd_net_),
            .in1(N__63694),
            .in2(N__63687),
            .in3(N__63415),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n268 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18267 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_23_27_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_23_27_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_23_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_7_lut_LC_23_27_5  (
            .in0(_gnd_net_),
            .in1(N__63412),
            .in2(N__63406),
            .in3(N__63139),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n317 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18268 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_23_27_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_23_27_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_23_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_8_lut_LC_23_27_6  (
            .in0(_gnd_net_),
            .in1(N__63110),
            .in2(N__62854),
            .in3(N__62836),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n366 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18269 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_23_27_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_23_27_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_23_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_9_lut_LC_23_27_7  (
            .in0(_gnd_net_),
            .in1(N__66937),
            .in2(N__66920),
            .in3(N__66643),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n415 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18270 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18271 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_23_28_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_23_28_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_23_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_10_lut_LC_23_28_0  (
            .in0(_gnd_net_),
            .in1(N__66598),
            .in2(N__66388),
            .in3(N__66370),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n464 ),
            .ltout(),
            .carryin(bfn_23_28_0_),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18272 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_23_28_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_23_28_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_23_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_11_lut_LC_23_28_1  (
            .in0(_gnd_net_),
            .in1(N__66367),
            .in2(N__66360),
            .in3(N__66109),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n513 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18272 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18273 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_23_28_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_23_28_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_23_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_12_lut_LC_23_28_2  (
            .in0(_gnd_net_),
            .in1(N__66106),
            .in2(N__66100),
            .in3(N__65854),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n562 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18273 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18274 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_23_28_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_23_28_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_23_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_13_lut_LC_23_28_3  (
            .in0(_gnd_net_),
            .in1(N__65851),
            .in2(N__65843),
            .in3(N__65620),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n611 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18274 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18275 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_23_28_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_23_28_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_23_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_14_lut_LC_23_28_4  (
            .in0(_gnd_net_),
            .in1(N__65617),
            .in2(N__65610),
            .in3(N__65392),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n660 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18275 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18276 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_23_28_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_23_28_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_23_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_15_lut_LC_23_28_5  (
            .in0(_gnd_net_),
            .in1(N__65389),
            .in2(N__65227),
            .in3(N__65206),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n709 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18276 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18277 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_23_28_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_23_28_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_23_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.Error_sub_temp_31__I_0_add_568_16_lut_LC_23_28_6  (
            .in0(_gnd_net_),
            .in1(N__65193),
            .in2(N__65038),
            .in3(N__67000),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n766 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_Q_Current_Control.n18277 ),
            .carryout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_LUT4_0_LC_23_28_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_LUT4_0_LC_23_28_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_LUT4_0_LC_23_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_LUT4_0_LC_23_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66997),
            .lcout(\foc.u_DQ_Current_Control.u_Q_Current_Control.n767_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_19_LC_24_14_4 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_19_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_19_LC_24_14_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_19_LC_24_14_4  (
            .in0(N__66964),
            .in1(N__68594),
            .in2(N__68549),
            .in3(N__68649),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_15_LC_24_14_6 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_15_LC_24_14_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_15_LC_24_14_6 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_15_LC_24_14_6  (
            .in0(N__67516),
            .in1(N__67964),
            .in2(N__67900),
            .in3(N__68942),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_17_LC_24_14_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_17_LC_24_14_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_17_LC_24_14_7 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_17_LC_24_14_7  (
            .in0(N__68862),
            .in1(N__68721),
            .in2(N__66967),
            .in3(N__68793),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n20098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13232_4_lut_LC_24_15_0 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13232_4_lut_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13232_4_lut_LC_24_15_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13232_4_lut_LC_24_15_0  (
            .in0(N__66943),
            .in1(N__68460),
            .in2(N__68179),
            .in3(N__67547),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13251_4_lut_LC_24_15_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13251_4_lut_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13251_4_lut_LC_24_15_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i13251_4_lut_LC_24_15_1  (
            .in0(N__68099),
            .in1(N__67970),
            .in2(N__66958),
            .in3(N__68047),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n15188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_LC_24_15_2 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_LC_24_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_LC_24_15_2  (
            .in0(N__68861),
            .in1(N__67885),
            .in2(N__66955),
            .in3(N__68936),
            .lcout(),
            .ltout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_27_LC_24_15_3 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_27_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_27_LC_24_15_3 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_27_LC_24_15_3  (
            .in0(N__68720),
            .in1(N__68792),
            .in2(N__66952),
            .in3(N__68648),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12921_2_lut_LC_24_15_5 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12921_2_lut_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12921_2_lut_LC_24_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i12921_2_lut_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(N__67611),
            .in2(_gnd_net_),
            .in3(N__67677),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n14851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_14_LC_24_15_7 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_14_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_14_LC_24_15_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.i1_4_lut_adj_14_LC_24_15_7  (
            .in0(N__68100),
            .in1(N__68048),
            .in2(N__68180),
            .in3(N__67522),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.u_Saturate_Output.n19690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_2_lut_LC_24_16_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_2_lut_LC_24_16_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_2_lut_LC_24_16_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_2_lut_LC_24_16_0  (
            .in0(N__67503),
            .in1(N__67485),
            .in2(N__67474),
            .in3(_gnd_net_),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20184 ),
            .ltout(),
            .carryin(bfn_24_16_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_3_lut_LC_24_16_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_3_lut_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_3_lut_LC_24_16_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_3_lut_LC_24_16_1  (
            .in0(N__67216),
            .in1(N__67203),
            .in2(N__67192),
            .in3(N__67177),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20186 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15568 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_4_lut_LC_24_16_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_4_lut_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_4_lut_LC_24_16_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_4_lut_LC_24_16_2  (
            .in0(N__67174),
            .in1(N__67161),
            .in2(N__67150),
            .in3(N__67135),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20188 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15569 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_5_lut_LC_24_16_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_5_lut_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_5_lut_LC_24_16_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_5_lut_LC_24_16_3  (
            .in0(N__67132),
            .in1(N__67116),
            .in2(N__67105),
            .in3(N__67090),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20190 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15570 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_6_lut_LC_24_16_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_6_lut_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_6_lut_LC_24_16_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_6_lut_LC_24_16_4  (
            .in0(N__67087),
            .in1(N__67077),
            .in2(N__67066),
            .in3(N__67051),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20192 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15571 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_lut_LC_24_16_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_lut_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_lut_LC_24_16_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_lut_LC_24_16_5  (
            .in0(N__67048),
            .in1(N__67032),
            .in2(N__67021),
            .in3(N__67003),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20194 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15572 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_0_LC_24_16_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_0_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_0_LC_24_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_0_LC_24_16_6  (
            .in0(_gnd_net_),
            .in1(N__68418),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_1_LC_24_16_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_1_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_1_LC_24_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_7_THRU_CRY_1_LC_24_16_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__68434),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_0_THRU_CO ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15573_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_8_lut_LC_24_17_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_8_lut_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_8_lut_LC_24_17_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_8_lut_LC_24_17_0  (
            .in0(N__67861),
            .in1(N__67855),
            .in2(N__67842),
            .in3(N__67825),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20196 ),
            .ltout(),
            .carryin(bfn_24_17_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_9_lut_LC_24_17_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_9_lut_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_9_lut_LC_24_17_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_9_lut_LC_24_17_1  (
            .in0(N__67822),
            .in1(N__67809),
            .in2(N__67798),
            .in3(N__67768),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.n20198 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15574 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_10_lut_LC_24_17_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_10_lut_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_10_lut_LC_24_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_10_lut_LC_24_17_2  (
            .in0(_gnd_net_),
            .in1(N__67758),
            .in2(N__67747),
            .in3(N__67717),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_9 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15575 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_11_lut_LC_24_17_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_11_lut_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_11_lut_LC_24_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_11_lut_LC_24_17_3  (
            .in0(_gnd_net_),
            .in1(N__67714),
            .in2(N__67695),
            .in3(N__67654),
            .lcout(\foc.preSatVoltage_10_adj_2311 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15576 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_12_lut_LC_24_17_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_12_lut_LC_24_17_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_12_lut_LC_24_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_12_lut_LC_24_17_4  (
            .in0(_gnd_net_),
            .in1(N__67650),
            .in2(N__67633),
            .in3(N__67591),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_11 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15577 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_13_lut_LC_24_17_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_13_lut_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_13_lut_LC_24_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_13_lut_LC_24_17_5  (
            .in0(_gnd_net_),
            .in1(N__67581),
            .in2(N__67570),
            .in3(N__67525),
            .lcout(\foc.preSatVoltage_12_adj_2330 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15578 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_lut_LC_24_17_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_lut_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_lut_LC_24_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_lut_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(N__68496),
            .in2(N__68479),
            .in3(N__68440),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_13 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15579 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_THRU_CRY_0_LC_24_17_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_THRU_CRY_0_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_THRU_CRY_0_LC_24_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_14_THRU_CRY_0_LC_24_17_7  (
            .in0(_gnd_net_),
            .in1(N__68422),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15580 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15580_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_15_lut_LC_24_18_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_15_lut_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_15_lut_LC_24_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_15_lut_LC_24_18_0  (
            .in0(_gnd_net_),
            .in1(N__68214),
            .in2(N__68203),
            .in3(N__68146),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_14 ),
            .ltout(),
            .carryin(bfn_24_18_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_16_lut_LC_24_18_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_16_lut_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_16_lut_LC_24_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_16_lut_LC_24_18_1  (
            .in0(_gnd_net_),
            .in1(N__68136),
            .in2(N__68125),
            .in3(N__68083),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_15 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15581 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_17_lut_LC_24_18_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_17_lut_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_17_lut_LC_24_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_17_lut_LC_24_18_2  (
            .in0(_gnd_net_),
            .in1(N__68076),
            .in2(N__68065),
            .in3(N__68020),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_16 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15582 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_18_lut_LC_24_18_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_18_lut_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_18_lut_LC_24_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_18_lut_LC_24_18_3  (
            .in0(_gnd_net_),
            .in1(N__68013),
            .in2(N__67996),
            .in3(N__67936),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_17 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15583 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_19_lut_LC_24_18_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_19_lut_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_19_lut_LC_24_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_19_lut_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__67929),
            .in2(N__67915),
            .in3(N__67864),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_18 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15584 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_20_lut_LC_24_18_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_20_lut_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_20_lut_LC_24_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_20_lut_LC_24_18_5  (
            .in0(_gnd_net_),
            .in1(N__68977),
            .in2(N__68961),
            .in3(N__68914),
            .lcout(\foc.preSatVoltage_19_adj_2329 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15585 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_21_lut_LC_24_18_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_21_lut_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_21_lut_LC_24_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_21_lut_LC_24_18_6  (
            .in0(_gnd_net_),
            .in1(N__68911),
            .in2(N__68890),
            .in3(N__68842),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_20 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15586 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_22_lut_LC_24_18_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_22_lut_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_22_lut_LC_24_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_22_lut_LC_24_18_7  (
            .in0(_gnd_net_),
            .in1(N__68829),
            .in2(N__68818),
            .in3(N__68773),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_21 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15587 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_23_lut_LC_24_19_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_23_lut_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_23_lut_LC_24_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_23_lut_LC_24_19_0  (
            .in0(_gnd_net_),
            .in1(N__68769),
            .in2(N__68746),
            .in3(N__68701),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_22 ),
            .ltout(),
            .carryin(bfn_24_19_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_24_lut_LC_24_19_1 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_24_lut_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_24_lut_LC_24_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_24_lut_LC_24_19_1  (
            .in0(_gnd_net_),
            .in1(N__68697),
            .in2(N__68674),
            .in3(N__68626),
            .lcout(\foc.preSatVoltage_23_adj_2328 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15589 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_25_lut_LC_24_19_2 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_25_lut_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_25_lut_LC_24_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_25_lut_LC_24_19_2  (
            .in0(_gnd_net_),
            .in1(N__69059),
            .in2(N__68623),
            .in3(N__68572),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_24 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15590 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_26_lut_LC_24_19_3 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_26_lut_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_26_lut_LC_24_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_26_lut_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(N__68569),
            .in2(N__69071),
            .in3(N__68518),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_25 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15591 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_27_lut_LC_24_19_4 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_27_lut_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_27_lut_LC_24_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_27_lut_LC_24_19_4  (
            .in0(_gnd_net_),
            .in1(N__69063),
            .in2(N__68515),
            .in3(N__69268),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_26 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15592 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_28_lut_LC_24_19_5 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_28_lut_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_28_lut_LC_24_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_28_lut_LC_24_19_5  (
            .in0(_gnd_net_),
            .in1(N__69265),
            .in2(N__69072),
            .in3(N__69226),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_27 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15593 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_29_lut_LC_24_19_6 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_29_lut_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_29_lut_LC_24_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_29_lut_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(N__69067),
            .in2(N__69223),
            .in3(N__69175),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_28 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15594 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_30_lut_LC_24_19_7 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_30_lut_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_30_lut_LC_24_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_30_lut_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(N__69172),
            .in2(N__69073),
            .in3(N__69130),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_29 ),
            .ltout(),
            .carryin(\foc.u_DQ_Current_Control.u_D_Current_Control.n15595 ),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_31_lut_LC_24_20_0 .C_ON=1'b1;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_31_lut_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_31_lut_LC_24_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_31_lut_LC_24_20_0  (
            .in0(_gnd_net_),
            .in1(N__69043),
            .in2(N__69127),
            .in3(N__69076),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.preSatVoltage_30 ),
            .ltout(),
            .carryin(bfn_24_20_0_),
            .carryout(\foc.u_DQ_Current_Control.u_D_Current_Control.n15597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_32_lut_LC_24_20_1 .C_ON=1'b0;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_32_lut_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_32_lut_LC_24_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \foc.u_DQ_Current_Control.u_D_Current_Control.add_547_32_lut_LC_24_20_1  (
            .in0(N__69044),
            .in1(N__69025),
            .in2(_gnd_net_),
            .in3(N__69013),
            .lcout(\foc.u_DQ_Current_Control.u_D_Current_Control.Voltage_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
