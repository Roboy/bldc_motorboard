-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 18:04:00

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46223\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.data_in_frame_0_3\ : std_logic;
signal \c0.n9186_cascade_\ : std_logic;
signal \c0.n8857_cascade_\ : std_logic;
signal \c0.n8725_cascade_\ : std_logic;
signal \c0.n8063_cascade_\ : std_logic;
signal \c0.n20_adj_2547_cascade_\ : std_logic;
signal \c0.n9317\ : std_logic;
signal \c0.n8063\ : std_logic;
signal \c0.n17650\ : std_logic;
signal \c0.n8645_cascade_\ : std_logic;
signal \c0.n9186\ : std_logic;
signal \c0.n30_adj_2489_cascade_\ : std_logic;
signal \c0.n18_adj_2545\ : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal \c0.n16405\ : std_logic;
signal \c0.n16406\ : std_logic;
signal \c0.n16407\ : std_logic;
signal \c0.n16408\ : std_logic;
signal \c0.n16409\ : std_logic;
signal \c0.n16410\ : std_logic;
signal \c0.n16411\ : std_logic;
signal \c0.data_out_frame2_0_0\ : std_logic;
signal data_out_frame2_7_2 : std_logic;
signal \c0.data_out_frame2_0_6\ : std_logic;
signal \c0.n18546_cascade_\ : std_logic;
signal data_out_frame2_11_5 : std_logic;
signal \c0.n18474\ : std_logic;
signal \c0.n18534_cascade_\ : std_logic;
signal data_out_frame2_17_5 : std_logic;
signal \c0.n18537_cascade_\ : std_logic;
signal \c0.n17803\ : std_logic;
signal \c0.n18080\ : std_logic;
signal \c0.n18384_cascade_\ : std_logic;
signal \c0.n22_adj_2523\ : std_logic;
signal \c0.n18387_cascade_\ : std_logic;
signal \c0.n5_adj_2463\ : std_logic;
signal data_out_frame2_16_5 : std_logic;
signal data_out_frame2_9_5 : std_logic;
signal data_out_frame2_6_2 : std_logic;
signal data_out_frame2_16_2 : std_logic;
signal \c0.n18486_cascade_\ : std_logic;
signal \c0.n18489_cascade_\ : std_logic;
signal \c0.n18084\ : std_logic;
signal \c0.n18366_cascade_\ : std_logic;
signal \c0.n6_adj_2466\ : std_logic;
signal \c0.n22_adj_2529\ : std_logic;
signal \c0.n18369_cascade_\ : std_logic;
signal data_out_frame2_7_5 : std_logic;
signal \c0.n5_adj_2503_cascade_\ : std_logic;
signal data_out_frame2_14_2 : std_logic;
signal \c0.n18606_cascade_\ : std_logic;
signal \c0.n18570_cascade_\ : std_logic;
signal \c0.n17779\ : std_logic;
signal \c0.n17773_cascade_\ : std_logic;
signal \c0.n18074\ : std_logic;
signal \c0.n18432_cascade_\ : std_logic;
signal \c0.n18435_cascade_\ : std_logic;
signal \c0.n17836\ : std_logic;
signal \c0.n18360_cascade_\ : std_logic;
signal \c0.n6_adj_2504\ : std_logic;
signal \c0.n18471_cascade_\ : std_logic;
signal \c0.n18363\ : std_logic;
signal \c0.n22_adj_2530_cascade_\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \c0.tx2.n16372\ : std_logic;
signal \c0.tx2.n16373\ : std_logic;
signal \c0.tx2.n16374\ : std_logic;
signal \c0.tx2.n16375\ : std_logic;
signal \c0.tx2.n16376\ : std_logic;
signal \c0.tx2.n16377\ : std_logic;
signal \c0.tx2.n16378\ : std_logic;
signal \c0.tx2.n16379\ : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal \c0.tx2.n17953\ : std_logic;
signal \c0.tx2.n18013\ : std_logic;
signal \c0.tx2.n17939\ : std_logic;
signal n316 : std_logic;
signal \c0.n17507_cascade_\ : std_logic;
signal \c0.data_in_frame_0_4\ : std_logic;
signal \c0.n17507\ : std_logic;
signal \c0.n17476_cascade_\ : std_logic;
signal \c0.n17476\ : std_logic;
signal \c0.n17478_cascade_\ : std_logic;
signal \c0.n17629_cascade_\ : std_logic;
signal \c0.n16_adj_2546\ : std_logic;
signal \c0.n9254\ : std_logic;
signal \c0.n9254_cascade_\ : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.n8976\ : std_logic;
signal \c0.data_in_frame_1_3\ : std_logic;
signal \c0.n5_adj_2515\ : std_logic;
signal \c0.data_out_frame2_0_5\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal \c0.n2607\ : std_logic;
signal \c0.n17513\ : std_logic;
signal \c0.n2602\ : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal \c0.n9_adj_2500\ : std_logic;
signal \c0.n9_adj_2507\ : std_logic;
signal \c0.n17325_cascade_\ : std_logic;
signal \c0.n8_adj_2459_cascade_\ : std_logic;
signal \c0.n2604\ : std_logic;
signal \c0.n11_adj_2460\ : std_logic;
signal \c0.n9605\ : std_logic;
signal \c0.n9900\ : std_logic;
signal \c0.n17806\ : std_logic;
signal data_out_frame2_18_5 : std_logic;
signal data_out_frame2_13_2 : std_logic;
signal \c0.n18492\ : std_logic;
signal \c0.n17827\ : std_logic;
signal data_out_frame2_12_5 : std_logic;
signal \c0.n9043_cascade_\ : std_logic;
signal data_out_frame2_14_6 : std_logic;
signal data_out_frame2_10_6 : std_logic;
signal data_out_frame2_11_0 : std_logic;
signal data_out_frame2_6_6 : std_logic;
signal data_out_frame2_7_6 : std_logic;
signal data_out_frame2_8_5 : std_logic;
signal data_out_frame2_15_1 : std_logic;
signal data_out_frame2_11_6 : std_logic;
signal data_out_frame2_15_6 : std_logic;
signal data_out_frame2_5_2 : std_logic;
signal data_out_frame2_15_2 : std_logic;
signal data_out_frame2_15_0 : std_logic;
signal data_out_frame2_8_6 : std_logic;
signal \c0.n18564\ : std_logic;
signal data_out_frame2_16_1 : std_logic;
signal data_out_frame2_17_1 : std_logic;
signal data_out_frame2_18_0 : std_logic;
signal data_out_frame2_10_3 : std_logic;
signal data_out_frame2_14_4 : std_logic;
signal \c0.n5_adj_2495\ : std_logic;
signal data_out_frame2_5_5 : std_logic;
signal \c0.n6_adj_2496\ : std_logic;
signal data_out_frame2_11_3 : std_logic;
signal \c0.n17629\ : std_logic;
signal \c0.n8725\ : std_logic;
signal data_out_frame2_10_0 : std_logic;
signal data_out_frame2_17_0 : std_logic;
signal data_out_frame2_16_0 : std_logic;
signal \c0.n18600\ : std_logic;
signal data_out_frame2_5_0 : std_logic;
signal \c0.n5_adj_2477_cascade_\ : std_logic;
signal \c0.n6_adj_2436\ : std_logic;
signal data_out_frame2_18_1 : std_logic;
signal \c0.n18468\ : std_logic;
signal data_out_frame2_5_1 : std_logic;
signal data_out_frame2_10_2 : std_logic;
signal data_out_frame2_11_2 : std_logic;
signal data_out_frame2_12_0 : std_logic;
signal \c0.n17794\ : std_logic;
signal \c0.n18078\ : std_logic;
signal \c0.n18408_cascade_\ : std_logic;
signal \c0.n6_adj_2506\ : std_logic;
signal \c0.n18411_cascade_\ : std_logic;
signal data_out_frame2_18_6 : std_logic;
signal \c0.n18552_cascade_\ : std_logic;
signal \c0.n18555_cascade_\ : std_logic;
signal \c0.n22_adj_2521\ : std_logic;
signal n317 : std_logic;
signal n318 : std_logic;
signal n319 : std_logic;
signal n321 : std_logic;
signal \r_Clock_Count_0_adj_2634\ : std_logic;
signal \r_Clock_Count_2_adj_2632\ : std_logic;
signal \r_Clock_Count_4_adj_2630\ : std_logic;
signal \r_Clock_Count_3_adj_2631\ : std_logic;
signal \r_Clock_Count_5_adj_2629\ : std_logic;
signal \c0.tx2.n10_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \c0.tx2.r_Clock_Count_8\ : std_logic;
signal \c0.tx2.n16452\ : std_logic;
signal \c0.tx2.r_SM_Main_2_N_2323_1_cascade_\ : std_logic;
signal n320 : std_logic;
signal n10244 : std_logic;
signal \r_Clock_Count_1_adj_2633\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_2354\ : std_logic;
signal \c0.tx2.n12306_cascade_\ : std_logic;
signal \c0.n12_adj_2492\ : std_logic;
signal \c0.data_in_frame_0_7\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal \c0.n17553_cascade_\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal \c0.n17406_cascade_\ : std_logic;
signal data_in_frame_5_5 : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal \c0.data_in_frame_1_5\ : std_logic;
signal \n9419_cascade_\ : std_logic;
signal \c0.n25_adj_2491\ : std_logic;
signal \n1396_cascade_\ : std_logic;
signal \n2589_cascade_\ : std_logic;
signal n2589 : std_logic;
signal \c0.n18558\ : std_logic;
signal \c0.n17797\ : std_logic;
signal \c0.n17424\ : std_logic;
signal \c0.n17569\ : std_logic;
signal \c0.n10_adj_2505\ : std_logic;
signal \c0.n9028\ : std_logic;
signal \c0.n8061_cascade_\ : std_logic;
signal \c0.data_in_frame_6_4\ : std_logic;
signal n2595 : std_logic;
signal \c0.data_in_frame_0_0\ : std_logic;
signal \c0.n2839\ : std_logic;
signal \c0.n9151_cascade_\ : std_logic;
signal \c0.n17588_cascade_\ : std_logic;
signal data_in_frame_8_5 : std_logic;
signal \c0.n6_adj_2429\ : std_logic;
signal \c0.data_out_frame2_20_5\ : std_logic;
signal data_out_frame2_12_2 : std_logic;
signal data_out_frame2_13_1 : std_logic;
signal data_out_frame2_12_1 : std_logic;
signal data_out_frame2_7_0 : std_logic;
signal \n9606_cascade_\ : std_logic;
signal data_out_frame2_10_5 : std_logic;
signal data_out_frame2_13_5 : std_logic;
signal data_out_frame2_9_0 : std_logic;
signal data_out_frame2_6_1 : std_logic;
signal data_out_frame2_17_2 : std_logic;
signal data_out_frame2_5_7 : std_logic;
signal data_out_frame2_6_5 : std_logic;
signal data_out_frame2_6_0 : std_logic;
signal data_out_frame2_7_1 : std_logic;
signal data_out_frame2_16_6 : std_logic;
signal data_out_frame2_11_7 : std_logic;
signal data_out_frame2_9_1 : std_logic;
signal data_out_frame2_8_1 : std_logic;
signal \c0.n17833\ : std_logic;
signal data_out_frame2_19_0 : std_logic;
signal \c0.n18603\ : std_logic;
signal \c0.n22_adj_2510\ : std_logic;
signal data_out_frame2_14_7 : std_logic;
signal data_out_frame2_15_7 : std_logic;
signal data_out_frame2_12_7 : std_logic;
signal \c0.n18582_cascade_\ : std_logic;
signal data_out_frame2_13_7 : std_logic;
signal data_out_frame2_9_2 : std_logic;
signal data_out_frame2_8_2 : std_logic;
signal \c0.n18504\ : std_logic;
signal \c0.n17824\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.n18612_cascade_\ : std_logic;
signal \c0.tx2.n18615\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal data_out_frame2_17_6 : std_logic;
signal data_out_frame2_13_4 : std_logic;
signal \c0.n12\ : std_logic;
signal \c0.n11_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal \c0.tx2.n18450\ : std_logic;
signal \c0.tx2.n18453\ : std_logic;
signal data_out_frame2_5_3 : std_logic;
signal data_out_frame2_7_3 : std_logic;
signal \c0.n5_adj_2509\ : std_logic;
signal \c0.byte_transmit_counter2_5\ : std_logic;
signal \c0.byte_transmit_counter2_6\ : std_logic;
signal \c0.n18_adj_2544_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_7\ : std_logic;
signal \c0.n19_adj_2540_cascade_\ : std_logic;
signal \c0.tx2_transmit_N_2287\ : std_logic;
signal \c0.tx2_transmit_N_2287_cascade_\ : std_logic;
signal \c0.n19_adj_2540\ : std_logic;
signal \c0.n67_cascade_\ : std_logic;
signal \c0.n13530\ : std_logic;
signal \c0.n17656\ : std_logic;
signal \c0.n20_adj_2427\ : std_logic;
signal \c0.n10_adj_2428_cascade_\ : std_logic;
signal \c0.n17442\ : std_logic;
signal \c0.n17553\ : std_logic;
signal \c0.n17442_cascade_\ : std_logic;
signal \c0.n17550\ : std_logic;
signal \c0.data_in_frame_4_0\ : std_logic;
signal \c0.n8874\ : std_logic;
signal \c0.data_in_frame_1_4\ : std_logic;
signal \c0.n8874_cascade_\ : std_logic;
signal \c0.n9349\ : std_logic;
signal \c0.n9368_cascade_\ : std_logic;
signal \c0.n23_adj_2426\ : std_logic;
signal \c0.data_in_frame_1_6\ : std_logic;
signal \c0.n17632\ : std_logic;
signal \c0.n17485\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal \c0.n17406\ : std_logic;
signal \c0.n12_adj_2449_cascade_\ : std_logic;
signal n2598 : std_logic;
signal \c0.n23_adj_2462\ : std_logic;
signal \c0.n24_adj_2454_cascade_\ : std_logic;
signal data_in_frame_5_3 : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal \c0.data_in_frame_7_7\ : std_logic;
signal n2584 : std_logic;
signal \c0.n9151\ : std_logic;
signal \n2584_cascade_\ : std_logic;
signal \c0.n21_adj_2465\ : std_logic;
signal n9419 : std_logic;
signal \c0.n8061\ : std_logic;
signal \c0.n8857\ : std_logic;
signal \c0.n18_adj_2468\ : std_logic;
signal \c0.n26_adj_2469_cascade_\ : std_logic;
signal \c0.n30\ : std_logic;
signal data_out_frame2_6_7 : std_logic;
signal \c0.n5_adj_2501\ : std_logic;
signal \c0.n17534\ : std_logic;
signal \c0.n8674\ : std_logic;
signal \c0.n9163\ : std_logic;
signal \c0.n17470\ : std_logic;
signal n9148 : std_logic;
signal \n9148_cascade_\ : std_logic;
signal \c0.n22_adj_2508\ : std_logic;
signal \c0.n12_adj_2542\ : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal \c0.n9058\ : std_logic;
signal \c0.n17467\ : std_logic;
signal \c0.data_in_frame_4_3\ : std_logic;
signal \c0.n17562\ : std_logic;
signal data_in_frame_8_7 : std_logic;
signal \c0.n17647_cascade_\ : std_logic;
signal \c0.n12_adj_2549\ : std_logic;
signal data_in_8_5 : std_logic;
signal \c0.n17602\ : std_logic;
signal \c0.n30_adj_2489\ : std_logic;
signal \c0.n9345\ : std_logic;
signal \c0.n9345_cascade_\ : std_logic;
signal \c0.n10_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_6\ : std_logic;
signal \c0.n17647\ : std_logic;
signal \c0.n8995\ : std_logic;
signal \c0.n6_adj_2550\ : std_logic;
signal \c0.data_out_frame2_20_0\ : std_logic;
signal \c0.n6_adj_2502_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_2\ : std_logic;
signal \c0.data_out_frame2_19_5\ : std_logic;
signal data_out_frame2_14_0 : std_logic;
signal data_out_frame2_18_2 : std_logic;
signal data_out_frame2_5_6 : std_logic;
signal data_out_frame2_6_3 : std_logic;
signal data_out_frame2_12_6 : std_logic;
signal data_out_frame2_13_6 : std_logic;
signal data_out_frame2_8_0 : std_logic;
signal data_out_frame2_10_7 : std_logic;
signal data_out_frame2_15_4 : std_logic;
signal data_out_frame2_12_4 : std_logic;
signal \c0.n17535_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_6\ : std_logic;
signal \c0.n9240\ : std_logic;
signal \c0.n9240_cascade_\ : std_logic;
signal \c0.n9131\ : std_logic;
signal \c0.n17409_cascade_\ : std_logic;
signal \c0.n10_adj_2470\ : std_logic;
signal \c0.data_out_frame2_20_1\ : std_logic;
signal \c0.data_out_frame2_19_1\ : std_logic;
signal \c0.n6_adj_2464\ : std_logic;
signal \c0.n18423_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal data_out_frame2_18_7 : std_logic;
signal \c0.data_out_frame2_19_7\ : std_logic;
signal \c0.n18576_cascade_\ : std_logic;
signal data_out_frame2_17_7 : std_logic;
signal \c0.n18579_cascade_\ : std_logic;
signal \c0.n22_adj_2520\ : std_logic;
signal \c0.n17788\ : std_logic;
signal \c0.n18420\ : std_logic;
signal \c0.n4_adj_2480\ : std_logic;
signal tx_enable : std_logic;
signal tx2_o : std_logic;
signal tx2_enable : std_logic;
signal \c0.tx2.n4\ : std_logic;
signal \c0.tx2.n9568_cascade_\ : std_logic;
signal \c0.tx2.tx2_active\ : std_logic;
signal \c0.tx2.n23\ : std_logic;
signal \c0.r_SM_Main_2_N_2326_0\ : std_logic;
signal \c0.tx2.n17990\ : std_logic;
signal \c0.tx2.r_SM_Main_2_N_2323_1\ : std_logic;
signal \c0.tx2.n12_cascade_\ : std_logic;
signal \r_SM_Main_2_adj_2628\ : std_logic;
signal \c0.tx2.r_SM_Main_0\ : std_logic;
signal \c0.tx2.r_SM_Main_1\ : std_logic;
signal \c0.tx2.n6812_cascade_\ : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.n17697_cascade_\ : std_logic;
signal data_in_0_4 : std_logic;
signal data_in_frame_5_0 : std_logic;
signal \c0.n9306\ : std_logic;
signal \c0.data_in_frame_1_2\ : std_logic;
signal \c0.data_in_frame_6_1\ : std_logic;
signal \c0.n9328\ : std_logic;
signal \c0.n8645\ : std_logic;
signal n9100 : std_logic;
signal \c0.data_in_frame_4_5\ : std_logic;
signal \c0.data_in_frame_0_5\ : std_logic;
signal \c0.data_in_frame_4_4\ : std_logic;
signal \c0.n9176\ : std_logic;
signal \c0.data_in_frame_4_2\ : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal \c0.n10_adj_2430_cascade_\ : std_logic;
signal \c0.data_in_frame_4_1\ : std_logic;
signal \c0.n8695_cascade_\ : std_logic;
signal \c0.n8867\ : std_logic;
signal \c0.data_in_frame_0_6\ : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal data_in_5_0 : std_logic;
signal data_in_7_6 : std_logic;
signal n2593 : std_logic;
signal \n2593_cascade_\ : std_logic;
signal \c0.n22_adj_2461\ : std_logic;
signal n2586 : std_logic;
signal \c0.n9279\ : std_logic;
signal \n2590_cascade_\ : std_logic;
signal \c0.n10_adj_2450\ : std_logic;
signal data_in_6_3 : std_logic;
signal n2596 : std_logic;
signal \c0.n17529\ : std_logic;
signal \n2596_cascade_\ : std_logic;
signal \c0.n10_adj_2498\ : std_logic;
signal \c0.data_in_frame_7_3\ : std_logic;
signal n2588 : std_logic;
signal \c0.n8687\ : std_logic;
signal n2585 : std_logic;
signal \c0.n17\ : std_logic;
signal n2590 : std_logic;
signal \c0.data_in_frame_7_1\ : std_logic;
signal \c0.data_in_frame_1_0\ : std_logic;
signal \c0.data_in_frame_4_6\ : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.data_in_frame_4_7\ : std_logic;
signal \c0.n17403\ : std_logic;
signal \c0.n17403_cascade_\ : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal n9283 : std_logic;
signal \n9283_cascade_\ : std_logic;
signal data_out_frame2_16_7 : std_logic;
signal \c0.n9219\ : std_logic;
signal \c0.n8695\ : std_logic;
signal \c0.data_in_frame_6_6\ : std_logic;
signal \c0.n9208\ : std_logic;
signal \c0.n22_cascade_\ : std_logic;
signal n16_adj_2656 : std_logic;
signal \c0.n17519\ : std_logic;
signal \c0.n24_cascade_\ : std_logic;
signal \c0.n11_adj_2453\ : std_logic;
signal data_in_frame_8_2 : std_logic;
signal data_in_frame_8_1 : std_logic;
signal \c0.data_in_frame_6_3\ : std_logic;
signal \c0.n17605\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.data_in_frame_7_6\ : std_logic;
signal \c0.n9144\ : std_logic;
signal \c0.n8064\ : std_logic;
signal \c0.n17582_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_7\ : std_logic;
signal n2560 : std_logic;
signal \c0.n17588\ : std_logic;
signal \c0.n17582\ : std_logic;
signal \n2560_cascade_\ : std_logic;
signal n17585 : std_logic;
signal \c0.n17648\ : std_logic;
signal \c0.n18_cascade_\ : std_logic;
signal \c0.n17418\ : std_logic;
signal n2572 : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \c0.tx.n16357\ : std_logic;
signal \c0.tx.n16358\ : std_logic;
signal \c0.tx.n16359\ : std_logic;
signal \c0.tx.n16360\ : std_logic;
signal \c0.tx.n16361\ : std_logic;
signal \c0.tx.n16362\ : std_logic;
signal \c0.tx.n16363\ : std_logic;
signal \c0.tx.n16364\ : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal \c0.n31\ : std_logic;
signal data_out_frame2_9_6 : std_logic;
signal data_out_frame2_15_3 : std_logic;
signal data_out_frame2_14_3 : std_logic;
signal \c0.n18516_cascade_\ : std_logic;
signal data_out_frame2_13_3 : std_logic;
signal data_out_frame2_11_1 : std_logic;
signal data_out_frame2_10_1 : std_logic;
signal \c0.n18480\ : std_logic;
signal \c0.n136\ : std_logic;
signal \c0.n1_adj_2443\ : std_logic;
signal \c0.n14631_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_2\ : std_logic;
signal \c0.n17482\ : std_logic;
signal data_out_frame2_9_3 : std_logic;
signal data_out_frame2_8_3 : std_logic;
signal \c0.n18522\ : std_logic;
signal \c0.data_out_frame2_0_7\ : std_logic;
signal \c0.n18076\ : std_logic;
signal data_out_frame2_9_7 : std_logic;
signal data_out_frame2_8_7 : std_logic;
signal \c0.n18588\ : std_logic;
signal \c0.n17785\ : std_logic;
signal \bfn_5_29_0_\ : std_logic;
signal n16319 : std_logic;
signal n16320 : std_logic;
signal n16321 : std_logic;
signal n16322 : std_logic;
signal n16323 : std_logic;
signal n16324 : std_logic;
signal n16325 : std_logic;
signal n16326 : std_logic;
signal \bfn_5_30_0_\ : std_logic;
signal n16327 : std_logic;
signal n16328 : std_logic;
signal n16329 : std_logic;
signal n16330 : std_logic;
signal n16331 : std_logic;
signal n16332 : std_logic;
signal n16333 : std_logic;
signal n16334 : std_logic;
signal \bfn_5_31_0_\ : std_logic;
signal n16335 : std_logic;
signal n16336 : std_logic;
signal n16337 : std_logic;
signal n16338 : std_logic;
signal n16339 : std_logic;
signal n16340 : std_logic;
signal n16341 : std_logic;
signal n16342 : std_logic;
signal \bfn_5_32_0_\ : std_logic;
signal n16343 : std_logic;
signal n16344 : std_logic;
signal n16345 : std_logic;
signal n16346 : std_logic;
signal n16347 : std_logic;
signal n16348 : std_logic;
signal n16349 : std_logic;
signal data_in_5_3 : std_logic;
signal \c0.n17715_cascade_\ : std_logic;
signal data_out_frame2_15_5 : std_logic;
signal \c0.n18540\ : std_logic;
signal \c0.data_in_1_0\ : std_logic;
signal \c0.data_in_0_0\ : std_logic;
signal data_in_3_7 : std_logic;
signal \c0.n6_adj_2473\ : std_logic;
signal data_in_8_0 : std_logic;
signal \c0.n81\ : std_logic;
signal data_in_6_0 : std_logic;
signal \c0.data_in_frame_6_0\ : std_logic;
signal n2599 : std_logic;
signal \n2599_cascade_\ : std_logic;
signal \c0.n20_adj_2452\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n12_adj_2472_cascade_\ : std_logic;
signal \c0.n17765\ : std_logic;
signal \c0.n8556_cascade_\ : std_logic;
signal \c0.n7_cascade_\ : std_logic;
signal \c0.n6_adj_2478\ : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.n8460\ : std_logic;
signal \c0.n17745\ : std_logic;
signal \c0.n16_adj_2485_cascade_\ : std_logic;
signal data_in_frame_10_6 : std_logic;
signal \n63_adj_2642_cascade_\ : std_logic;
signal n16468 : std_logic;
signal data_in_7_0 : std_logic;
signal \c0.n4_adj_2512_cascade_\ : std_logic;
signal n2591 : std_logic;
signal \c0.n8751\ : std_logic;
signal \c0.n17532\ : std_logic;
signal \n2591_cascade_\ : std_logic;
signal \c0.n9324\ : std_logic;
signal \c0.n17533\ : std_logic;
signal \c0.n2605\ : std_logic;
signal n2570 : std_logic;
signal \n2570_cascade_\ : std_logic;
signal \c0.n8556\ : std_logic;
signal \c0.n17_adj_2514_cascade_\ : std_logic;
signal \c0.data_in_frame_6_2\ : std_logic;
signal \FRAME_MATCHER_next_state_31_N_2026_1_cascade_\ : std_logic;
signal n2567 : std_logic;
signal \c0.n8658\ : std_logic;
signal data_in_frame_5_1 : std_logic;
signal \c0.n17516\ : std_logic;
signal \c0.n2601_cascade_\ : std_logic;
signal n2597 : std_logic;
signal \c0.n9039\ : std_logic;
signal \c0.n17522\ : std_logic;
signal \c0.n2606\ : std_logic;
signal \c0.n17428_cascade_\ : std_logic;
signal \c0.n11_adj_2494\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n17575\ : std_logic;
signal \c0.n9103\ : std_logic;
signal data_in_frame_5_2 : std_logic;
signal data_in_frame_5_6 : std_logic;
signal \c0.n17430\ : std_logic;
signal data_in_frame_5_4 : std_logic;
signal \c0.n2603\ : std_logic;
signal n2568 : std_logic;
signal \c0.n17538\ : std_logic;
signal \c0.n9355\ : std_logic;
signal \n2568_cascade_\ : std_logic;
signal \c0.n17541\ : std_logic;
signal \c0.n21_cascade_\ : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n27_cascade_\ : std_logic;
signal \c0.n5_adj_2438\ : std_logic;
signal \c0.data_in_frame_6_7\ : std_logic;
signal \c0.n4_adj_2548\ : std_logic;
signal data_in_frame_8_4 : std_logic;
signal n19_adj_2651 : std_logic;
signal data_in_frame_8_3 : std_logic;
signal n9380 : std_logic;
signal n9054 : std_logic;
signal \n6_adj_2604_cascade_\ : std_logic;
signal data_in_frame_7_0 : std_logic;
signal \c0.data_in_frame_1_7\ : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.n17614\ : std_logic;
signal \c0.n8666\ : std_logic;
signal data_out_frame2_14_1 : std_logic;
signal n18104 : std_logic;
signal n18097 : std_logic;
signal n18103 : std_logic;
signal data_in_7_3 : std_logic;
signal n18054 : std_logic;
signal data_out_frame2_10_4 : std_logic;
signal data_out_frame2_11_4 : std_logic;
signal data_out_frame2_14_5 : std_logic;
signal \c0.data_in_frame_10_0\ : std_logic;
signal \c0.n14631\ : std_logic;
signal data_out_frame2_12_3 : std_logic;
signal data_in_20_2 : std_logic;
signal \c0.n17815\ : std_logic;
signal \c0.n17818\ : std_logic;
signal \c0.n6_adj_2432\ : std_logic;
signal \c0.n18372_cascade_\ : std_logic;
signal \c0.n18375_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal data_out_frame2_18_3 : std_logic;
signal \c0.data_out_frame2_19_3\ : std_logic;
signal data_out_frame2_16_3 : std_logic;
signal \c0.n18510_cascade_\ : std_logic;
signal data_out_frame2_17_3 : std_logic;
signal \c0.data_out_frame2_20_3\ : std_logic;
signal \c0.n18513_cascade_\ : std_logic;
signal \c0.n22_adj_2527\ : std_logic;
signal n9652 : std_logic;
signal n9922 : std_logic;
signal \r_Bit_Index_2_adj_2635\ : std_logic;
signal \c0.n17559\ : std_logic;
signal n9135 : std_logic;
signal \c0.data_out_frame2_0_3\ : std_logic;
signal \c0.n18082\ : std_logic;
signal \r_Bit_Index_1_adj_2636\ : std_logic;
signal \r_Bit_Index_0_adj_2637\ : std_logic;
signal n4980 : std_logic;
signal \bfn_6_30_0_\ : std_logic;
signal n225 : std_logic;
signal \c0.rx.n16365\ : std_logic;
signal \c0.rx.n16366\ : std_logic;
signal \c0.rx.n16367\ : std_logic;
signal \c0.rx.n16368\ : std_logic;
signal \c0.rx.n16369\ : std_logic;
signal \c0.rx.n16370\ : std_logic;
signal \c0.rx.n16371\ : std_logic;
signal n224 : std_logic;
signal n226 : std_logic;
signal n221 : std_logic;
signal n223 : std_logic;
signal \c0.rx.n17999\ : std_logic;
signal \c0.n18444\ : std_logic;
signal \c0.n9\ : std_logic;
signal data_out_frame2_18_4 : std_logic;
signal \c0.data_out_frame2_19_4\ : std_logic;
signal data_out_frame2_16_4 : std_logic;
signal \c0.n18528_cascade_\ : std_logic;
signal data_out_frame2_17_4 : std_logic;
signal \c0.n134\ : std_logic;
signal \c0.n18531_cascade_\ : std_logic;
signal data_out_frame2_5_4 : std_logic;
signal \c0.n17955_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.data_out_frame2_0_4\ : std_logic;
signal \c0.n18456_cascade_\ : std_logic;
signal \c0.n18447\ : std_logic;
signal \c0.n18459_cascade_\ : std_logic;
signal \c0.n22_adj_2525\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.n15_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.tx2.n7727\ : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_4_7 : std_logic;
signal data_in_4_5 : std_logic;
signal data_in_3_5 : std_logic;
signal \c0.n28_adj_2475_cascade_\ : std_logic;
signal \c0.n8_adj_2474\ : std_logic;
signal \c0.n8559\ : std_logic;
signal \c0.data_in_2_0\ : std_logic;
signal data_in_0_1 : std_logic;
signal data_in_1_7 : std_logic;
signal data_in_2_5 : std_logic;
signal \c0.n17_adj_2486\ : std_logic;
signal \c0.data_in_1_3\ : std_logic;
signal \c0.data_in_0_3\ : std_logic;
signal data_in_4_3 : std_logic;
signal data_in_3_3 : std_logic;
signal \c0.data_in_frame_7_4\ : std_logic;
signal n2587 : std_logic;
signal \c0.data_in_7_4\ : std_logic;
signal \c0.data_in_6_4\ : std_logic;
signal data_in_5_4 : std_logic;
signal \c0.data_in_4_4\ : std_logic;
signal n17952 : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.data_in_3_4\ : std_logic;
signal \c0.n17743\ : std_logic;
signal data_in_4_0 : std_logic;
signal \c0.data_in_3_0\ : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_2_6 : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_9_1 : std_logic;
signal \c0.data_in_frame_7_5\ : std_logic;
signal data_in_frame_8_6 : std_logic;
signal \c0.n17473\ : std_logic;
signal \c0.data_in_4_6\ : std_logic;
signal data_in_frame_5_7 : std_logic;
signal \c0.n9368\ : std_logic;
signal \c0.n9365\ : std_logic;
signal \c0.n2600_cascade_\ : std_logic;
signal \c0.n9334\ : std_logic;
signal \c0.n10_adj_2493\ : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.n8572\ : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.n4_adj_2512\ : std_logic;
signal n2594 : std_logic;
signal \n2573_cascade_\ : std_logic;
signal n17481 : std_logic;
signal \c0.n9043\ : std_logic;
signal \c0.n8886\ : std_logic;
signal \c0.n15927\ : std_logic;
signal \c0.n17594\ : std_logic;
signal \c0.n17412\ : std_logic;
signal \n2565_cascade_\ : std_logic;
signal n2574 : std_logic;
signal n17547 : std_logic;
signal \c0.n23_cascade_\ : std_logic;
signal \c0.n17536\ : std_logic;
signal \c0.n28\ : std_logic;
signal data_in_frame_8_0 : std_logic;
signal data_in_frame_1_1 : std_logic;
signal \c0.data_in_frame_10_4\ : std_logic;
signal n2563 : std_logic;
signal \c0.data_in_frame_7_2\ : std_logic;
signal \c0.n8062\ : std_logic;
signal \n2563_cascade_\ : std_logic;
signal \c0.n9204\ : std_logic;
signal \c0.n8890\ : std_logic;
signal \c0.n17592_cascade_\ : std_logic;
signal \c0.n26\ : std_logic;
signal data_in_10_1 : std_logic;
signal \c0.n17544\ : std_logic;
signal \c0.n8056\ : std_logic;
signal \n2566_cascade_\ : std_logic;
signal n2561 : std_logic;
signal \c0.n19\ : std_logic;
signal data_in_9_0 : std_logic;
signal \c0.data_in_frame_9_0\ : std_logic;
signal n2575 : std_logic;
signal \c0.n17504\ : std_logic;
signal \c0.n6_adj_2541_cascade_\ : std_logic;
signal \c0.n17591\ : std_logic;
signal \c0.data_out_frame2_20_4\ : std_logic;
signal \c0.n17488\ : std_logic;
signal data_in_frame_9_6 : std_logic;
signal n17479 : std_logic;
signal n9051 : std_logic;
signal n6_adj_2583 : std_logic;
signal \c0.data_out_frame2_19_2\ : std_logic;
signal \c0.data_in_frame_0_1\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.data_in_frame_0_2\ : std_logic;
signal \c0.n10_adj_2536\ : std_logic;
signal n18101 : std_logic;
signal data_in_8_3 : std_logic;
signal \n8517_cascade_\ : std_logic;
signal n17366 : std_logic;
signal data_in_9_3 : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal \r_Clock_Count_3\ : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.tx.n10_cascade_\ : std_logic;
signal \r_Clock_Count_1\ : std_logic;
signal data_in_5_5 : std_logic;
signal data_in_19_0 : std_logic;
signal data_in_10_0 : std_logic;
signal rx_data_4 : std_logic;
signal data_in_15_2 : std_logic;
signal data_in_14_2 : std_logic;
signal data_in_4_2 : std_logic;
signal data_in_9_7 : std_logic;
signal data_in_8_7 : std_logic;
signal data_out_frame2_13_0 : std_logic;
signal data_in_18_5 : std_logic;
signal \n8562_cascade_\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.rx.n2_cascade_\ : std_logic;
signal \c0.rx.n2\ : std_logic;
signal \r_Clock_Count_0_adj_2624\ : std_logic;
signal \r_Clock_Count_1_adj_2623\ : std_logic;
signal \c0.rx.n79\ : std_logic;
signal \c0.rx.n18597\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \c0.rx.n13537\ : std_logic;
signal \c0.rx.n4_adj_2424\ : std_logic;
signal \c0.rx.n17381\ : std_logic;
signal \c0.rx.n18003_cascade_\ : std_logic;
signal \n13880_cascade_\ : std_logic;
signal \c0.rx.n10193\ : std_logic;
signal \r_Clock_Count_2_adj_2622\ : std_logic;
signal \c0.rx.n124\ : std_logic;
signal \r_Clock_Count_3_adj_2621\ : std_logic;
signal \c0.rx.n97_cascade_\ : std_logic;
signal \c0.rx.n17345\ : std_logic;
signal n13880 : std_logic;
signal n222 : std_logic;
signal \r_Clock_Count_4_adj_2620\ : std_logic;
signal n3 : std_logic;
signal \c0.rx.n18001\ : std_logic;
signal \n17856_cascade_\ : std_logic;
signal n17855 : std_logic;
signal \LED_c\ : std_logic;
signal \c0.rx.n112\ : std_logic;
signal data_out_frame2_7_4 : std_logic;
signal data_out_frame2_6_4 : std_logic;
signal \c0.n5_adj_2425\ : std_logic;
signal data_out_frame2_9_4 : std_logic;
signal data_out_frame2_8_4 : std_logic;
signal \c0.n8\ : std_logic;
signal \c0.data_out_frame2_0_1\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.n18086\ : std_logic;
signal data_in_10_7 : std_logic;
signal data_in_11_7 : std_logic;
signal data_in_12_7 : std_logic;
signal data_in_13_7 : std_logic;
signal data_in_14_7 : std_logic;
signal data_in_16_7 : std_logic;
signal data_in_15_7 : std_logic;
signal n2564 : std_logic;
signal data_in_14_1 : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_1_1 : std_logic;
signal data_in_13_1 : std_logic;
signal data_in_12_1 : std_logic;
signal data_in_11_1 : std_logic;
signal data_in_6_6 : std_logic;
signal data_in_5_6 : std_logic;
signal n9606 : std_logic;
signal data_out_frame2_7_7 : std_logic;
signal \c0.data_in_frame_9_7\ : std_logic;
signal \c0.n17433\ : std_logic;
signal data_in_7_7 : std_logic;
signal n2573 : std_logic;
signal \c0.data_in_frame_9_2\ : std_logic;
signal n2565 : std_logic;
signal \c0.data_in_frame_10_2\ : std_logic;
signal n2566 : std_logic;
signal n1396 : std_logic;
signal n2571 : std_logic;
signal \c0.data_in_frame_9_4\ : std_logic;
signal data_in_17_7 : std_logic;
signal n7364 : std_logic;
signal data_in_6_2 : std_logic;
signal data_in_5_2 : std_logic;
signal \c0.data_in_frame_10_5\ : std_logic;
signal n2562 : std_logic;
signal data_in_10_5 : std_logic;
signal data_in_9_5 : std_logic;
signal data_in_12_5 : std_logic;
signal data_in_11_5 : std_logic;
signal n18098 : std_logic;
signal \c0.n142\ : std_logic;
signal \c0.n1\ : std_logic;
signal \FRAME_MATCHER_next_state_1\ : std_logic;
signal \c0.FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n1_adj_2437\ : std_logic;
signal \r_SM_Main_2_N_2323_1_cascade_\ : std_logic;
signal \n17757_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_2\ : std_logic;
signal \c0.FRAME_MATCHER_state_1\ : std_logic;
signal \c0.n157\ : std_logic;
signal n18010 : std_logic;
signal n9390 : std_logic;
signal \n9390_cascade_\ : std_logic;
signal \n17681_cascade_\ : std_logic;
signal n16466 : std_logic;
signal n17356 : std_logic;
signal n18102 : std_logic;
signal \r_Clock_Count_2\ : std_logic;
signal n13601 : std_logic;
signal data_in_7_2 : std_logic;
signal n13597 : std_logic;
signal rx_data_6 : std_logic;
signal data_in_16_2 : std_logic;
signal n4 : std_logic;
signal rx_data_3 : std_logic;
signal n4_adj_2582 : std_logic;
signal data_in_20_6 : std_logic;
signal data_in_8_2 : std_logic;
signal n8567 : std_logic;
signal data_in_11_2 : std_logic;
signal data_in_13_2 : std_logic;
signal data_in_12_2 : std_logic;
signal \FRAME_MATCHER_next_state_31_N_2026_1\ : std_logic;
signal n63_adj_2642 : std_logic;
signal n63 : std_logic;
signal \FRAME_MATCHER_next_state_0\ : std_logic;
signal data_in_17_5 : std_logic;
signal \c0.rx.r_SM_Main_2_N_2386_0\ : std_logic;
signal \c0.rx.n18066\ : std_logic;
signal rand_data_0 : std_logic;
signal \bfn_9_29_0_\ : std_logic;
signal rand_data_1 : std_logic;
signal n16412 : std_logic;
signal rand_data_2 : std_logic;
signal n16413 : std_logic;
signal rand_data_3 : std_logic;
signal n16414 : std_logic;
signal rand_data_4 : std_logic;
signal n16415 : std_logic;
signal rand_data_5 : std_logic;
signal n16416 : std_logic;
signal rand_data_6 : std_logic;
signal rand_setpoint_6 : std_logic;
signal n16417 : std_logic;
signal rand_data_7 : std_logic;
signal rand_setpoint_7 : std_logic;
signal n16418 : std_logic;
signal n16419 : std_logic;
signal rand_data_8 : std_logic;
signal \bfn_9_30_0_\ : std_logic;
signal rand_data_9 : std_logic;
signal n16420 : std_logic;
signal rand_data_10 : std_logic;
signal n16421 : std_logic;
signal rand_data_11 : std_logic;
signal n16422 : std_logic;
signal rand_data_12 : std_logic;
signal n16423 : std_logic;
signal rand_data_13 : std_logic;
signal n16424 : std_logic;
signal rand_data_14 : std_logic;
signal n16425 : std_logic;
signal rand_data_15 : std_logic;
signal n16426 : std_logic;
signal n16427 : std_logic;
signal rand_data_16 : std_logic;
signal \bfn_9_31_0_\ : std_logic;
signal rand_data_17 : std_logic;
signal n16428 : std_logic;
signal rand_data_18 : std_logic;
signal n16429 : std_logic;
signal rand_data_19 : std_logic;
signal n16430 : std_logic;
signal rand_data_20 : std_logic;
signal n16431 : std_logic;
signal rand_data_21 : std_logic;
signal n16432 : std_logic;
signal rand_data_22 : std_logic;
signal n16433 : std_logic;
signal rand_data_23 : std_logic;
signal n16434 : std_logic;
signal n16435 : std_logic;
signal rand_data_24 : std_logic;
signal \bfn_9_32_0_\ : std_logic;
signal rand_data_25 : std_logic;
signal n16436 : std_logic;
signal rand_data_26 : std_logic;
signal n16437 : std_logic;
signal rand_data_27 : std_logic;
signal n16438 : std_logic;
signal rand_data_28 : std_logic;
signal n16439 : std_logic;
signal rand_data_29 : std_logic;
signal n16440 : std_logic;
signal rand_data_30 : std_logic;
signal n16441 : std_logic;
signal rand_data_31 : std_logic;
signal n16442 : std_logic;
signal data_in_1_5 : std_logic;
signal data_in_7_5 : std_logic;
signal data_in_6_5 : std_logic;
signal data_in_8_1 : std_logic;
signal \c0.data_in_7_1\ : std_logic;
signal data_in_10_3 : std_logic;
signal data_in_6_7 : std_logic;
signal data_in_5_7 : std_logic;
signal \c0.data_in_frame_10_1\ : std_logic;
signal \c0.data_in_frame_10_3\ : std_logic;
signal \c0.n6\ : std_logic;
signal data_in_11_0 : std_logic;
signal n7086 : std_logic;
signal data_in_15_1 : std_logic;
signal \c0.data_in_frame_9_1\ : std_logic;
signal \c0.data_in_frame_10_7\ : std_logic;
signal \c0.data_in_frame_9_5\ : std_logic;
signal \c0.data_in_frame_9_3\ : std_logic;
signal \c0.n8989\ : std_logic;
signal data_in_10_2 : std_logic;
signal data_in_9_2 : std_logic;
signal data_in_18_7 : std_logic;
signal rx_data_7 : std_logic;
signal data_in_16_3 : std_logic;
signal data_in_15_3 : std_logic;
signal data_in_20_7 : std_logic;
signal data_in_19_7 : std_logic;
signal n12123 : std_logic;
signal n7080 : std_logic;
signal n17767 : std_logic;
signal \c0.tx.n17\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal \n1_cascade_\ : std_logic;
signal \n3_adj_2650_cascade_\ : std_logic;
signal tx_o_adj_2584 : std_logic;
signal \c0.n17556_cascade_\ : std_logic;
signal data_in_1_4 : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_2_3 : std_logic;
signal data_in_3_2 : std_logic;
signal \c0.n16_adj_2513\ : std_logic;
signal data_in_18_0 : std_logic;
signal n9796 : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal n12_adj_2618 : std_logic;
signal n22 : std_logic;
signal n17950 : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal \c0.n6_adj_2448\ : std_logic;
signal data_in_19_6 : std_logic;
signal data_in_18_6 : std_logic;
signal rx_data_1 : std_logic;
signal rand_setpoint_2 : std_logic;
signal data_in_19_5 : std_logic;
signal rx_data_5 : std_logic;
signal data_in_20_5 : std_logic;
signal \c0.n17911\ : std_logic;
signal \c0.n5_adj_2488\ : std_logic;
signal \c0.n18498\ : std_logic;
signal \c0.n2_adj_2487_cascade_\ : std_logic;
signal n4_adj_2649 : std_logic;
signal n8562 : std_logic;
signal \n4_adj_2649_cascade_\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal rx_data_0 : std_logic;
signal data_in_20_0 : std_logic;
signal data_in_17_6 : std_logic;
signal data_in_16_6 : std_logic;
signal rand_setpoint_4 : std_logic;
signal data_in_15_6 : std_logic;
signal rand_setpoint_11 : std_logic;
signal rand_setpoint_25 : std_logic;
signal rand_setpoint_30 : std_logic;
signal rand_setpoint_31 : std_logic;
signal rand_setpoint_10 : std_logic;
signal \r_Clock_Count_5_adj_2619\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.n97\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2380_2_cascade_\ : std_logic;
signal \c0.rx.n18000_cascade_\ : std_logic;
signal \c0.rx.n18594\ : std_logic;
signal rand_setpoint_27 : std_logic;
signal \c0.n17966_cascade_\ : std_logic;
signal rand_setpoint_29 : std_logic;
signal \c0.n17970_cascade_\ : std_logic;
signal rand_setpoint_24 : std_logic;
signal \c0.n17957_cascade_\ : std_logic;
signal rand_setpoint_22 : std_logic;
signal data_in_19_2 : std_logic;
signal data_in_20_4 : std_logic;
signal data_in_19_4 : std_logic;
signal data_in_18_4 : std_logic;
signal data_in_18_2 : std_logic;
signal data_in_17_2 : std_logic;
signal data_in_8_4 : std_logic;
signal data_in_9_4 : std_logic;
signal data_in_10_4 : std_logic;
signal data_in_11_4 : std_logic;
signal data_in_12_4 : std_logic;
signal data_in_13_4 : std_logic;
signal data_in_14_4 : std_logic;
signal data_in_11_3 : std_logic;
signal data_in_15_4 : std_logic;
signal data_in_17_4 : std_logic;
signal data_in_16_4 : std_logic;
signal data_in_4_1 : std_logic;
signal \c0.n18089_cascade_\ : std_logic;
signal \c0.n18429_cascade_\ : std_logic;
signal \tx_data_7_N_keep\ : std_logic;
signal \c0.n18017_cascade_\ : std_logic;
signal \c0.n18426\ : std_logic;
signal data_in_17_3 : std_logic;
signal \c0.n5_adj_2499\ : std_logic;
signal \c0.n18378_cascade_\ : std_logic;
signal \c0.n18381_cascade_\ : std_logic;
signal \tx_data_2_N_keep\ : std_logic;
signal data_in_20_3 : std_logic;
signal data_in_13_5 : std_logic;
signal data_in_19_3 : std_logic;
signal data_in_18_3 : std_logic;
signal data_in_12_0 : std_logic;
signal data_in_12_3 : std_logic;
signal n18462 : std_logic;
signal n18465 : std_logic;
signal data_in_9_6 : std_logic;
signal data_in_8_6 : std_logic;
signal data_in_16_5 : std_logic;
signal data_in_14_3 : std_logic;
signal data_in_13_3 : std_logic;
signal \n17737_cascade_\ : std_logic;
signal n17312 : std_logic;
signal \n17312_cascade_\ : std_logic;
signal \n14_adj_2615_cascade_\ : std_logic;
signal data_in_17_1 : std_logic;
signal data_in_16_1 : std_logic;
signal n17757 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal data_in_18_1 : std_logic;
signal n18438 : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal n18441 : std_logic;
signal data_in_13_0 : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal data_in_20_1 : std_logic;
signal data_in_19_1 : std_logic;
signal data_in_17_0 : std_logic;
signal data_in_16_0 : std_logic;
signal \c0.n18501\ : std_logic;
signal \tx_data_0_N_keep_cascade_\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal data_in_15_5 : std_logic;
signal data_in_14_5 : std_logic;
signal n4958 : std_logic;
signal \r_Bit_Index_2_adj_2625\ : std_logic;
signal \n4958_cascade_\ : std_logic;
signal \n9920_cascade_\ : std_logic;
signal \r_Bit_Index_1_adj_2626\ : std_logic;
signal data_in_15_0 : std_logic;
signal data_in_14_0 : std_logic;
signal rand_setpoint_1 : std_logic;
signal rand_setpoint_0 : std_logic;
signal \c0.n8953_cascade_\ : std_logic;
signal rand_setpoint_5 : std_logic;
signal \c0.n5\ : std_logic;
signal \c0.n17972\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2380_2\ : std_logic;
signal \c0.rx.n17351\ : std_logic;
signal \c0.rx.r_SM_Main_0\ : std_logic;
signal \c0.rx.n17376\ : std_logic;
signal \c0.data_out_6__2__N_803_cascade_\ : std_logic;
signal rand_setpoint_18 : std_logic;
signal \c0.n2216_cascade_\ : std_logic;
signal \c0.data_out_6_2\ : std_logic;
signal rand_setpoint_26 : std_logic;
signal \c0.data_out_6__2__N_803\ : std_logic;
signal \c0.n17964_cascade_\ : std_logic;
signal \c0.n17525_cascade_\ : std_logic;
signal \c0.rx.n9553\ : std_logic;
signal \c0.rx.r_SM_Main_2\ : std_logic;
signal \c0.rx.r_SM_Main_1\ : std_logic;
signal \c0.data_in_6_1\ : std_logic;
signal data_in_5_1 : std_logic;
signal data_in_10_6 : std_logic;
signal data_in_11_6 : std_logic;
signal \c0.n17755\ : std_logic;
signal \c0.n25_adj_2517\ : std_logic;
signal \c0.n1314_cascade_\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \c0.n16305\ : std_logic;
signal \c0.n7273\ : std_logic;
signal \c0.n16306\ : std_logic;
signal \c0.n7272\ : std_logic;
signal \c0.n16307\ : std_logic;
signal \c0.n16308\ : std_logic;
signal \c0.n16309\ : std_logic;
signal \c0.n7269\ : std_logic;
signal \c0.n16310\ : std_logic;
signal \c0.n16311\ : std_logic;
signal \c0.n16312\ : std_logic;
signal \c0.n18011\ : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal \c0.n7266\ : std_logic;
signal \c0.n16313\ : std_logic;
signal \c0.n7265\ : std_logic;
signal \c0.n16314\ : std_logic;
signal \c0.n16315\ : std_logic;
signal \c0.n16316\ : std_logic;
signal \c0.n16317\ : std_logic;
signal \c0.n16318\ : std_logic;
signal \r_SM_Main_2_N_2323_1\ : std_logic;
signal \n4_adj_2653_cascade_\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.n17349\ : std_logic;
signal \c0.n17937\ : std_logic;
signal \c0.n18390_cascade_\ : std_logic;
signal \c0.n18393_cascade_\ : std_logic;
signal \tx_data_3_N_keep\ : std_logic;
signal \c0.n18095\ : std_logic;
signal n9646 : std_logic;
signal n9920 : std_logic;
signal \r_Bit_Index_0_adj_2627\ : std_logic;
signal \c0.data_out_6__7__N_675_cascade_\ : std_logic;
signal rand_setpoint_15 : std_logic;
signal \c0.n17928_cascade_\ : std_logic;
signal rand_setpoint_14 : std_logic;
signal \c0.n17465\ : std_logic;
signal \c0.n17906_cascade_\ : std_logic;
signal \c0.n17921\ : std_logic;
signal \c0.data_out_10_6\ : std_logic;
signal \c0.n2_adj_2483\ : std_logic;
signal \c0.n17389\ : std_logic;
signal \c0.n17389_cascade_\ : std_logic;
signal \c0.n17600_cascade_\ : std_logic;
signal \c0.n9658\ : std_logic;
signal \c0.n17398_cascade_\ : std_logic;
signal rand_setpoint_20 : std_logic;
signal \c0.n2146_cascade_\ : std_logic;
signal \c0.data_out_5__3__N_964\ : std_logic;
signal \c0.data_out_5__3__N_964_cascade_\ : std_logic;
signal \c0.data_out_6__3__N_785_cascade_\ : std_logic;
signal rand_setpoint_19 : std_logic;
signal \c0.n2181_cascade_\ : std_logic;
signal \data_out_6__6__N_729\ : std_logic;
signal data_out_2_0 : std_logic;
signal \data_out_6__7__N_678\ : std_logic;
signal \n96_cascade_\ : std_logic;
signal \n47_cascade_\ : std_logic;
signal n2615 : std_logic;
signal \n41_cascade_\ : std_logic;
signal n17958 : std_logic;
signal n43 : std_logic;
signal \c0.n7271\ : std_logic;
signal \c0.n18105\ : std_logic;
signal \c0.n18012\ : std_logic;
signal \c0.n17936\ : std_logic;
signal \c0.n7275\ : std_logic;
signal \c0.n7274\ : std_logic;
signal \c0.n18008\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal delay_counter_0 : std_logic;
signal delay_counter_13 : std_logic;
signal delay_counter_14 : std_logic;
signal \c0.n7264\ : std_logic;
signal \n29_cascade_\ : std_logic;
signal data_in_12_6 : std_logic;
signal \c0.n149_cascade_\ : std_logic;
signal \c0.n93\ : std_logic;
signal \n8529_cascade_\ : std_logic;
signal \c0.n8550_cascade_\ : std_logic;
signal n121_adj_2606 : std_logic;
signal n8529 : std_logic;
signal \n121_adj_2606_cascade_\ : std_logic;
signal n13_adj_2652 : std_logic;
signal \c0.n251\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \c0.n16350\ : std_logic;
signal \c0.n16351\ : std_logic;
signal \c0.n16352\ : std_logic;
signal \c0.n16353\ : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal \tx_transmit_N_2239_5\ : std_logic;
signal \c0.n16354\ : std_logic;
signal \c0.n16355\ : std_logic;
signal byte_transmit_counter_7 : std_logic;
signal \c0.n16356\ : std_logic;
signal \tx_transmit_N_2239_7\ : std_logic;
signal data_out_3_4 : std_logic;
signal \c0.n18093_cascade_\ : std_logic;
signal \c0.n18399_cascade_\ : std_logic;
signal \tx_transmit_N_2239_4\ : std_logic;
signal \c0.n5_adj_2447\ : std_logic;
signal \c0.n17941_cascade_\ : std_logic;
signal \c0.n18396\ : std_logic;
signal \c0.n18068\ : std_logic;
signal \c0.n5_adj_2490\ : std_logic;
signal \c0.data_out_10_4\ : std_logic;
signal \c0.n18067\ : std_logic;
signal \c0.n18092\ : std_logic;
signal \c0.n18094\ : std_logic;
signal \c0.n18096\ : std_logic;
signal \c0.n18088\ : std_logic;
signal \c0.n8634\ : std_logic;
signal \c0.n9276_cascade_\ : std_logic;
signal \c0.data_out_7__1__N_626\ : std_logic;
signal \c0.n17623_cascade_\ : std_logic;
signal rand_setpoint_8 : std_logic;
signal \c0.n17916_cascade_\ : std_logic;
signal \c0.data_out_7_0\ : std_logic;
signal \c0.n8486\ : std_logic;
signal \c0.n8486_cascade_\ : std_logic;
signal \c0.n16450\ : std_logic;
signal n4_adj_2612 : std_logic;
signal rand_setpoint_13 : std_logic;
signal \c0.n17925_cascade_\ : std_logic;
signal rand_setpoint_12 : std_logic;
signal \c0.n17931_cascade_\ : std_logic;
signal \c0.n17400\ : std_logic;
signal \c0.data_out_7__4__N_550\ : std_logic;
signal \c0.data_out_7_4\ : std_logic;
signal \data_out_5__4__N_959\ : std_logic;
signal rand_setpoint_28 : std_logic;
signal \c0.n17967_cascade_\ : std_logic;
signal \c0.n6_adj_2467\ : std_logic;
signal \c0.n9276\ : std_logic;
signal \c0.n17662_cascade_\ : std_logic;
signal rand_setpoint_23 : std_logic;
signal \c0.n2041_cascade_\ : std_logic;
signal \c0.n17974\ : std_logic;
signal rand_setpoint_16 : std_logic;
signal \c0.n17693_cascade_\ : std_logic;
signal \c0.data_out_6_0\ : std_logic;
signal data_out_1_7 : std_logic;
signal \c0.n17578\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal n96 : std_logic;
signal n6878 : std_logic;
signal \n17672_cascade_\ : std_logic;
signal \c0.n113\ : std_logic;
signal n17364 : std_logic;
signal \c0.n18009\ : std_logic;
signal \c0.delay_counter_12\ : std_logic;
signal n119 : std_logic;
signal \UART_TRANSMITTER_state_7_N_1749_2_cascade_\ : std_logic;
signal n18032 : std_logic;
signal n8488 : std_logic;
signal n17709 : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.n17753\ : std_logic;
signal n29 : std_logic;
signal \c0.n7268\ : std_logic;
signal \c0.n1314\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.delay_counter_11\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.n10_adj_2532_cascade_\ : std_logic;
signal \c0.n14_adj_2533\ : std_logic;
signal n17306 : std_logic;
signal \n17306_cascade_\ : std_logic;
signal \c0.n17387\ : std_logic;
signal \c0.n6_adj_2534\ : std_logic;
signal \tx_data_4_N_keep\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \c0.n16_adj_2445_cascade_\ : std_logic;
signal \c0.n19_adj_2446_cascade_\ : std_logic;
signal \c0.n8550\ : std_logic;
signal \c0.n2650\ : std_logic;
signal \c0.tx_transmit_N_2239_0\ : std_logic;
signal \c0.tx_transmit_N_2239_1\ : std_logic;
signal \tx_transmit_N_2239_2\ : std_logic;
signal \c0.n97\ : std_logic;
signal \c0.tx_transmit\ : std_logic;
signal tx_active : std_logic;
signal n13415 : std_logic;
signal \tx_transmit_N_2239_3\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal n16485 : std_logic;
signal \c0.n7428\ : std_logic;
signal n14_adj_2615 : std_logic;
signal n9631 : std_logic;
signal \tx_transmit_N_2239_6\ : std_logic;
signal byte_transmit_counter_6 : std_logic;
signal \c0.n149\ : std_logic;
signal \c0.n17741\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \c0.n18071\ : std_logic;
signal \c0.n8_adj_2526_cascade_\ : std_logic;
signal \c0.n18072\ : std_logic;
signal \c0.n17644\ : std_logic;
signal \c0.data_out_7__2__N_574\ : std_logic;
signal \c0.data_out_7__2__N_574_cascade_\ : std_logic;
signal \c0.data_out_10_2\ : std_logic;
signal \c0.data_out_9_2\ : std_logic;
signal \c0.data_out_9_3\ : std_logic;
signal \c0.n18073_cascade_\ : std_logic;
signal rand_setpoint_3 : std_logic;
signal data_out_8_2 : std_logic;
signal \c0.data_out_6_4\ : std_logic;
signal \c0.n9091_cascade_\ : std_logic;
signal \c0.n17566_cascade_\ : std_logic;
signal \c0.data_out_6_3\ : std_logic;
signal \c0.n9195_cascade_\ : std_logic;
signal \c0.data_out_7__4__N_556\ : std_logic;
signal \c0.n18015\ : std_logic;
signal \c0.n8_adj_2516\ : std_logic;
signal \c0.data_out_6_7\ : std_logic;
signal \c0.n9195\ : std_logic;
signal \c0.n17668_cascade_\ : std_logic;
signal \c0.n8812\ : std_logic;
signal \c0.n8_adj_2511_cascade_\ : std_logic;
signal \c0.n17623\ : std_logic;
signal \c0.n8950\ : std_logic;
signal \c0.data_out_9_0\ : std_logic;
signal \c0.data_out_10_0\ : std_logic;
signal \c0.n18016\ : std_logic;
signal \c0.data_out_2_3\ : std_logic;
signal \c0.n4_adj_2543_cascade_\ : std_logic;
signal rand_setpoint_21 : std_logic;
signal \c0.n9656_cascade_\ : std_logic;
signal rand_setpoint_17 : std_logic;
signal \c0.n2251_cascade_\ : std_logic;
signal \c0.n17962\ : std_logic;
signal \c0.data_out_6__1__N_849\ : std_logic;
signal \c0.data_out_1_1\ : std_logic;
signal data_out_1_2 : std_logic;
signal \c0.n8767_cascade_\ : std_logic;
signal \c0.n17525\ : std_logic;
signal \c0.n17641\ : std_logic;
signal \c0.n17457_cascade_\ : std_logic;
signal \c0.n8964\ : std_logic;
signal \c0.n17415\ : std_logic;
signal \c0.data_out_6__3__N_788\ : std_logic;
signal \c0.n17415_cascade_\ : std_logic;
signal \c0.data_out_5_2\ : std_logic;
signal rand_setpoint_9 : std_logic;
signal \c0.n9518\ : std_logic;
signal \data_out_6__2__N_804\ : std_logic;
signal \c0.n17457\ : std_logic;
signal \c0.n17654\ : std_logic;
signal \c0.n18061\ : std_logic;
signal \c0.data_out_7__5__N_543\ : std_logic;
signal \data_out_6__1__N_850\ : std_logic;
signal \c0.n2\ : std_logic;
signal \c0.n18060\ : std_logic;
signal data_out_0_5 : std_logic;
signal \c0.n18065_cascade_\ : std_logic;
signal \tx_data_5_N_keep\ : std_logic;
signal \c0.n18014\ : std_logic;
signal \tx_data_1_N_keep\ : std_logic;
signal \c0.n17943\ : std_logic;
signal \c0.n5_adj_2481_cascade_\ : std_logic;
signal \c0.n18091\ : std_logic;
signal \c0.n18402_cascade_\ : std_logic;
signal \c0.n2_adj_2476\ : std_logic;
signal \c0.n18405\ : std_logic;
signal \c0.data_out_5_1\ : std_logic;
signal \c0.n45_adj_2518_cascade_\ : std_logic;
signal \c0.n1_adj_2522\ : std_logic;
signal \c0.n46_cascade_\ : std_logic;
signal \c0.n44_adj_2524\ : std_logic;
signal \c0.n8_adj_2531\ : std_logic;
signal \c0.n18069_cascade_\ : std_logic;
signal \c0.n18070\ : std_logic;
signal rx_data_ready : std_logic;
signal data_in_14_6 : std_logic;
signal data_in_13_6 : std_logic;
signal \c0.n17445\ : std_logic;
signal \c0.n17510\ : std_logic;
signal \c0.data_out_9_1\ : std_logic;
signal data_out_8_1 : std_logic;
signal \c0.n8_adj_2519\ : std_logic;
signal \c0.n8_adj_2535\ : std_logic;
signal \c0.n17398\ : std_logic;
signal \c0.n9091\ : std_logic;
signal \c0.data_out_9_4\ : std_logic;
signal \c0.data_out_6_1\ : std_logic;
signal \c0.n17499\ : std_logic;
signal \c0.n6_adj_2451\ : std_logic;
signal \c0.data_out_10_5\ : std_logic;
signal \c0.n18064\ : std_logic;
signal \c0.n17668\ : std_logic;
signal \c0.n9087\ : std_logic;
signal \c0.n8_adj_2528_cascade_\ : std_logic;
signal \c0.data_out_10_1\ : std_logic;
signal \c0.n17556\ : std_logic;
signal \c0.data_out_6__7__N_675\ : std_logic;
signal \c0.data_out_10_7\ : std_logic;
signal \c0.n8600\ : std_logic;
signal \c0.data_out_5_3\ : std_logic;
signal \c0.n17635_cascade_\ : std_logic;
signal \c0.n17922\ : std_logic;
signal \c0.data_out_7__7__N_519\ : std_logic;
signal \c0.data_out_7_5\ : std_logic;
signal \c0.n17492\ : std_logic;
signal \c0.n17635\ : std_logic;
signal \c0.n17492_cascade_\ : std_logic;
signal \c0.data_out_10_3\ : std_logic;
signal \c0.data_out_7_2\ : std_logic;
signal \c0.n17600\ : std_logic;
signal \c0.data_out_9_6\ : std_logic;
signal \c0.data_out_7_1\ : std_logic;
signal \c0.n17454\ : std_logic;
signal \c0.data_out_6_5\ : std_logic;
signal \c0.data_out_6__5__N_752\ : std_logic;
signal \c0.n17454_cascade_\ : std_logic;
signal \c0.data_out_9_5\ : std_logic;
signal \c0.n8_adj_2537\ : std_logic;
signal \c0.n17626\ : std_logic;
signal \c0.n17608\ : std_logic;
signal \c0.n8970\ : std_logic;
signal \c0.n17662\ : std_logic;
signal data_out_8_6 : std_logic;
signal \c0.n17665\ : std_logic;
signal \c0.n12_adj_2482_cascade_\ : std_logic;
signal \c0.data_out_7_3\ : std_logic;
signal \data_out_10__7__N_114\ : std_logic;
signal \c0.data_out_9_7\ : std_logic;
signal data_out_8_7 : std_logic;
signal \c0.n8_adj_2538\ : std_logic;
signal \c0.data_out_0_6\ : std_logic;
signal data_out_0_3 : std_logic;
signal data_out_0_1 : std_logic;
signal data_out_0_0 : std_logic;
signal \c0.n8926\ : std_logic;
signal \c0.n8767\ : std_logic;
signal \c0.n8926_cascade_\ : std_logic;
signal n2720 : std_logic;
signal \UART_TRANSMITTER_state_0\ : std_logic;
signal n4430 : std_logic;
signal data_out_1_6 : std_logic;
signal data_out_3_5 : std_logic;
signal \UART_TRANSMITTER_state_1\ : std_logic;
signal n9519 : std_logic;
signal \data_out_5__7__N_931\ : std_logic;
signal \c0.data_out_6__4__N_765\ : std_logic;
signal \c0.n1_adj_2484\ : std_logic;
signal \c0.n18414_cascade_\ : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal \c0.n18417_cascade_\ : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal n7734 : std_logic;
signal \tx_data_6_N_keep_cascade_\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.data_out_7__6__N_530\ : std_logic;
signal \c0.n17949\ : std_logic;
signal data_out_3_6 : std_logic;
signal \c0.n18090\ : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.data_out_7_6\ : std_logic;
signal \c0.n5_adj_2444\ : std_logic;
signal \c0.n8_adj_2539\ : std_logic;
signal byte_transmit_counter_2 : std_logic;
signal \c0.n18062\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n18063\ : std_logic;
signal data_out_8_0 : std_logic;
signal \c0.data_out_7_7\ : std_logic;
signal \c0.n17638\ : std_logic;
signal n26 : std_logic;
signal \bfn_16_29_0_\ : std_logic;
signal n25 : std_logic;
signal n16380 : std_logic;
signal n24 : std_logic;
signal n16381 : std_logic;
signal n23 : std_logic;
signal n16382 : std_logic;
signal n22_adj_2655 : std_logic;
signal n16383 : std_logic;
signal n21 : std_logic;
signal n16384 : std_logic;
signal n20 : std_logic;
signal n16385 : std_logic;
signal n19 : std_logic;
signal n16386 : std_logic;
signal n16387 : std_logic;
signal n18 : std_logic;
signal \bfn_16_30_0_\ : std_logic;
signal n17 : std_logic;
signal n16388 : std_logic;
signal n16 : std_logic;
signal n16389 : std_logic;
signal n15 : std_logic;
signal n16390 : std_logic;
signal n14 : std_logic;
signal n16391 : std_logic;
signal n13 : std_logic;
signal n16392 : std_logic;
signal n12 : std_logic;
signal n16393 : std_logic;
signal n11 : std_logic;
signal n16394 : std_logic;
signal n16395 : std_logic;
signal n10 : std_logic;
signal \bfn_16_31_0_\ : std_logic;
signal n9 : std_logic;
signal n16396 : std_logic;
signal n8_adj_2617 : std_logic;
signal n16397 : std_logic;
signal n7 : std_logic;
signal n16398 : std_logic;
signal n6 : std_logic;
signal n16399 : std_logic;
signal blink_counter_21 : std_logic;
signal n16400 : std_logic;
signal blink_counter_22 : std_logic;
signal n16401 : std_logic;
signal blink_counter_23 : std_logic;
signal n16402 : std_logic;
signal n16403 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_16_32_0_\ : std_logic;
signal n16404 : std_logic;
signal blink_counter_25 : std_logic;
signal \CLK_c\ : std_logic;
signal \c0.data_out_5__5__N_950\ : std_logic;
signal \c0.n17438\ : std_logic;
signal \c0.data_out_6__3__N_781\ : std_logic;
signal \c0.n17653\ : std_logic;
signal \c0.n17976\ : std_logic;
signal \c0.n8953\ : std_logic;
signal data_out_8_5 : std_logic;
signal \c0.data_out_6_6\ : std_logic;
signal \c0.n8922\ : std_logic;
signal data_out_8_4 : std_logic;
signal data_out_8_3 : std_logic;
signal \c0.n17620\ : std_logic;
signal \c0.n17611\ : std_logic;
signal \c0.n17659\ : std_logic;
signal \c0.n8777\ : std_logic;
signal \UART_TRANSMITTER_state_2\ : std_logic;
signal \c0.n17918\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50526\,
            DIN => \N__50525\,
            DOUT => \N__50524\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50526\,
            PADOUT => \N__50525\,
            PADIN => \N__50524\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30263\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50517\,
            DIN => \N__50516\,
            DOUT => \N__50515\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50517\,
            PADOUT => \N__50516\,
            PADIN => \N__50515\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50508\,
            DIN => \N__50507\,
            DOUT => \N__50506\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50508\,
            PADOUT => \N__50507\,
            PADIN => \N__50506\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__50364\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50499\,
            DIN => \N__50498\,
            DOUT => \N__50497\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50499\,
            PADOUT => \N__50498\,
            PADIN => \N__50497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21152\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21122\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50490\,
            DIN => \N__50489\,
            DOUT => \N__50488\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50490\,
            PADOUT => \N__50489\,
            PADIN => \N__50488\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37175\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__21161\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50481\,
            DIN => \N__50480\,
            DOUT => \N__50479\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50481\,
            PADOUT => \N__50480\,
            PADIN => \N__50479\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__12591\ : InMux
    port map (
            O => \N__50462\,
            I => n16404
        );

    \I__12590\ : InMux
    port map (
            O => \N__50459\,
            I => \N__50456\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__50456\,
            I => \N__50453\
        );

    \I__12588\ : Span4Mux_v
    port map (
            O => \N__50453\,
            I => \N__50450\
        );

    \I__12587\ : Span4Mux_h
    port map (
            O => \N__50450\,
            I => \N__50447\
        );

    \I__12586\ : Span4Mux_h
    port map (
            O => \N__50447\,
            I => \N__50443\
        );

    \I__12585\ : InMux
    port map (
            O => \N__50446\,
            I => \N__50440\
        );

    \I__12584\ : Odrv4
    port map (
            O => \N__50443\,
            I => blink_counter_25
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__50440\,
            I => blink_counter_25
        );

    \I__12582\ : ClkMux
    port map (
            O => \N__50435\,
            I => \N__49880\
        );

    \I__12581\ : ClkMux
    port map (
            O => \N__50434\,
            I => \N__49880\
        );

    \I__12580\ : ClkMux
    port map (
            O => \N__50433\,
            I => \N__49880\
        );

    \I__12579\ : ClkMux
    port map (
            O => \N__50432\,
            I => \N__49880\
        );

    \I__12578\ : ClkMux
    port map (
            O => \N__50431\,
            I => \N__49880\
        );

    \I__12577\ : ClkMux
    port map (
            O => \N__50430\,
            I => \N__49880\
        );

    \I__12576\ : ClkMux
    port map (
            O => \N__50429\,
            I => \N__49880\
        );

    \I__12575\ : ClkMux
    port map (
            O => \N__50428\,
            I => \N__49880\
        );

    \I__12574\ : ClkMux
    port map (
            O => \N__50427\,
            I => \N__49880\
        );

    \I__12573\ : ClkMux
    port map (
            O => \N__50426\,
            I => \N__49880\
        );

    \I__12572\ : ClkMux
    port map (
            O => \N__50425\,
            I => \N__49880\
        );

    \I__12571\ : ClkMux
    port map (
            O => \N__50424\,
            I => \N__49880\
        );

    \I__12570\ : ClkMux
    port map (
            O => \N__50423\,
            I => \N__49880\
        );

    \I__12569\ : ClkMux
    port map (
            O => \N__50422\,
            I => \N__49880\
        );

    \I__12568\ : ClkMux
    port map (
            O => \N__50421\,
            I => \N__49880\
        );

    \I__12567\ : ClkMux
    port map (
            O => \N__50420\,
            I => \N__49880\
        );

    \I__12566\ : ClkMux
    port map (
            O => \N__50419\,
            I => \N__49880\
        );

    \I__12565\ : ClkMux
    port map (
            O => \N__50418\,
            I => \N__49880\
        );

    \I__12564\ : ClkMux
    port map (
            O => \N__50417\,
            I => \N__49880\
        );

    \I__12563\ : ClkMux
    port map (
            O => \N__50416\,
            I => \N__49880\
        );

    \I__12562\ : ClkMux
    port map (
            O => \N__50415\,
            I => \N__49880\
        );

    \I__12561\ : ClkMux
    port map (
            O => \N__50414\,
            I => \N__49880\
        );

    \I__12560\ : ClkMux
    port map (
            O => \N__50413\,
            I => \N__49880\
        );

    \I__12559\ : ClkMux
    port map (
            O => \N__50412\,
            I => \N__49880\
        );

    \I__12558\ : ClkMux
    port map (
            O => \N__50411\,
            I => \N__49880\
        );

    \I__12557\ : ClkMux
    port map (
            O => \N__50410\,
            I => \N__49880\
        );

    \I__12556\ : ClkMux
    port map (
            O => \N__50409\,
            I => \N__49880\
        );

    \I__12555\ : ClkMux
    port map (
            O => \N__50408\,
            I => \N__49880\
        );

    \I__12554\ : ClkMux
    port map (
            O => \N__50407\,
            I => \N__49880\
        );

    \I__12553\ : ClkMux
    port map (
            O => \N__50406\,
            I => \N__49880\
        );

    \I__12552\ : ClkMux
    port map (
            O => \N__50405\,
            I => \N__49880\
        );

    \I__12551\ : ClkMux
    port map (
            O => \N__50404\,
            I => \N__49880\
        );

    \I__12550\ : ClkMux
    port map (
            O => \N__50403\,
            I => \N__49880\
        );

    \I__12549\ : ClkMux
    port map (
            O => \N__50402\,
            I => \N__49880\
        );

    \I__12548\ : ClkMux
    port map (
            O => \N__50401\,
            I => \N__49880\
        );

    \I__12547\ : ClkMux
    port map (
            O => \N__50400\,
            I => \N__49880\
        );

    \I__12546\ : ClkMux
    port map (
            O => \N__50399\,
            I => \N__49880\
        );

    \I__12545\ : ClkMux
    port map (
            O => \N__50398\,
            I => \N__49880\
        );

    \I__12544\ : ClkMux
    port map (
            O => \N__50397\,
            I => \N__49880\
        );

    \I__12543\ : ClkMux
    port map (
            O => \N__50396\,
            I => \N__49880\
        );

    \I__12542\ : ClkMux
    port map (
            O => \N__50395\,
            I => \N__49880\
        );

    \I__12541\ : ClkMux
    port map (
            O => \N__50394\,
            I => \N__49880\
        );

    \I__12540\ : ClkMux
    port map (
            O => \N__50393\,
            I => \N__49880\
        );

    \I__12539\ : ClkMux
    port map (
            O => \N__50392\,
            I => \N__49880\
        );

    \I__12538\ : ClkMux
    port map (
            O => \N__50391\,
            I => \N__49880\
        );

    \I__12537\ : ClkMux
    port map (
            O => \N__50390\,
            I => \N__49880\
        );

    \I__12536\ : ClkMux
    port map (
            O => \N__50389\,
            I => \N__49880\
        );

    \I__12535\ : ClkMux
    port map (
            O => \N__50388\,
            I => \N__49880\
        );

    \I__12534\ : ClkMux
    port map (
            O => \N__50387\,
            I => \N__49880\
        );

    \I__12533\ : ClkMux
    port map (
            O => \N__50386\,
            I => \N__49880\
        );

    \I__12532\ : ClkMux
    port map (
            O => \N__50385\,
            I => \N__49880\
        );

    \I__12531\ : ClkMux
    port map (
            O => \N__50384\,
            I => \N__49880\
        );

    \I__12530\ : ClkMux
    port map (
            O => \N__50383\,
            I => \N__49880\
        );

    \I__12529\ : ClkMux
    port map (
            O => \N__50382\,
            I => \N__49880\
        );

    \I__12528\ : ClkMux
    port map (
            O => \N__50381\,
            I => \N__49880\
        );

    \I__12527\ : ClkMux
    port map (
            O => \N__50380\,
            I => \N__49880\
        );

    \I__12526\ : ClkMux
    port map (
            O => \N__50379\,
            I => \N__49880\
        );

    \I__12525\ : ClkMux
    port map (
            O => \N__50378\,
            I => \N__49880\
        );

    \I__12524\ : ClkMux
    port map (
            O => \N__50377\,
            I => \N__49880\
        );

    \I__12523\ : ClkMux
    port map (
            O => \N__50376\,
            I => \N__49880\
        );

    \I__12522\ : ClkMux
    port map (
            O => \N__50375\,
            I => \N__49880\
        );

    \I__12521\ : ClkMux
    port map (
            O => \N__50374\,
            I => \N__49880\
        );

    \I__12520\ : ClkMux
    port map (
            O => \N__50373\,
            I => \N__49880\
        );

    \I__12519\ : ClkMux
    port map (
            O => \N__50372\,
            I => \N__49880\
        );

    \I__12518\ : ClkMux
    port map (
            O => \N__50371\,
            I => \N__49880\
        );

    \I__12517\ : ClkMux
    port map (
            O => \N__50370\,
            I => \N__49880\
        );

    \I__12516\ : ClkMux
    port map (
            O => \N__50369\,
            I => \N__49880\
        );

    \I__12515\ : ClkMux
    port map (
            O => \N__50368\,
            I => \N__49880\
        );

    \I__12514\ : ClkMux
    port map (
            O => \N__50367\,
            I => \N__49880\
        );

    \I__12513\ : ClkMux
    port map (
            O => \N__50366\,
            I => \N__49880\
        );

    \I__12512\ : ClkMux
    port map (
            O => \N__50365\,
            I => \N__49880\
        );

    \I__12511\ : ClkMux
    port map (
            O => \N__50364\,
            I => \N__49880\
        );

    \I__12510\ : ClkMux
    port map (
            O => \N__50363\,
            I => \N__49880\
        );

    \I__12509\ : ClkMux
    port map (
            O => \N__50362\,
            I => \N__49880\
        );

    \I__12508\ : ClkMux
    port map (
            O => \N__50361\,
            I => \N__49880\
        );

    \I__12507\ : ClkMux
    port map (
            O => \N__50360\,
            I => \N__49880\
        );

    \I__12506\ : ClkMux
    port map (
            O => \N__50359\,
            I => \N__49880\
        );

    \I__12505\ : ClkMux
    port map (
            O => \N__50358\,
            I => \N__49880\
        );

    \I__12504\ : ClkMux
    port map (
            O => \N__50357\,
            I => \N__49880\
        );

    \I__12503\ : ClkMux
    port map (
            O => \N__50356\,
            I => \N__49880\
        );

    \I__12502\ : ClkMux
    port map (
            O => \N__50355\,
            I => \N__49880\
        );

    \I__12501\ : ClkMux
    port map (
            O => \N__50354\,
            I => \N__49880\
        );

    \I__12500\ : ClkMux
    port map (
            O => \N__50353\,
            I => \N__49880\
        );

    \I__12499\ : ClkMux
    port map (
            O => \N__50352\,
            I => \N__49880\
        );

    \I__12498\ : ClkMux
    port map (
            O => \N__50351\,
            I => \N__49880\
        );

    \I__12497\ : ClkMux
    port map (
            O => \N__50350\,
            I => \N__49880\
        );

    \I__12496\ : ClkMux
    port map (
            O => \N__50349\,
            I => \N__49880\
        );

    \I__12495\ : ClkMux
    port map (
            O => \N__50348\,
            I => \N__49880\
        );

    \I__12494\ : ClkMux
    port map (
            O => \N__50347\,
            I => \N__49880\
        );

    \I__12493\ : ClkMux
    port map (
            O => \N__50346\,
            I => \N__49880\
        );

    \I__12492\ : ClkMux
    port map (
            O => \N__50345\,
            I => \N__49880\
        );

    \I__12491\ : ClkMux
    port map (
            O => \N__50344\,
            I => \N__49880\
        );

    \I__12490\ : ClkMux
    port map (
            O => \N__50343\,
            I => \N__49880\
        );

    \I__12489\ : ClkMux
    port map (
            O => \N__50342\,
            I => \N__49880\
        );

    \I__12488\ : ClkMux
    port map (
            O => \N__50341\,
            I => \N__49880\
        );

    \I__12487\ : ClkMux
    port map (
            O => \N__50340\,
            I => \N__49880\
        );

    \I__12486\ : ClkMux
    port map (
            O => \N__50339\,
            I => \N__49880\
        );

    \I__12485\ : ClkMux
    port map (
            O => \N__50338\,
            I => \N__49880\
        );

    \I__12484\ : ClkMux
    port map (
            O => \N__50337\,
            I => \N__49880\
        );

    \I__12483\ : ClkMux
    port map (
            O => \N__50336\,
            I => \N__49880\
        );

    \I__12482\ : ClkMux
    port map (
            O => \N__50335\,
            I => \N__49880\
        );

    \I__12481\ : ClkMux
    port map (
            O => \N__50334\,
            I => \N__49880\
        );

    \I__12480\ : ClkMux
    port map (
            O => \N__50333\,
            I => \N__49880\
        );

    \I__12479\ : ClkMux
    port map (
            O => \N__50332\,
            I => \N__49880\
        );

    \I__12478\ : ClkMux
    port map (
            O => \N__50331\,
            I => \N__49880\
        );

    \I__12477\ : ClkMux
    port map (
            O => \N__50330\,
            I => \N__49880\
        );

    \I__12476\ : ClkMux
    port map (
            O => \N__50329\,
            I => \N__49880\
        );

    \I__12475\ : ClkMux
    port map (
            O => \N__50328\,
            I => \N__49880\
        );

    \I__12474\ : ClkMux
    port map (
            O => \N__50327\,
            I => \N__49880\
        );

    \I__12473\ : ClkMux
    port map (
            O => \N__50326\,
            I => \N__49880\
        );

    \I__12472\ : ClkMux
    port map (
            O => \N__50325\,
            I => \N__49880\
        );

    \I__12471\ : ClkMux
    port map (
            O => \N__50324\,
            I => \N__49880\
        );

    \I__12470\ : ClkMux
    port map (
            O => \N__50323\,
            I => \N__49880\
        );

    \I__12469\ : ClkMux
    port map (
            O => \N__50322\,
            I => \N__49880\
        );

    \I__12468\ : ClkMux
    port map (
            O => \N__50321\,
            I => \N__49880\
        );

    \I__12467\ : ClkMux
    port map (
            O => \N__50320\,
            I => \N__49880\
        );

    \I__12466\ : ClkMux
    port map (
            O => \N__50319\,
            I => \N__49880\
        );

    \I__12465\ : ClkMux
    port map (
            O => \N__50318\,
            I => \N__49880\
        );

    \I__12464\ : ClkMux
    port map (
            O => \N__50317\,
            I => \N__49880\
        );

    \I__12463\ : ClkMux
    port map (
            O => \N__50316\,
            I => \N__49880\
        );

    \I__12462\ : ClkMux
    port map (
            O => \N__50315\,
            I => \N__49880\
        );

    \I__12461\ : ClkMux
    port map (
            O => \N__50314\,
            I => \N__49880\
        );

    \I__12460\ : ClkMux
    port map (
            O => \N__50313\,
            I => \N__49880\
        );

    \I__12459\ : ClkMux
    port map (
            O => \N__50312\,
            I => \N__49880\
        );

    \I__12458\ : ClkMux
    port map (
            O => \N__50311\,
            I => \N__49880\
        );

    \I__12457\ : ClkMux
    port map (
            O => \N__50310\,
            I => \N__49880\
        );

    \I__12456\ : ClkMux
    port map (
            O => \N__50309\,
            I => \N__49880\
        );

    \I__12455\ : ClkMux
    port map (
            O => \N__50308\,
            I => \N__49880\
        );

    \I__12454\ : ClkMux
    port map (
            O => \N__50307\,
            I => \N__49880\
        );

    \I__12453\ : ClkMux
    port map (
            O => \N__50306\,
            I => \N__49880\
        );

    \I__12452\ : ClkMux
    port map (
            O => \N__50305\,
            I => \N__49880\
        );

    \I__12451\ : ClkMux
    port map (
            O => \N__50304\,
            I => \N__49880\
        );

    \I__12450\ : ClkMux
    port map (
            O => \N__50303\,
            I => \N__49880\
        );

    \I__12449\ : ClkMux
    port map (
            O => \N__50302\,
            I => \N__49880\
        );

    \I__12448\ : ClkMux
    port map (
            O => \N__50301\,
            I => \N__49880\
        );

    \I__12447\ : ClkMux
    port map (
            O => \N__50300\,
            I => \N__49880\
        );

    \I__12446\ : ClkMux
    port map (
            O => \N__50299\,
            I => \N__49880\
        );

    \I__12445\ : ClkMux
    port map (
            O => \N__50298\,
            I => \N__49880\
        );

    \I__12444\ : ClkMux
    port map (
            O => \N__50297\,
            I => \N__49880\
        );

    \I__12443\ : ClkMux
    port map (
            O => \N__50296\,
            I => \N__49880\
        );

    \I__12442\ : ClkMux
    port map (
            O => \N__50295\,
            I => \N__49880\
        );

    \I__12441\ : ClkMux
    port map (
            O => \N__50294\,
            I => \N__49880\
        );

    \I__12440\ : ClkMux
    port map (
            O => \N__50293\,
            I => \N__49880\
        );

    \I__12439\ : ClkMux
    port map (
            O => \N__50292\,
            I => \N__49880\
        );

    \I__12438\ : ClkMux
    port map (
            O => \N__50291\,
            I => \N__49880\
        );

    \I__12437\ : ClkMux
    port map (
            O => \N__50290\,
            I => \N__49880\
        );

    \I__12436\ : ClkMux
    port map (
            O => \N__50289\,
            I => \N__49880\
        );

    \I__12435\ : ClkMux
    port map (
            O => \N__50288\,
            I => \N__49880\
        );

    \I__12434\ : ClkMux
    port map (
            O => \N__50287\,
            I => \N__49880\
        );

    \I__12433\ : ClkMux
    port map (
            O => \N__50286\,
            I => \N__49880\
        );

    \I__12432\ : ClkMux
    port map (
            O => \N__50285\,
            I => \N__49880\
        );

    \I__12431\ : ClkMux
    port map (
            O => \N__50284\,
            I => \N__49880\
        );

    \I__12430\ : ClkMux
    port map (
            O => \N__50283\,
            I => \N__49880\
        );

    \I__12429\ : ClkMux
    port map (
            O => \N__50282\,
            I => \N__49880\
        );

    \I__12428\ : ClkMux
    port map (
            O => \N__50281\,
            I => \N__49880\
        );

    \I__12427\ : ClkMux
    port map (
            O => \N__50280\,
            I => \N__49880\
        );

    \I__12426\ : ClkMux
    port map (
            O => \N__50279\,
            I => \N__49880\
        );

    \I__12425\ : ClkMux
    port map (
            O => \N__50278\,
            I => \N__49880\
        );

    \I__12424\ : ClkMux
    port map (
            O => \N__50277\,
            I => \N__49880\
        );

    \I__12423\ : ClkMux
    port map (
            O => \N__50276\,
            I => \N__49880\
        );

    \I__12422\ : ClkMux
    port map (
            O => \N__50275\,
            I => \N__49880\
        );

    \I__12421\ : ClkMux
    port map (
            O => \N__50274\,
            I => \N__49880\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__50273\,
            I => \N__49880\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__50272\,
            I => \N__49880\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__50271\,
            I => \N__49880\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__50270\,
            I => \N__49880\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__50269\,
            I => \N__49880\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__50268\,
            I => \N__49880\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__50267\,
            I => \N__49880\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__50266\,
            I => \N__49880\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__50265\,
            I => \N__49880\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__50264\,
            I => \N__49880\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__50263\,
            I => \N__49880\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__50262\,
            I => \N__49880\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__50261\,
            I => \N__49880\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__50260\,
            I => \N__49880\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__50259\,
            I => \N__49880\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__50258\,
            I => \N__49880\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__50257\,
            I => \N__49880\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__50256\,
            I => \N__49880\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__50255\,
            I => \N__49880\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__50254\,
            I => \N__49880\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__50253\,
            I => \N__49880\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__50252\,
            I => \N__49880\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__50251\,
            I => \N__49880\
        );

    \I__12397\ : GlobalMux
    port map (
            O => \N__49880\,
            I => \N__49877\
        );

    \I__12396\ : gio2CtrlBuf
    port map (
            O => \N__49877\,
            I => \CLK_c\
        );

    \I__12395\ : InMux
    port map (
            O => \N__49874\,
            I => \N__49869\
        );

    \I__12394\ : InMux
    port map (
            O => \N__49873\,
            I => \N__49863\
        );

    \I__12393\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49860\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__49869\,
            I => \N__49857\
        );

    \I__12391\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49854\
        );

    \I__12390\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49850\
        );

    \I__12389\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49847\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__49863\,
            I => \N__49843\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__49860\,
            I => \N__49836\
        );

    \I__12386\ : Span4Mux_h
    port map (
            O => \N__49857\,
            I => \N__49836\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__49854\,
            I => \N__49836\
        );

    \I__12384\ : InMux
    port map (
            O => \N__49853\,
            I => \N__49833\
        );

    \I__12383\ : LocalMux
    port map (
            O => \N__49850\,
            I => \N__49830\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__49847\,
            I => \N__49827\
        );

    \I__12381\ : InMux
    port map (
            O => \N__49846\,
            I => \N__49824\
        );

    \I__12380\ : Span4Mux_h
    port map (
            O => \N__49843\,
            I => \N__49819\
        );

    \I__12379\ : Span4Mux_v
    port map (
            O => \N__49836\,
            I => \N__49819\
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__49833\,
            I => \c0.data_out_5__5__N_950\
        );

    \I__12377\ : Odrv4
    port map (
            O => \N__49830\,
            I => \c0.data_out_5__5__N_950\
        );

    \I__12376\ : Odrv4
    port map (
            O => \N__49827\,
            I => \c0.data_out_5__5__N_950\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__49824\,
            I => \c0.data_out_5__5__N_950\
        );

    \I__12374\ : Odrv4
    port map (
            O => \N__49819\,
            I => \c0.data_out_5__5__N_950\
        );

    \I__12373\ : InMux
    port map (
            O => \N__49808\,
            I => \N__49804\
        );

    \I__12372\ : InMux
    port map (
            O => \N__49807\,
            I => \N__49801\
        );

    \I__12371\ : LocalMux
    port map (
            O => \N__49804\,
            I => \N__49798\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__49801\,
            I => \c0.n17438\
        );

    \I__12369\ : Odrv4
    port map (
            O => \N__49798\,
            I => \c0.n17438\
        );

    \I__12368\ : CascadeMux
    port map (
            O => \N__49793\,
            I => \N__49787\
        );

    \I__12367\ : InMux
    port map (
            O => \N__49792\,
            I => \N__49784\
        );

    \I__12366\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49780\
        );

    \I__12365\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49777\
        );

    \I__12364\ : InMux
    port map (
            O => \N__49787\,
            I => \N__49774\
        );

    \I__12363\ : LocalMux
    port map (
            O => \N__49784\,
            I => \N__49771\
        );

    \I__12362\ : InMux
    port map (
            O => \N__49783\,
            I => \N__49768\
        );

    \I__12361\ : LocalMux
    port map (
            O => \N__49780\,
            I => \N__49763\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__49777\,
            I => \N__49763\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__49774\,
            I => \N__49760\
        );

    \I__12358\ : Span4Mux_h
    port map (
            O => \N__49771\,
            I => \N__49755\
        );

    \I__12357\ : LocalMux
    port map (
            O => \N__49768\,
            I => \N__49755\
        );

    \I__12356\ : Odrv12
    port map (
            O => \N__49763\,
            I => \c0.data_out_6__3__N_781\
        );

    \I__12355\ : Odrv4
    port map (
            O => \N__49760\,
            I => \c0.data_out_6__3__N_781\
        );

    \I__12354\ : Odrv4
    port map (
            O => \N__49755\,
            I => \c0.data_out_6__3__N_781\
        );

    \I__12353\ : InMux
    port map (
            O => \N__49748\,
            I => \N__49745\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__49745\,
            I => \N__49741\
        );

    \I__12351\ : InMux
    port map (
            O => \N__49744\,
            I => \N__49738\
        );

    \I__12350\ : Span4Mux_h
    port map (
            O => \N__49741\,
            I => \N__49733\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__49738\,
            I => \N__49733\
        );

    \I__12348\ : Odrv4
    port map (
            O => \N__49733\,
            I => \c0.n17653\
        );

    \I__12347\ : InMux
    port map (
            O => \N__49730\,
            I => \N__49727\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__49727\,
            I => \N__49724\
        );

    \I__12345\ : Odrv4
    port map (
            O => \N__49724\,
            I => \c0.n17976\
        );

    \I__12344\ : InMux
    port map (
            O => \N__49721\,
            I => \N__49718\
        );

    \I__12343\ : LocalMux
    port map (
            O => \N__49718\,
            I => \N__49715\
        );

    \I__12342\ : Span4Mux_h
    port map (
            O => \N__49715\,
            I => \N__49712\
        );

    \I__12341\ : Odrv4
    port map (
            O => \N__49712\,
            I => \c0.n8953\
        );

    \I__12340\ : CascadeMux
    port map (
            O => \N__49709\,
            I => \N__49703\
        );

    \I__12339\ : InMux
    port map (
            O => \N__49708\,
            I => \N__49698\
        );

    \I__12338\ : InMux
    port map (
            O => \N__49707\,
            I => \N__49698\
        );

    \I__12337\ : InMux
    port map (
            O => \N__49706\,
            I => \N__49694\
        );

    \I__12336\ : InMux
    port map (
            O => \N__49703\,
            I => \N__49691\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__49698\,
            I => \N__49688\
        );

    \I__12334\ : InMux
    port map (
            O => \N__49697\,
            I => \N__49685\
        );

    \I__12333\ : LocalMux
    port map (
            O => \N__49694\,
            I => \N__49682\
        );

    \I__12332\ : LocalMux
    port map (
            O => \N__49691\,
            I => \N__49679\
        );

    \I__12331\ : Span4Mux_s3_v
    port map (
            O => \N__49688\,
            I => \N__49676\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__49685\,
            I => data_out_8_5
        );

    \I__12329\ : Odrv4
    port map (
            O => \N__49682\,
            I => data_out_8_5
        );

    \I__12328\ : Odrv12
    port map (
            O => \N__49679\,
            I => data_out_8_5
        );

    \I__12327\ : Odrv4
    port map (
            O => \N__49676\,
            I => data_out_8_5
        );

    \I__12326\ : InMux
    port map (
            O => \N__49667\,
            I => \N__49664\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__49664\,
            I => \N__49660\
        );

    \I__12324\ : InMux
    port map (
            O => \N__49663\,
            I => \N__49657\
        );

    \I__12323\ : Span4Mux_v
    port map (
            O => \N__49660\,
            I => \N__49652\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__49657\,
            I => \N__49652\
        );

    \I__12321\ : Span4Mux_h
    port map (
            O => \N__49652\,
            I => \N__49648\
        );

    \I__12320\ : InMux
    port map (
            O => \N__49651\,
            I => \N__49645\
        );

    \I__12319\ : Span4Mux_v
    port map (
            O => \N__49648\,
            I => \N__49642\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__49645\,
            I => \c0.data_out_6_6\
        );

    \I__12317\ : Odrv4
    port map (
            O => \N__49642\,
            I => \c0.data_out_6_6\
        );

    \I__12316\ : InMux
    port map (
            O => \N__49637\,
            I => \N__49634\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__49634\,
            I => \N__49630\
        );

    \I__12314\ : InMux
    port map (
            O => \N__49633\,
            I => \N__49627\
        );

    \I__12313\ : Span12Mux_h
    port map (
            O => \N__49630\,
            I => \N__49624\
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__49627\,
            I => \N__49621\
        );

    \I__12311\ : Odrv12
    port map (
            O => \N__49624\,
            I => \c0.n8922\
        );

    \I__12310\ : Odrv4
    port map (
            O => \N__49621\,
            I => \c0.n8922\
        );

    \I__12309\ : InMux
    port map (
            O => \N__49616\,
            I => \N__49612\
        );

    \I__12308\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49607\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__49612\,
            I => \N__49604\
        );

    \I__12306\ : InMux
    port map (
            O => \N__49611\,
            I => \N__49598\
        );

    \I__12305\ : InMux
    port map (
            O => \N__49610\,
            I => \N__49598\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__49607\,
            I => \N__49595\
        );

    \I__12303\ : Span4Mux_h
    port map (
            O => \N__49604\,
            I => \N__49592\
        );

    \I__12302\ : InMux
    port map (
            O => \N__49603\,
            I => \N__49589\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__49598\,
            I => \N__49586\
        );

    \I__12300\ : Span4Mux_h
    port map (
            O => \N__49595\,
            I => \N__49581\
        );

    \I__12299\ : Span4Mux_h
    port map (
            O => \N__49592\,
            I => \N__49581\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__49589\,
            I => data_out_8_4
        );

    \I__12297\ : Odrv12
    port map (
            O => \N__49586\,
            I => data_out_8_4
        );

    \I__12296\ : Odrv4
    port map (
            O => \N__49581\,
            I => data_out_8_4
        );

    \I__12295\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49571\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__49571\,
            I => \N__49568\
        );

    \I__12293\ : Span4Mux_h
    port map (
            O => \N__49568\,
            I => \N__49562\
        );

    \I__12292\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49555\
        );

    \I__12291\ : InMux
    port map (
            O => \N__49566\,
            I => \N__49555\
        );

    \I__12290\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49555\
        );

    \I__12289\ : Odrv4
    port map (
            O => \N__49562\,
            I => data_out_8_3
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__49555\,
            I => data_out_8_3
        );

    \I__12287\ : InMux
    port map (
            O => \N__49550\,
            I => \N__49546\
        );

    \I__12286\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49543\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49540\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__49543\,
            I => \N__49537\
        );

    \I__12283\ : Span4Mux_s3_v
    port map (
            O => \N__49540\,
            I => \N__49534\
        );

    \I__12282\ : Span4Mux_h
    port map (
            O => \N__49537\,
            I => \N__49531\
        );

    \I__12281\ : Odrv4
    port map (
            O => \N__49534\,
            I => \c0.n17620\
        );

    \I__12280\ : Odrv4
    port map (
            O => \N__49531\,
            I => \c0.n17620\
        );

    \I__12279\ : InMux
    port map (
            O => \N__49526\,
            I => \N__49523\
        );

    \I__12278\ : LocalMux
    port map (
            O => \N__49523\,
            I => \N__49520\
        );

    \I__12277\ : Span4Mux_h
    port map (
            O => \N__49520\,
            I => \N__49516\
        );

    \I__12276\ : InMux
    port map (
            O => \N__49519\,
            I => \N__49513\
        );

    \I__12275\ : Span4Mux_h
    port map (
            O => \N__49516\,
            I => \N__49510\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__49513\,
            I => \c0.n17611\
        );

    \I__12273\ : Odrv4
    port map (
            O => \N__49510\,
            I => \c0.n17611\
        );

    \I__12272\ : InMux
    port map (
            O => \N__49505\,
            I => \N__49501\
        );

    \I__12271\ : InMux
    port map (
            O => \N__49504\,
            I => \N__49498\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__49501\,
            I => \N__49493\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__49498\,
            I => \N__49493\
        );

    \I__12268\ : Span4Mux_h
    port map (
            O => \N__49493\,
            I => \N__49490\
        );

    \I__12267\ : Odrv4
    port map (
            O => \N__49490\,
            I => \c0.n17659\
        );

    \I__12266\ : CascadeMux
    port map (
            O => \N__49487\,
            I => \N__49483\
        );

    \I__12265\ : CascadeMux
    port map (
            O => \N__49486\,
            I => \N__49480\
        );

    \I__12264\ : InMux
    port map (
            O => \N__49483\,
            I => \N__49477\
        );

    \I__12263\ : InMux
    port map (
            O => \N__49480\,
            I => \N__49473\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49470\
        );

    \I__12261\ : InMux
    port map (
            O => \N__49476\,
            I => \N__49467\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49464\
        );

    \I__12259\ : Span4Mux_h
    port map (
            O => \N__49470\,
            I => \N__49461\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__49467\,
            I => \N__49456\
        );

    \I__12257\ : Span4Mux_h
    port map (
            O => \N__49464\,
            I => \N__49456\
        );

    \I__12256\ : Odrv4
    port map (
            O => \N__49461\,
            I => \c0.n8777\
        );

    \I__12255\ : Odrv4
    port map (
            O => \N__49456\,
            I => \c0.n8777\
        );

    \I__12254\ : InMux
    port map (
            O => \N__49451\,
            I => \N__49437\
        );

    \I__12253\ : InMux
    port map (
            O => \N__49450\,
            I => \N__49437\
        );

    \I__12252\ : CascadeMux
    port map (
            O => \N__49449\,
            I => \N__49432\
        );

    \I__12251\ : InMux
    port map (
            O => \N__49448\,
            I => \N__49427\
        );

    \I__12250\ : InMux
    port map (
            O => \N__49447\,
            I => \N__49427\
        );

    \I__12249\ : InMux
    port map (
            O => \N__49446\,
            I => \N__49424\
        );

    \I__12248\ : CascadeMux
    port map (
            O => \N__49445\,
            I => \N__49411\
        );

    \I__12247\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49404\
        );

    \I__12246\ : InMux
    port map (
            O => \N__49443\,
            I => \N__49404\
        );

    \I__12245\ : InMux
    port map (
            O => \N__49442\,
            I => \N__49404\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__49437\,
            I => \N__49401\
        );

    \I__12243\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49398\
        );

    \I__12242\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49392\
        );

    \I__12241\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49392\
        );

    \I__12240\ : LocalMux
    port map (
            O => \N__49427\,
            I => \N__49389\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__49424\,
            I => \N__49386\
        );

    \I__12238\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49378\
        );

    \I__12237\ : InMux
    port map (
            O => \N__49422\,
            I => \N__49378\
        );

    \I__12236\ : InMux
    port map (
            O => \N__49421\,
            I => \N__49371\
        );

    \I__12235\ : InMux
    port map (
            O => \N__49420\,
            I => \N__49371\
        );

    \I__12234\ : InMux
    port map (
            O => \N__49419\,
            I => \N__49371\
        );

    \I__12233\ : InMux
    port map (
            O => \N__49418\,
            I => \N__49368\
        );

    \I__12232\ : InMux
    port map (
            O => \N__49417\,
            I => \N__49365\
        );

    \I__12231\ : InMux
    port map (
            O => \N__49416\,
            I => \N__49356\
        );

    \I__12230\ : InMux
    port map (
            O => \N__49415\,
            I => \N__49356\
        );

    \I__12229\ : InMux
    port map (
            O => \N__49414\,
            I => \N__49356\
        );

    \I__12228\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49353\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__49404\,
            I => \N__49350\
        );

    \I__12226\ : Span4Mux_s3_v
    port map (
            O => \N__49401\,
            I => \N__49347\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__49398\,
            I => \N__49344\
        );

    \I__12224\ : InMux
    port map (
            O => \N__49397\,
            I => \N__49341\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__49392\,
            I => \N__49334\
        );

    \I__12222\ : Span4Mux_s3_v
    port map (
            O => \N__49389\,
            I => \N__49334\
        );

    \I__12221\ : Span4Mux_s3_v
    port map (
            O => \N__49386\,
            I => \N__49334\
        );

    \I__12220\ : InMux
    port map (
            O => \N__49385\,
            I => \N__49329\
        );

    \I__12219\ : InMux
    port map (
            O => \N__49384\,
            I => \N__49329\
        );

    \I__12218\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49318\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__49378\,
            I => \N__49309\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__49371\,
            I => \N__49309\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__49368\,
            I => \N__49309\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__49365\,
            I => \N__49309\
        );

    \I__12213\ : CascadeMux
    port map (
            O => \N__49364\,
            I => \N__49305\
        );

    \I__12212\ : CascadeMux
    port map (
            O => \N__49363\,
            I => \N__49301\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__49356\,
            I => \N__49298\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__49353\,
            I => \N__49295\
        );

    \I__12209\ : Span4Mux_s3_v
    port map (
            O => \N__49350\,
            I => \N__49292\
        );

    \I__12208\ : Span4Mux_h
    port map (
            O => \N__49347\,
            I => \N__49282\
        );

    \I__12207\ : Span4Mux_h
    port map (
            O => \N__49344\,
            I => \N__49282\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__49341\,
            I => \N__49282\
        );

    \I__12205\ : Span4Mux_h
    port map (
            O => \N__49334\,
            I => \N__49277\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__49329\,
            I => \N__49277\
        );

    \I__12203\ : InMux
    port map (
            O => \N__49328\,
            I => \N__49272\
        );

    \I__12202\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49272\
        );

    \I__12201\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49267\
        );

    \I__12200\ : InMux
    port map (
            O => \N__49325\,
            I => \N__49267\
        );

    \I__12199\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49264\
        );

    \I__12198\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49257\
        );

    \I__12197\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49257\
        );

    \I__12196\ : InMux
    port map (
            O => \N__49321\,
            I => \N__49257\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__49318\,
            I => \N__49248\
        );

    \I__12194\ : Span4Mux_s3_v
    port map (
            O => \N__49309\,
            I => \N__49248\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__49308\,
            I => \N__49245\
        );

    \I__12192\ : InMux
    port map (
            O => \N__49305\,
            I => \N__49237\
        );

    \I__12191\ : InMux
    port map (
            O => \N__49304\,
            I => \N__49237\
        );

    \I__12190\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49237\
        );

    \I__12189\ : Span4Mux_s3_v
    port map (
            O => \N__49298\,
            I => \N__49230\
        );

    \I__12188\ : Span4Mux_s3_v
    port map (
            O => \N__49295\,
            I => \N__49230\
        );

    \I__12187\ : Span4Mux_h
    port map (
            O => \N__49292\,
            I => \N__49230\
        );

    \I__12186\ : InMux
    port map (
            O => \N__49291\,
            I => \N__49223\
        );

    \I__12185\ : InMux
    port map (
            O => \N__49290\,
            I => \N__49223\
        );

    \I__12184\ : InMux
    port map (
            O => \N__49289\,
            I => \N__49223\
        );

    \I__12183\ : Sp12to4
    port map (
            O => \N__49282\,
            I => \N__49218\
        );

    \I__12182\ : Sp12to4
    port map (
            O => \N__49277\,
            I => \N__49218\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__49272\,
            I => \N__49209\
        );

    \I__12180\ : LocalMux
    port map (
            O => \N__49267\,
            I => \N__49209\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__49264\,
            I => \N__49209\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__49257\,
            I => \N__49209\
        );

    \I__12177\ : InMux
    port map (
            O => \N__49256\,
            I => \N__49204\
        );

    \I__12176\ : InMux
    port map (
            O => \N__49255\,
            I => \N__49204\
        );

    \I__12175\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49199\
        );

    \I__12174\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49199\
        );

    \I__12173\ : Span4Mux_v
    port map (
            O => \N__49248\,
            I => \N__49196\
        );

    \I__12172\ : InMux
    port map (
            O => \N__49245\,
            I => \N__49191\
        );

    \I__12171\ : InMux
    port map (
            O => \N__49244\,
            I => \N__49191\
        );

    \I__12170\ : LocalMux
    port map (
            O => \N__49237\,
            I => \N__49184\
        );

    \I__12169\ : Span4Mux_v
    port map (
            O => \N__49230\,
            I => \N__49184\
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__49223\,
            I => \N__49184\
        );

    \I__12167\ : Span12Mux_s10_v
    port map (
            O => \N__49218\,
            I => \N__49181\
        );

    \I__12166\ : Span12Mux_s5_v
    port map (
            O => \N__49209\,
            I => \N__49176\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__49204\,
            I => \N__49176\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__49199\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12163\ : Odrv4
    port map (
            O => \N__49196\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__49191\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12161\ : Odrv4
    port map (
            O => \N__49184\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12160\ : Odrv12
    port map (
            O => \N__49181\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12159\ : Odrv12
    port map (
            O => \N__49176\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__12158\ : InMux
    port map (
            O => \N__49163\,
            I => \N__49160\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__49160\,
            I => \N__49157\
        );

    \I__12156\ : Span4Mux_h
    port map (
            O => \N__49157\,
            I => \N__49154\
        );

    \I__12155\ : Odrv4
    port map (
            O => \N__49154\,
            I => \c0.n17918\
        );

    \I__12154\ : InMux
    port map (
            O => \N__49151\,
            I => \bfn_16_31_0_\
        );

    \I__12153\ : InMux
    port map (
            O => \N__49148\,
            I => \N__49145\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__49145\,
            I => n9
        );

    \I__12151\ : InMux
    port map (
            O => \N__49142\,
            I => n16396
        );

    \I__12150\ : InMux
    port map (
            O => \N__49139\,
            I => \N__49136\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__49136\,
            I => n8_adj_2617
        );

    \I__12148\ : InMux
    port map (
            O => \N__49133\,
            I => n16397
        );

    \I__12147\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49127\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__49127\,
            I => n7
        );

    \I__12145\ : InMux
    port map (
            O => \N__49124\,
            I => n16398
        );

    \I__12144\ : InMux
    port map (
            O => \N__49121\,
            I => \N__49118\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__49118\,
            I => n6
        );

    \I__12142\ : InMux
    port map (
            O => \N__49115\,
            I => n16399
        );

    \I__12141\ : CascadeMux
    port map (
            O => \N__49112\,
            I => \N__49108\
        );

    \I__12140\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49103\
        );

    \I__12139\ : InMux
    port map (
            O => \N__49108\,
            I => \N__49103\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__49103\,
            I => \N__49099\
        );

    \I__12137\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49096\
        );

    \I__12136\ : Odrv12
    port map (
            O => \N__49099\,
            I => blink_counter_21
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__49096\,
            I => blink_counter_21
        );

    \I__12134\ : InMux
    port map (
            O => \N__49091\,
            I => n16400
        );

    \I__12133\ : InMux
    port map (
            O => \N__49088\,
            I => \N__49082\
        );

    \I__12132\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49082\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__49082\,
            I => \N__49079\
        );

    \I__12130\ : Span12Mux_h
    port map (
            O => \N__49079\,
            I => \N__49075\
        );

    \I__12129\ : InMux
    port map (
            O => \N__49078\,
            I => \N__49072\
        );

    \I__12128\ : Odrv12
    port map (
            O => \N__49075\,
            I => blink_counter_22
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__49072\,
            I => blink_counter_22
        );

    \I__12126\ : InMux
    port map (
            O => \N__49067\,
            I => n16401
        );

    \I__12125\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49058\
        );

    \I__12124\ : InMux
    port map (
            O => \N__49063\,
            I => \N__49058\
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__49058\,
            I => \N__49054\
        );

    \I__12122\ : InMux
    port map (
            O => \N__49057\,
            I => \N__49051\
        );

    \I__12121\ : Odrv12
    port map (
            O => \N__49054\,
            I => blink_counter_23
        );

    \I__12120\ : LocalMux
    port map (
            O => \N__49051\,
            I => blink_counter_23
        );

    \I__12119\ : InMux
    port map (
            O => \N__49046\,
            I => n16402
        );

    \I__12118\ : CascadeMux
    port map (
            O => \N__49043\,
            I => \N__49040\
        );

    \I__12117\ : InMux
    port map (
            O => \N__49040\,
            I => \N__49034\
        );

    \I__12116\ : InMux
    port map (
            O => \N__49039\,
            I => \N__49034\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__49034\,
            I => \N__49031\
        );

    \I__12114\ : Span4Mux_v
    port map (
            O => \N__49031\,
            I => \N__49028\
        );

    \I__12113\ : Span4Mux_h
    port map (
            O => \N__49028\,
            I => \N__49025\
        );

    \I__12112\ : Span4Mux_h
    port map (
            O => \N__49025\,
            I => \N__49021\
        );

    \I__12111\ : InMux
    port map (
            O => \N__49024\,
            I => \N__49018\
        );

    \I__12110\ : Odrv4
    port map (
            O => \N__49021\,
            I => blink_counter_24
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__49018\,
            I => blink_counter_24
        );

    \I__12108\ : InMux
    port map (
            O => \N__49013\,
            I => \bfn_16_32_0_\
        );

    \I__12107\ : InMux
    port map (
            O => \N__49010\,
            I => \N__49007\
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__49007\,
            I => n18
        );

    \I__12105\ : InMux
    port map (
            O => \N__49004\,
            I => \bfn_16_30_0_\
        );

    \I__12104\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48998\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__48998\,
            I => n17
        );

    \I__12102\ : InMux
    port map (
            O => \N__48995\,
            I => n16388
        );

    \I__12101\ : InMux
    port map (
            O => \N__48992\,
            I => \N__48989\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__48989\,
            I => n16
        );

    \I__12099\ : InMux
    port map (
            O => \N__48986\,
            I => n16389
        );

    \I__12098\ : InMux
    port map (
            O => \N__48983\,
            I => \N__48980\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__48980\,
            I => n15
        );

    \I__12096\ : InMux
    port map (
            O => \N__48977\,
            I => n16390
        );

    \I__12095\ : InMux
    port map (
            O => \N__48974\,
            I => \N__48971\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__48971\,
            I => n14
        );

    \I__12093\ : InMux
    port map (
            O => \N__48968\,
            I => n16391
        );

    \I__12092\ : InMux
    port map (
            O => \N__48965\,
            I => \N__48962\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__48962\,
            I => n13
        );

    \I__12090\ : InMux
    port map (
            O => \N__48959\,
            I => n16392
        );

    \I__12089\ : InMux
    port map (
            O => \N__48956\,
            I => \N__48953\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__48953\,
            I => n12
        );

    \I__12087\ : InMux
    port map (
            O => \N__48950\,
            I => n16393
        );

    \I__12086\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48944\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__48944\,
            I => n11
        );

    \I__12084\ : InMux
    port map (
            O => \N__48941\,
            I => n16394
        );

    \I__12083\ : InMux
    port map (
            O => \N__48938\,
            I => \N__48935\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__48935\,
            I => n10
        );

    \I__12081\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48929\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__48929\,
            I => n26
        );

    \I__12079\ : InMux
    port map (
            O => \N__48926\,
            I => \bfn_16_29_0_\
        );

    \I__12078\ : InMux
    port map (
            O => \N__48923\,
            I => \N__48920\
        );

    \I__12077\ : LocalMux
    port map (
            O => \N__48920\,
            I => n25
        );

    \I__12076\ : InMux
    port map (
            O => \N__48917\,
            I => n16380
        );

    \I__12075\ : InMux
    port map (
            O => \N__48914\,
            I => \N__48911\
        );

    \I__12074\ : LocalMux
    port map (
            O => \N__48911\,
            I => n24
        );

    \I__12073\ : InMux
    port map (
            O => \N__48908\,
            I => n16381
        );

    \I__12072\ : InMux
    port map (
            O => \N__48905\,
            I => \N__48902\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__48902\,
            I => n23
        );

    \I__12070\ : InMux
    port map (
            O => \N__48899\,
            I => n16382
        );

    \I__12069\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48893\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__48893\,
            I => n22_adj_2655
        );

    \I__12067\ : InMux
    port map (
            O => \N__48890\,
            I => n16383
        );

    \I__12066\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48884\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__48884\,
            I => n21
        );

    \I__12064\ : InMux
    port map (
            O => \N__48881\,
            I => n16384
        );

    \I__12063\ : InMux
    port map (
            O => \N__48878\,
            I => \N__48875\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__48875\,
            I => n20
        );

    \I__12061\ : InMux
    port map (
            O => \N__48872\,
            I => n16385
        );

    \I__12060\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48866\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__48866\,
            I => n19
        );

    \I__12058\ : InMux
    port map (
            O => \N__48863\,
            I => n16386
        );

    \I__12057\ : InMux
    port map (
            O => \N__48860\,
            I => \N__48857\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__48857\,
            I => \N__48854\
        );

    \I__12055\ : Span4Mux_v
    port map (
            O => \N__48854\,
            I => \N__48851\
        );

    \I__12054\ : Odrv4
    port map (
            O => \N__48851\,
            I => \c0.n1_adj_2484\
        );

    \I__12053\ : CascadeMux
    port map (
            O => \N__48848\,
            I => \c0.n18414_cascade_\
        );

    \I__12052\ : InMux
    port map (
            O => \N__48845\,
            I => \N__48841\
        );

    \I__12051\ : InMux
    port map (
            O => \N__48844\,
            I => \N__48834\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__48841\,
            I => \N__48830\
        );

    \I__12049\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48825\
        );

    \I__12048\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48825\
        );

    \I__12047\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48822\
        );

    \I__12046\ : InMux
    port map (
            O => \N__48837\,
            I => \N__48819\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__48834\,
            I => \N__48816\
        );

    \I__12044\ : CascadeMux
    port map (
            O => \N__48833\,
            I => \N__48812\
        );

    \I__12043\ : Span4Mux_h
    port map (
            O => \N__48830\,
            I => \N__48808\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__48825\,
            I => \N__48805\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__48822\,
            I => \N__48801\
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__48819\,
            I => \N__48798\
        );

    \I__12039\ : Span4Mux_h
    port map (
            O => \N__48816\,
            I => \N__48795\
        );

    \I__12038\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48792\
        );

    \I__12037\ : InMux
    port map (
            O => \N__48812\,
            I => \N__48787\
        );

    \I__12036\ : InMux
    port map (
            O => \N__48811\,
            I => \N__48787\
        );

    \I__12035\ : Span4Mux_v
    port map (
            O => \N__48808\,
            I => \N__48782\
        );

    \I__12034\ : Span4Mux_h
    port map (
            O => \N__48805\,
            I => \N__48782\
        );

    \I__12033\ : InMux
    port map (
            O => \N__48804\,
            I => \N__48779\
        );

    \I__12032\ : Odrv4
    port map (
            O => \N__48801\,
            I => byte_transmit_counter_4
        );

    \I__12031\ : Odrv4
    port map (
            O => \N__48798\,
            I => byte_transmit_counter_4
        );

    \I__12030\ : Odrv4
    port map (
            O => \N__48795\,
            I => byte_transmit_counter_4
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__48792\,
            I => byte_transmit_counter_4
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__48787\,
            I => byte_transmit_counter_4
        );

    \I__12027\ : Odrv4
    port map (
            O => \N__48782\,
            I => byte_transmit_counter_4
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__48779\,
            I => byte_transmit_counter_4
        );

    \I__12025\ : CascadeMux
    port map (
            O => \N__48764\,
            I => \c0.n18417_cascade_\
        );

    \I__12024\ : CascadeMux
    port map (
            O => \N__48761\,
            I => \N__48756\
        );

    \I__12023\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48751\
        );

    \I__12022\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48748\
        );

    \I__12021\ : InMux
    port map (
            O => \N__48756\,
            I => \N__48745\
        );

    \I__12020\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48742\
        );

    \I__12019\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48739\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__48751\,
            I => \N__48733\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__48748\,
            I => \N__48730\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__48745\,
            I => \N__48725\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__48742\,
            I => \N__48725\
        );

    \I__12014\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48721\
        );

    \I__12013\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48717\
        );

    \I__12012\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48712\
        );

    \I__12011\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48712\
        );

    \I__12010\ : Span4Mux_h
    port map (
            O => \N__48733\,
            I => \N__48705\
        );

    \I__12009\ : Span4Mux_h
    port map (
            O => \N__48730\,
            I => \N__48705\
        );

    \I__12008\ : Span4Mux_h
    port map (
            O => \N__48725\,
            I => \N__48705\
        );

    \I__12007\ : InMux
    port map (
            O => \N__48724\,
            I => \N__48702\
        );

    \I__12006\ : Span4Mux_h
    port map (
            O => \N__48721\,
            I => \N__48699\
        );

    \I__12005\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48696\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__48717\,
            I => byte_transmit_counter_3
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__48712\,
            I => byte_transmit_counter_3
        );

    \I__12002\ : Odrv4
    port map (
            O => \N__48705\,
            I => byte_transmit_counter_3
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__48702\,
            I => byte_transmit_counter_3
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__48699\,
            I => byte_transmit_counter_3
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__48696\,
            I => byte_transmit_counter_3
        );

    \I__11998\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48679\
        );

    \I__11997\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48676\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__48679\,
            I => \N__48671\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__48676\,
            I => \N__48668\
        );

    \I__11994\ : InMux
    port map (
            O => \N__48675\,
            I => \N__48665\
        );

    \I__11993\ : InMux
    port map (
            O => \N__48674\,
            I => \N__48662\
        );

    \I__11992\ : Span4Mux_h
    port map (
            O => \N__48671\,
            I => \N__48657\
        );

    \I__11991\ : Span4Mux_v
    port map (
            O => \N__48668\,
            I => \N__48652\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__48665\,
            I => \N__48652\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48649\
        );

    \I__11988\ : InMux
    port map (
            O => \N__48661\,
            I => \N__48643\
        );

    \I__11987\ : InMux
    port map (
            O => \N__48660\,
            I => \N__48643\
        );

    \I__11986\ : Span4Mux_v
    port map (
            O => \N__48657\,
            I => \N__48635\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__48652\,
            I => \N__48635\
        );

    \I__11984\ : Span4Mux_h
    port map (
            O => \N__48649\,
            I => \N__48635\
        );

    \I__11983\ : InMux
    port map (
            O => \N__48648\,
            I => \N__48632\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__48643\,
            I => \N__48629\
        );

    \I__11981\ : InMux
    port map (
            O => \N__48642\,
            I => \N__48626\
        );

    \I__11980\ : Odrv4
    port map (
            O => \N__48635\,
            I => n7734
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__48632\,
            I => n7734
        );

    \I__11978\ : Odrv12
    port map (
            O => \N__48629\,
            I => n7734
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__48626\,
            I => n7734
        );

    \I__11976\ : CascadeMux
    port map (
            O => \N__48617\,
            I => \tx_data_6_N_keep_cascade_\
        );

    \I__11975\ : InMux
    port map (
            O => \N__48614\,
            I => \N__48611\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__48611\,
            I => \N__48608\
        );

    \I__11973\ : Span4Mux_h
    port map (
            O => \N__48608\,
            I => \N__48604\
        );

    \I__11972\ : InMux
    port map (
            O => \N__48607\,
            I => \N__48601\
        );

    \I__11971\ : Span4Mux_h
    port map (
            O => \N__48604\,
            I => \N__48598\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__48601\,
            I => \r_Tx_Data_6\
        );

    \I__11969\ : Odrv4
    port map (
            O => \N__48598\,
            I => \r_Tx_Data_6\
        );

    \I__11968\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48586\
        );

    \I__11967\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48583\
        );

    \I__11966\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48580\
        );

    \I__11965\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48577\
        );

    \I__11964\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48574\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__48586\,
            I => \N__48571\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__48583\,
            I => \N__48564\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__48580\,
            I => \N__48564\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__48577\,
            I => \N__48561\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__48574\,
            I => \N__48556\
        );

    \I__11958\ : Span4Mux_h
    port map (
            O => \N__48571\,
            I => \N__48556\
        );

    \I__11957\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48553\
        );

    \I__11956\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48550\
        );

    \I__11955\ : Span4Mux_h
    port map (
            O => \N__48564\,
            I => \N__48547\
        );

    \I__11954\ : Span4Mux_h
    port map (
            O => \N__48561\,
            I => \N__48542\
        );

    \I__11953\ : Span4Mux_h
    port map (
            O => \N__48556\,
            I => \N__48542\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__48553\,
            I => \c0.data_out_7__6__N_530\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__48550\,
            I => \c0.data_out_7__6__N_530\
        );

    \I__11950\ : Odrv4
    port map (
            O => \N__48547\,
            I => \c0.data_out_7__6__N_530\
        );

    \I__11949\ : Odrv4
    port map (
            O => \N__48542\,
            I => \c0.data_out_7__6__N_530\
        );

    \I__11948\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48530\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__48530\,
            I => \c0.n17949\
        );

    \I__11946\ : CascadeMux
    port map (
            O => \N__48527\,
            I => \N__48523\
        );

    \I__11945\ : InMux
    port map (
            O => \N__48526\,
            I => \N__48519\
        );

    \I__11944\ : InMux
    port map (
            O => \N__48523\,
            I => \N__48516\
        );

    \I__11943\ : InMux
    port map (
            O => \N__48522\,
            I => \N__48513\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__48519\,
            I => \N__48510\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__48516\,
            I => \N__48507\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__48513\,
            I => \N__48504\
        );

    \I__11939\ : Span4Mux_v
    port map (
            O => \N__48510\,
            I => \N__48496\
        );

    \I__11938\ : Span4Mux_v
    port map (
            O => \N__48507\,
            I => \N__48496\
        );

    \I__11937\ : Span4Mux_v
    port map (
            O => \N__48504\,
            I => \N__48493\
        );

    \I__11936\ : InMux
    port map (
            O => \N__48503\,
            I => \N__48486\
        );

    \I__11935\ : InMux
    port map (
            O => \N__48502\,
            I => \N__48486\
        );

    \I__11934\ : InMux
    port map (
            O => \N__48501\,
            I => \N__48486\
        );

    \I__11933\ : Odrv4
    port map (
            O => \N__48496\,
            I => data_out_3_6
        );

    \I__11932\ : Odrv4
    port map (
            O => \N__48493\,
            I => data_out_3_6
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__48486\,
            I => data_out_3_6
        );

    \I__11930\ : InMux
    port map (
            O => \N__48479\,
            I => \N__48476\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__48476\,
            I => \c0.n18090\
        );

    \I__11928\ : InMux
    port map (
            O => \N__48473\,
            I => \N__48470\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__48470\,
            I => \N__48454\
        );

    \I__11926\ : InMux
    port map (
            O => \N__48469\,
            I => \N__48447\
        );

    \I__11925\ : InMux
    port map (
            O => \N__48468\,
            I => \N__48447\
        );

    \I__11924\ : InMux
    port map (
            O => \N__48467\,
            I => \N__48447\
        );

    \I__11923\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48440\
        );

    \I__11922\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48440\
        );

    \I__11921\ : InMux
    port map (
            O => \N__48464\,
            I => \N__48440\
        );

    \I__11920\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48433\
        );

    \I__11919\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48433\
        );

    \I__11918\ : InMux
    port map (
            O => \N__48461\,
            I => \N__48433\
        );

    \I__11917\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48422\
        );

    \I__11916\ : InMux
    port map (
            O => \N__48459\,
            I => \N__48404\
        );

    \I__11915\ : InMux
    port map (
            O => \N__48458\,
            I => \N__48404\
        );

    \I__11914\ : InMux
    port map (
            O => \N__48457\,
            I => \N__48404\
        );

    \I__11913\ : Span4Mux_s3_v
    port map (
            O => \N__48454\,
            I => \N__48385\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__48447\,
            I => \N__48385\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__48440\,
            I => \N__48385\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__48433\,
            I => \N__48385\
        );

    \I__11909\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48378\
        );

    \I__11908\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48378\
        );

    \I__11907\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48378\
        );

    \I__11906\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48373\
        );

    \I__11905\ : InMux
    port map (
            O => \N__48428\,
            I => \N__48368\
        );

    \I__11904\ : InMux
    port map (
            O => \N__48427\,
            I => \N__48368\
        );

    \I__11903\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48365\
        );

    \I__11902\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48362\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48359\
        );

    \I__11900\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48354\
        );

    \I__11899\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48354\
        );

    \I__11898\ : InMux
    port map (
            O => \N__48419\,
            I => \N__48349\
        );

    \I__11897\ : InMux
    port map (
            O => \N__48418\,
            I => \N__48349\
        );

    \I__11896\ : InMux
    port map (
            O => \N__48417\,
            I => \N__48344\
        );

    \I__11895\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48344\
        );

    \I__11894\ : InMux
    port map (
            O => \N__48415\,
            I => \N__48333\
        );

    \I__11893\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48333\
        );

    \I__11892\ : InMux
    port map (
            O => \N__48413\,
            I => \N__48333\
        );

    \I__11891\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48333\
        );

    \I__11890\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48333\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__48404\,
            I => \N__48330\
        );

    \I__11888\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48325\
        );

    \I__11887\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48325\
        );

    \I__11886\ : InMux
    port map (
            O => \N__48401\,
            I => \N__48318\
        );

    \I__11885\ : InMux
    port map (
            O => \N__48400\,
            I => \N__48318\
        );

    \I__11884\ : InMux
    port map (
            O => \N__48399\,
            I => \N__48318\
        );

    \I__11883\ : CascadeMux
    port map (
            O => \N__48398\,
            I => \N__48315\
        );

    \I__11882\ : InMux
    port map (
            O => \N__48397\,
            I => \N__48307\
        );

    \I__11881\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48307\
        );

    \I__11880\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48303\
        );

    \I__11879\ : InMux
    port map (
            O => \N__48394\,
            I => \N__48300\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__48385\,
            I => \N__48295\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48295\
        );

    \I__11876\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48292\
        );

    \I__11875\ : InMux
    port map (
            O => \N__48376\,
            I => \N__48289\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48284\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__48368\,
            I => \N__48284\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__48365\,
            I => \N__48281\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__48362\,
            I => \N__48274\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__48359\,
            I => \N__48274\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__48354\,
            I => \N__48274\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__48349\,
            I => \N__48261\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__48344\,
            I => \N__48261\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__48333\,
            I => \N__48261\
        );

    \I__11865\ : Span4Mux_h
    port map (
            O => \N__48330\,
            I => \N__48261\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__48325\,
            I => \N__48261\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__48318\,
            I => \N__48261\
        );

    \I__11862\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48258\
        );

    \I__11861\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48255\
        );

    \I__11860\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48250\
        );

    \I__11859\ : InMux
    port map (
            O => \N__48312\,
            I => \N__48250\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__48307\,
            I => \N__48247\
        );

    \I__11857\ : InMux
    port map (
            O => \N__48306\,
            I => \N__48244\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__48303\,
            I => \N__48237\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__48300\,
            I => \N__48237\
        );

    \I__11854\ : Span4Mux_h
    port map (
            O => \N__48295\,
            I => \N__48237\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__48292\,
            I => \N__48222\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__48289\,
            I => \N__48222\
        );

    \I__11851\ : Span4Mux_h
    port map (
            O => \N__48284\,
            I => \N__48222\
        );

    \I__11850\ : Span4Mux_v
    port map (
            O => \N__48281\,
            I => \N__48222\
        );

    \I__11849\ : Span4Mux_v
    port map (
            O => \N__48274\,
            I => \N__48222\
        );

    \I__11848\ : Span4Mux_v
    port map (
            O => \N__48261\,
            I => \N__48222\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__48258\,
            I => \N__48222\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__48255\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__48250\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11844\ : Odrv12
    port map (
            O => \N__48247\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__48244\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11842\ : Odrv4
    port map (
            O => \N__48237\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11841\ : Odrv4
    port map (
            O => \N__48222\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__11840\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48205\
        );

    \I__11839\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48202\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__48205\,
            I => \N__48199\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__48202\,
            I => \N__48195\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__48199\,
            I => \N__48192\
        );

    \I__11835\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48189\
        );

    \I__11834\ : Odrv4
    port map (
            O => \N__48195\,
            I => \c0.data_out_7_6\
        );

    \I__11833\ : Odrv4
    port map (
            O => \N__48192\,
            I => \c0.data_out_7_6\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__48189\,
            I => \c0.data_out_7_6\
        );

    \I__11831\ : CascadeMux
    port map (
            O => \N__48182\,
            I => \N__48179\
        );

    \I__11830\ : InMux
    port map (
            O => \N__48179\,
            I => \N__48176\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__48176\,
            I => \c0.n5_adj_2444\
        );

    \I__11828\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48170\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__48170\,
            I => \N__48167\
        );

    \I__11826\ : Odrv4
    port map (
            O => \N__48167\,
            I => \c0.n8_adj_2539\
        );

    \I__11825\ : CascadeMux
    port map (
            O => \N__48164\,
            I => \N__48160\
        );

    \I__11824\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48152\
        );

    \I__11823\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48145\
        );

    \I__11822\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48140\
        );

    \I__11821\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48140\
        );

    \I__11820\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48137\
        );

    \I__11819\ : CascadeMux
    port map (
            O => \N__48156\,
            I => \N__48130\
        );

    \I__11818\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48126\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__48152\,
            I => \N__48123\
        );

    \I__11816\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48116\
        );

    \I__11815\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48116\
        );

    \I__11814\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48116\
        );

    \I__11813\ : InMux
    port map (
            O => \N__48148\,
            I => \N__48113\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__48145\,
            I => \N__48103\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48100\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48097\
        );

    \I__11809\ : InMux
    port map (
            O => \N__48136\,
            I => \N__48092\
        );

    \I__11808\ : InMux
    port map (
            O => \N__48135\,
            I => \N__48092\
        );

    \I__11807\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48089\
        );

    \I__11806\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48082\
        );

    \I__11805\ : InMux
    port map (
            O => \N__48130\,
            I => \N__48082\
        );

    \I__11804\ : InMux
    port map (
            O => \N__48129\,
            I => \N__48082\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__48126\,
            I => \N__48077\
        );

    \I__11802\ : Span4Mux_v
    port map (
            O => \N__48123\,
            I => \N__48072\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__48116\,
            I => \N__48072\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48069\
        );

    \I__11799\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48066\
        );

    \I__11798\ : InMux
    port map (
            O => \N__48111\,
            I => \N__48061\
        );

    \I__11797\ : InMux
    port map (
            O => \N__48110\,
            I => \N__48061\
        );

    \I__11796\ : InMux
    port map (
            O => \N__48109\,
            I => \N__48056\
        );

    \I__11795\ : InMux
    port map (
            O => \N__48108\,
            I => \N__48056\
        );

    \I__11794\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48051\
        );

    \I__11793\ : InMux
    port map (
            O => \N__48106\,
            I => \N__48051\
        );

    \I__11792\ : Span4Mux_v
    port map (
            O => \N__48103\,
            I => \N__48038\
        );

    \I__11791\ : Span4Mux_h
    port map (
            O => \N__48100\,
            I => \N__48038\
        );

    \I__11790\ : Span4Mux_v
    port map (
            O => \N__48097\,
            I => \N__48038\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__48092\,
            I => \N__48038\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__48089\,
            I => \N__48038\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__48082\,
            I => \N__48038\
        );

    \I__11786\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48033\
        );

    \I__11785\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48033\
        );

    \I__11784\ : Span4Mux_v
    port map (
            O => \N__48077\,
            I => \N__48024\
        );

    \I__11783\ : Span4Mux_h
    port map (
            O => \N__48072\,
            I => \N__48024\
        );

    \I__11782\ : Span4Mux_v
    port map (
            O => \N__48069\,
            I => \N__48024\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__48066\,
            I => \N__48024\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__48061\,
            I => \N__48021\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__48056\,
            I => \N__48018\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__48051\,
            I => \N__48013\
        );

    \I__11777\ : Span4Mux_h
    port map (
            O => \N__48038\,
            I => \N__48013\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__48033\,
            I => \N__48008\
        );

    \I__11775\ : Span4Mux_h
    port map (
            O => \N__48024\,
            I => \N__48008\
        );

    \I__11774\ : Odrv4
    port map (
            O => \N__48021\,
            I => byte_transmit_counter_2
        );

    \I__11773\ : Odrv12
    port map (
            O => \N__48018\,
            I => byte_transmit_counter_2
        );

    \I__11772\ : Odrv4
    port map (
            O => \N__48013\,
            I => byte_transmit_counter_2
        );

    \I__11771\ : Odrv4
    port map (
            O => \N__48008\,
            I => byte_transmit_counter_2
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__47999\,
            I => \N__47996\
        );

    \I__11769\ : InMux
    port map (
            O => \N__47996\,
            I => \N__47993\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__47993\,
            I => \N__47990\
        );

    \I__11767\ : Odrv12
    port map (
            O => \N__47990\,
            I => \c0.n18062\
        );

    \I__11766\ : InMux
    port map (
            O => \N__47987\,
            I => \N__47978\
        );

    \I__11765\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47975\
        );

    \I__11764\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47964\
        );

    \I__11763\ : InMux
    port map (
            O => \N__47984\,
            I => \N__47961\
        );

    \I__11762\ : InMux
    port map (
            O => \N__47983\,
            I => \N__47958\
        );

    \I__11761\ : InMux
    port map (
            O => \N__47982\,
            I => \N__47953\
        );

    \I__11760\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47950\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__47978\,
            I => \N__47947\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__47975\,
            I => \N__47944\
        );

    \I__11757\ : InMux
    port map (
            O => \N__47974\,
            I => \N__47941\
        );

    \I__11756\ : InMux
    port map (
            O => \N__47973\,
            I => \N__47934\
        );

    \I__11755\ : InMux
    port map (
            O => \N__47972\,
            I => \N__47934\
        );

    \I__11754\ : InMux
    port map (
            O => \N__47971\,
            I => \N__47934\
        );

    \I__11753\ : InMux
    port map (
            O => \N__47970\,
            I => \N__47931\
        );

    \I__11752\ : CascadeMux
    port map (
            O => \N__47969\,
            I => \N__47927\
        );

    \I__11751\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47922\
        );

    \I__11750\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47922\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__47964\,
            I => \N__47919\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__47961\,
            I => \N__47916\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__47958\,
            I => \N__47913\
        );

    \I__11746\ : InMux
    port map (
            O => \N__47957\,
            I => \N__47908\
        );

    \I__11745\ : InMux
    port map (
            O => \N__47956\,
            I => \N__47908\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__47953\,
            I => \N__47903\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__47950\,
            I => \N__47903\
        );

    \I__11742\ : Span4Mux_h
    port map (
            O => \N__47947\,
            I => \N__47894\
        );

    \I__11741\ : Span4Mux_v
    port map (
            O => \N__47944\,
            I => \N__47894\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__47941\,
            I => \N__47894\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__47934\,
            I => \N__47894\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__47931\,
            I => \N__47891\
        );

    \I__11737\ : InMux
    port map (
            O => \N__47930\,
            I => \N__47887\
        );

    \I__11736\ : InMux
    port map (
            O => \N__47927\,
            I => \N__47884\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__47922\,
            I => \N__47881\
        );

    \I__11734\ : Span4Mux_h
    port map (
            O => \N__47919\,
            I => \N__47876\
        );

    \I__11733\ : Span4Mux_h
    port map (
            O => \N__47916\,
            I => \N__47876\
        );

    \I__11732\ : Span4Mux_h
    port map (
            O => \N__47913\,
            I => \N__47871\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__47908\,
            I => \N__47871\
        );

    \I__11730\ : Span4Mux_v
    port map (
            O => \N__47903\,
            I => \N__47864\
        );

    \I__11729\ : Span4Mux_h
    port map (
            O => \N__47894\,
            I => \N__47864\
        );

    \I__11728\ : Span4Mux_h
    port map (
            O => \N__47891\,
            I => \N__47864\
        );

    \I__11727\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47861\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__47887\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__47884\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11724\ : Odrv12
    port map (
            O => \N__47881\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11723\ : Odrv4
    port map (
            O => \N__47876\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11722\ : Odrv4
    port map (
            O => \N__47871\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__47864\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__47861\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__11719\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47843\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__47843\,
            I => \c0.n18063\
        );

    \I__11717\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47837\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__47837\,
            I => \N__47834\
        );

    \I__11715\ : Span4Mux_h
    port map (
            O => \N__47834\,
            I => \N__47830\
        );

    \I__11714\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47827\
        );

    \I__11713\ : Span4Mux_h
    port map (
            O => \N__47830\,
            I => \N__47822\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__47827\,
            I => \N__47819\
        );

    \I__11711\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47814\
        );

    \I__11710\ : InMux
    port map (
            O => \N__47825\,
            I => \N__47814\
        );

    \I__11709\ : Odrv4
    port map (
            O => \N__47822\,
            I => data_out_8_0
        );

    \I__11708\ : Odrv4
    port map (
            O => \N__47819\,
            I => data_out_8_0
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__47814\,
            I => data_out_8_0
        );

    \I__11706\ : InMux
    port map (
            O => \N__47807\,
            I => \N__47804\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__47804\,
            I => \N__47801\
        );

    \I__11704\ : Span4Mux_h
    port map (
            O => \N__47801\,
            I => \N__47796\
        );

    \I__11703\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47793\
        );

    \I__11702\ : InMux
    port map (
            O => \N__47799\,
            I => \N__47790\
        );

    \I__11701\ : Odrv4
    port map (
            O => \N__47796\,
            I => \c0.data_out_7_7\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__47793\,
            I => \c0.data_out_7_7\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__47790\,
            I => \c0.data_out_7_7\
        );

    \I__11698\ : CascadeMux
    port map (
            O => \N__47783\,
            I => \N__47780\
        );

    \I__11697\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47774\
        );

    \I__11696\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47774\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__47774\,
            I => \c0.n17638\
        );

    \I__11694\ : InMux
    port map (
            O => \N__47771\,
            I => \N__47763\
        );

    \I__11693\ : InMux
    port map (
            O => \N__47770\,
            I => \N__47760\
        );

    \I__11692\ : InMux
    port map (
            O => \N__47769\,
            I => \N__47757\
        );

    \I__11691\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47754\
        );

    \I__11690\ : InMux
    port map (
            O => \N__47767\,
            I => \N__47750\
        );

    \I__11689\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47747\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47744\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47741\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__47757\,
            I => \N__47736\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__47754\,
            I => \N__47736\
        );

    \I__11684\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47733\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__47750\,
            I => \N__47730\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__47747\,
            I => \N__47723\
        );

    \I__11681\ : Span4Mux_v
    port map (
            O => \N__47744\,
            I => \N__47723\
        );

    \I__11680\ : Span4Mux_v
    port map (
            O => \N__47741\,
            I => \N__47723\
        );

    \I__11679\ : Span4Mux_v
    port map (
            O => \N__47736\,
            I => \N__47720\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__47733\,
            I => \c0.data_out_0_6\
        );

    \I__11677\ : Odrv4
    port map (
            O => \N__47730\,
            I => \c0.data_out_0_6\
        );

    \I__11676\ : Odrv4
    port map (
            O => \N__47723\,
            I => \c0.data_out_0_6\
        );

    \I__11675\ : Odrv4
    port map (
            O => \N__47720\,
            I => \c0.data_out_0_6\
        );

    \I__11674\ : CascadeMux
    port map (
            O => \N__47711\,
            I => \N__47708\
        );

    \I__11673\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47705\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__47705\,
            I => \N__47700\
        );

    \I__11671\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47697\
        );

    \I__11670\ : InMux
    port map (
            O => \N__47703\,
            I => \N__47692\
        );

    \I__11669\ : Span4Mux_v
    port map (
            O => \N__47700\,
            I => \N__47687\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47687\
        );

    \I__11667\ : InMux
    port map (
            O => \N__47696\,
            I => \N__47684\
        );

    \I__11666\ : InMux
    port map (
            O => \N__47695\,
            I => \N__47681\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__47692\,
            I => \N__47674\
        );

    \I__11664\ : Span4Mux_h
    port map (
            O => \N__47687\,
            I => \N__47674\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__47684\,
            I => \N__47674\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__47681\,
            I => \N__47671\
        );

    \I__11661\ : Span4Mux_v
    port map (
            O => \N__47674\,
            I => \N__47664\
        );

    \I__11660\ : Span4Mux_h
    port map (
            O => \N__47671\,
            I => \N__47664\
        );

    \I__11659\ : InMux
    port map (
            O => \N__47670\,
            I => \N__47661\
        );

    \I__11658\ : InMux
    port map (
            O => \N__47669\,
            I => \N__47658\
        );

    \I__11657\ : Span4Mux_h
    port map (
            O => \N__47664\,
            I => \N__47655\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__47661\,
            I => data_out_0_3
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__47658\,
            I => data_out_0_3
        );

    \I__11654\ : Odrv4
    port map (
            O => \N__47655\,
            I => data_out_0_3
        );

    \I__11653\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47645\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__47645\,
            I => \N__47641\
        );

    \I__11651\ : InMux
    port map (
            O => \N__47644\,
            I => \N__47637\
        );

    \I__11650\ : Span4Mux_v
    port map (
            O => \N__47641\,
            I => \N__47632\
        );

    \I__11649\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47629\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47626\
        );

    \I__11647\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47623\
        );

    \I__11646\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47620\
        );

    \I__11645\ : Span4Mux_h
    port map (
            O => \N__47632\,
            I => \N__47616\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__47629\,
            I => \N__47613\
        );

    \I__11643\ : Span4Mux_v
    port map (
            O => \N__47626\,
            I => \N__47610\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__47623\,
            I => \N__47605\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__47620\,
            I => \N__47605\
        );

    \I__11640\ : InMux
    port map (
            O => \N__47619\,
            I => \N__47602\
        );

    \I__11639\ : Span4Mux_v
    port map (
            O => \N__47616\,
            I => \N__47599\
        );

    \I__11638\ : Span4Mux_v
    port map (
            O => \N__47613\,
            I => \N__47596\
        );

    \I__11637\ : Span4Mux_v
    port map (
            O => \N__47610\,
            I => \N__47591\
        );

    \I__11636\ : Span4Mux_v
    port map (
            O => \N__47605\,
            I => \N__47591\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__47602\,
            I => \N__47584\
        );

    \I__11634\ : Span4Mux_h
    port map (
            O => \N__47599\,
            I => \N__47584\
        );

    \I__11633\ : Span4Mux_v
    port map (
            O => \N__47596\,
            I => \N__47584\
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__47591\,
            I => data_out_0_1
        );

    \I__11631\ : Odrv4
    port map (
            O => \N__47584\,
            I => data_out_0_1
        );

    \I__11630\ : InMux
    port map (
            O => \N__47579\,
            I => \N__47574\
        );

    \I__11629\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47571\
        );

    \I__11628\ : InMux
    port map (
            O => \N__47577\,
            I => \N__47568\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__47574\,
            I => \N__47565\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__47571\,
            I => \N__47562\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__47568\,
            I => \N__47558\
        );

    \I__11624\ : Span4Mux_s2_v
    port map (
            O => \N__47565\,
            I => \N__47553\
        );

    \I__11623\ : Span4Mux_s2_v
    port map (
            O => \N__47562\,
            I => \N__47553\
        );

    \I__11622\ : InMux
    port map (
            O => \N__47561\,
            I => \N__47550\
        );

    \I__11621\ : Span4Mux_v
    port map (
            O => \N__47558\,
            I => \N__47547\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__47553\,
            I => \N__47544\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__47550\,
            I => data_out_0_0
        );

    \I__11618\ : Odrv4
    port map (
            O => \N__47547\,
            I => data_out_0_0
        );

    \I__11617\ : Odrv4
    port map (
            O => \N__47544\,
            I => data_out_0_0
        );

    \I__11616\ : CascadeMux
    port map (
            O => \N__47537\,
            I => \N__47534\
        );

    \I__11615\ : InMux
    port map (
            O => \N__47534\,
            I => \N__47530\
        );

    \I__11614\ : InMux
    port map (
            O => \N__47533\,
            I => \N__47526\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__47530\,
            I => \N__47523\
        );

    \I__11612\ : InMux
    port map (
            O => \N__47529\,
            I => \N__47520\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__47526\,
            I => \N__47513\
        );

    \I__11610\ : Span4Mux_s1_v
    port map (
            O => \N__47523\,
            I => \N__47513\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__47520\,
            I => \N__47513\
        );

    \I__11608\ : Span4Mux_v
    port map (
            O => \N__47513\,
            I => \N__47510\
        );

    \I__11607\ : Odrv4
    port map (
            O => \N__47510\,
            I => \c0.n8926\
        );

    \I__11606\ : InMux
    port map (
            O => \N__47507\,
            I => \N__47504\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__47504\,
            I => \c0.n8767\
        );

    \I__11604\ : CascadeMux
    port map (
            O => \N__47501\,
            I => \c0.n8926_cascade_\
        );

    \I__11603\ : CascadeMux
    port map (
            O => \N__47498\,
            I => \N__47495\
        );

    \I__11602\ : InMux
    port map (
            O => \N__47495\,
            I => \N__47489\
        );

    \I__11601\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47489\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__47489\,
            I => \N__47485\
        );

    \I__11599\ : InMux
    port map (
            O => \N__47488\,
            I => \N__47482\
        );

    \I__11598\ : Span4Mux_h
    port map (
            O => \N__47485\,
            I => \N__47477\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__47482\,
            I => \N__47477\
        );

    \I__11596\ : Span4Mux_h
    port map (
            O => \N__47477\,
            I => \N__47473\
        );

    \I__11595\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47470\
        );

    \I__11594\ : Odrv4
    port map (
            O => \N__47473\,
            I => n2720
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__47470\,
            I => n2720
        );

    \I__11592\ : CascadeMux
    port map (
            O => \N__47465\,
            I => \N__47462\
        );

    \I__11591\ : InMux
    port map (
            O => \N__47462\,
            I => \N__47458\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__47461\,
            I => \N__47455\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47431\
        );

    \I__11588\ : InMux
    port map (
            O => \N__47455\,
            I => \N__47428\
        );

    \I__11587\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47421\
        );

    \I__11586\ : InMux
    port map (
            O => \N__47453\,
            I => \N__47421\
        );

    \I__11585\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47421\
        );

    \I__11584\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47416\
        );

    \I__11583\ : InMux
    port map (
            O => \N__47450\,
            I => \N__47416\
        );

    \I__11582\ : CascadeMux
    port map (
            O => \N__47449\,
            I => \N__47406\
        );

    \I__11581\ : InMux
    port map (
            O => \N__47448\,
            I => \N__47386\
        );

    \I__11580\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47386\
        );

    \I__11579\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47386\
        );

    \I__11578\ : InMux
    port map (
            O => \N__47445\,
            I => \N__47386\
        );

    \I__11577\ : InMux
    port map (
            O => \N__47444\,
            I => \N__47386\
        );

    \I__11576\ : InMux
    port map (
            O => \N__47443\,
            I => \N__47375\
        );

    \I__11575\ : InMux
    port map (
            O => \N__47442\,
            I => \N__47375\
        );

    \I__11574\ : InMux
    port map (
            O => \N__47441\,
            I => \N__47375\
        );

    \I__11573\ : InMux
    port map (
            O => \N__47440\,
            I => \N__47375\
        );

    \I__11572\ : InMux
    port map (
            O => \N__47439\,
            I => \N__47375\
        );

    \I__11571\ : InMux
    port map (
            O => \N__47438\,
            I => \N__47368\
        );

    \I__11570\ : InMux
    port map (
            O => \N__47437\,
            I => \N__47368\
        );

    \I__11569\ : InMux
    port map (
            O => \N__47436\,
            I => \N__47368\
        );

    \I__11568\ : InMux
    port map (
            O => \N__47435\,
            I => \N__47363\
        );

    \I__11567\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47363\
        );

    \I__11566\ : Span4Mux_v
    port map (
            O => \N__47431\,
            I => \N__47356\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__47428\,
            I => \N__47356\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__47421\,
            I => \N__47356\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__47416\,
            I => \N__47353\
        );

    \I__11562\ : InMux
    port map (
            O => \N__47415\,
            I => \N__47348\
        );

    \I__11561\ : InMux
    port map (
            O => \N__47414\,
            I => \N__47348\
        );

    \I__11560\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47343\
        );

    \I__11559\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47343\
        );

    \I__11558\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47338\
        );

    \I__11557\ : InMux
    port map (
            O => \N__47410\,
            I => \N__47333\
        );

    \I__11556\ : InMux
    port map (
            O => \N__47409\,
            I => \N__47333\
        );

    \I__11555\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47330\
        );

    \I__11554\ : InMux
    port map (
            O => \N__47405\,
            I => \N__47327\
        );

    \I__11553\ : InMux
    port map (
            O => \N__47404\,
            I => \N__47322\
        );

    \I__11552\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47322\
        );

    \I__11551\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47317\
        );

    \I__11550\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47317\
        );

    \I__11549\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47312\
        );

    \I__11548\ : InMux
    port map (
            O => \N__47399\,
            I => \N__47312\
        );

    \I__11547\ : InMux
    port map (
            O => \N__47398\,
            I => \N__47307\
        );

    \I__11546\ : InMux
    port map (
            O => \N__47397\,
            I => \N__47307\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__47386\,
            I => \N__47302\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__47375\,
            I => \N__47302\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47284\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__47363\,
            I => \N__47284\
        );

    \I__11541\ : Span4Mux_s1_v
    port map (
            O => \N__47356\,
            I => \N__47284\
        );

    \I__11540\ : Span4Mux_s1_v
    port map (
            O => \N__47353\,
            I => \N__47284\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__47348\,
            I => \N__47284\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__47343\,
            I => \N__47280\
        );

    \I__11537\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47277\
        );

    \I__11536\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47272\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__47338\,
            I => \N__47259\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__47333\,
            I => \N__47259\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__47330\,
            I => \N__47259\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47259\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47259\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__47317\,
            I => \N__47259\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__47312\,
            I => \N__47252\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__47307\,
            I => \N__47252\
        );

    \I__11527\ : Span4Mux_s3_v
    port map (
            O => \N__47302\,
            I => \N__47252\
        );

    \I__11526\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47243\
        );

    \I__11525\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47243\
        );

    \I__11524\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47243\
        );

    \I__11523\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47243\
        );

    \I__11522\ : InMux
    port map (
            O => \N__47297\,
            I => \N__47237\
        );

    \I__11521\ : InMux
    port map (
            O => \N__47296\,
            I => \N__47230\
        );

    \I__11520\ : InMux
    port map (
            O => \N__47295\,
            I => \N__47230\
        );

    \I__11519\ : Span4Mux_v
    port map (
            O => \N__47284\,
            I => \N__47226\
        );

    \I__11518\ : InMux
    port map (
            O => \N__47283\,
            I => \N__47223\
        );

    \I__11517\ : Span4Mux_v
    port map (
            O => \N__47280\,
            I => \N__47220\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__47277\,
            I => \N__47217\
        );

    \I__11515\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47212\
        );

    \I__11514\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47212\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__47272\,
            I => \N__47203\
        );

    \I__11512\ : Span4Mux_s3_v
    port map (
            O => \N__47259\,
            I => \N__47203\
        );

    \I__11511\ : Span4Mux_h
    port map (
            O => \N__47252\,
            I => \N__47203\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__47243\,
            I => \N__47203\
        );

    \I__11509\ : InMux
    port map (
            O => \N__47242\,
            I => \N__47200\
        );

    \I__11508\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47197\
        );

    \I__11507\ : InMux
    port map (
            O => \N__47240\,
            I => \N__47194\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47191\
        );

    \I__11505\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47188\
        );

    \I__11504\ : InMux
    port map (
            O => \N__47235\,
            I => \N__47185\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__47230\,
            I => \N__47182\
        );

    \I__11502\ : InMux
    port map (
            O => \N__47229\,
            I => \N__47179\
        );

    \I__11501\ : Span4Mux_v
    port map (
            O => \N__47226\,
            I => \N__47170\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__47223\,
            I => \N__47170\
        );

    \I__11499\ : Span4Mux_v
    port map (
            O => \N__47220\,
            I => \N__47170\
        );

    \I__11498\ : Span4Mux_v
    port map (
            O => \N__47217\,
            I => \N__47170\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47163\
        );

    \I__11496\ : Span4Mux_v
    port map (
            O => \N__47203\,
            I => \N__47163\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__47200\,
            I => \N__47163\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__47197\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__47194\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11492\ : Odrv12
    port map (
            O => \N__47191\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__47188\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__47185\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11489\ : Odrv4
    port map (
            O => \N__47182\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__47179\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11487\ : Odrv4
    port map (
            O => \N__47170\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11486\ : Odrv4
    port map (
            O => \N__47163\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11485\ : SRMux
    port map (
            O => \N__47144\,
            I => \N__47138\
        );

    \I__11484\ : CascadeMux
    port map (
            O => \N__47143\,
            I => \N__47131\
        );

    \I__11483\ : CascadeMux
    port map (
            O => \N__47142\,
            I => \N__47128\
        );

    \I__11482\ : CascadeMux
    port map (
            O => \N__47141\,
            I => \N__47123\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__47138\,
            I => \N__47119\
        );

    \I__11480\ : InMux
    port map (
            O => \N__47137\,
            I => \N__47112\
        );

    \I__11479\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47112\
        );

    \I__11478\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47112\
        );

    \I__11477\ : CascadeMux
    port map (
            O => \N__47134\,
            I => \N__47107\
        );

    \I__11476\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47103\
        );

    \I__11475\ : InMux
    port map (
            O => \N__47128\,
            I => \N__47100\
        );

    \I__11474\ : CascadeMux
    port map (
            O => \N__47127\,
            I => \N__47097\
        );

    \I__11473\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47094\
        );

    \I__11472\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47089\
        );

    \I__11471\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47089\
        );

    \I__11470\ : Span4Mux_h
    port map (
            O => \N__47119\,
            I => \N__47086\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47083\
        );

    \I__11468\ : CascadeMux
    port map (
            O => \N__47111\,
            I => \N__47080\
        );

    \I__11467\ : InMux
    port map (
            O => \N__47110\,
            I => \N__47074\
        );

    \I__11466\ : InMux
    port map (
            O => \N__47107\,
            I => \N__47071\
        );

    \I__11465\ : InMux
    port map (
            O => \N__47106\,
            I => \N__47068\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__47103\,
            I => \N__47065\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47062\
        );

    \I__11462\ : InMux
    port map (
            O => \N__47097\,
            I => \N__47059\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__47094\,
            I => \N__47054\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47054\
        );

    \I__11459\ : Span4Mux_v
    port map (
            O => \N__47086\,
            I => \N__47049\
        );

    \I__11458\ : Span4Mux_s3_v
    port map (
            O => \N__47083\,
            I => \N__47049\
        );

    \I__11457\ : InMux
    port map (
            O => \N__47080\,
            I => \N__47044\
        );

    \I__11456\ : InMux
    port map (
            O => \N__47079\,
            I => \N__47044\
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__47078\,
            I => \N__47041\
        );

    \I__11454\ : CascadeMux
    port map (
            O => \N__47077\,
            I => \N__47036\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__47074\,
            I => \N__47033\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__47071\,
            I => \N__47030\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__47068\,
            I => \N__47027\
        );

    \I__11450\ : Span4Mux_h
    port map (
            O => \N__47065\,
            I => \N__47022\
        );

    \I__11449\ : Span4Mux_h
    port map (
            O => \N__47062\,
            I => \N__47022\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__47059\,
            I => \N__47019\
        );

    \I__11447\ : Span4Mux_s2_v
    port map (
            O => \N__47054\,
            I => \N__47016\
        );

    \I__11446\ : Sp12to4
    port map (
            O => \N__47049\,
            I => \N__47011\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__47044\,
            I => \N__47011\
        );

    \I__11444\ : InMux
    port map (
            O => \N__47041\,
            I => \N__47004\
        );

    \I__11443\ : InMux
    port map (
            O => \N__47040\,
            I => \N__47004\
        );

    \I__11442\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47004\
        );

    \I__11441\ : InMux
    port map (
            O => \N__47036\,
            I => \N__47001\
        );

    \I__11440\ : Span4Mux_s1_v
    port map (
            O => \N__47033\,
            I => \N__46992\
        );

    \I__11439\ : Span4Mux_h
    port map (
            O => \N__47030\,
            I => \N__46992\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__47027\,
            I => \N__46992\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__47022\,
            I => \N__46992\
        );

    \I__11436\ : Odrv12
    port map (
            O => \N__47019\,
            I => n4430
        );

    \I__11435\ : Odrv4
    port map (
            O => \N__47016\,
            I => n4430
        );

    \I__11434\ : Odrv12
    port map (
            O => \N__47011\,
            I => n4430
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__47004\,
            I => n4430
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__47001\,
            I => n4430
        );

    \I__11431\ : Odrv4
    port map (
            O => \N__46992\,
            I => n4430
        );

    \I__11430\ : InMux
    port map (
            O => \N__46979\,
            I => \N__46973\
        );

    \I__11429\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46970\
        );

    \I__11428\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46965\
        );

    \I__11427\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46965\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__46973\,
            I => \N__46962\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__46970\,
            I => data_out_1_6
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__46965\,
            I => data_out_1_6
        );

    \I__11423\ : Odrv12
    port map (
            O => \N__46962\,
            I => data_out_1_6
        );

    \I__11422\ : InMux
    port map (
            O => \N__46955\,
            I => \N__46951\
        );

    \I__11421\ : InMux
    port map (
            O => \N__46954\,
            I => \N__46946\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__46951\,
            I => \N__46943\
        );

    \I__11419\ : InMux
    port map (
            O => \N__46950\,
            I => \N__46940\
        );

    \I__11418\ : InMux
    port map (
            O => \N__46949\,
            I => \N__46937\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46934\
        );

    \I__11416\ : Span4Mux_h
    port map (
            O => \N__46943\,
            I => \N__46931\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__46940\,
            I => \N__46928\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__46937\,
            I => data_out_3_5
        );

    \I__11413\ : Odrv4
    port map (
            O => \N__46934\,
            I => data_out_3_5
        );

    \I__11412\ : Odrv4
    port map (
            O => \N__46931\,
            I => data_out_3_5
        );

    \I__11411\ : Odrv4
    port map (
            O => \N__46928\,
            I => data_out_3_5
        );

    \I__11410\ : CascadeMux
    port map (
            O => \N__46919\,
            I => \N__46911\
        );

    \I__11409\ : CascadeMux
    port map (
            O => \N__46918\,
            I => \N__46908\
        );

    \I__11408\ : CascadeMux
    port map (
            O => \N__46917\,
            I => \N__46904\
        );

    \I__11407\ : CascadeMux
    port map (
            O => \N__46916\,
            I => \N__46885\
        );

    \I__11406\ : CascadeMux
    port map (
            O => \N__46915\,
            I => \N__46874\
        );

    \I__11405\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46866\
        );

    \I__11404\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46863\
        );

    \I__11403\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46858\
        );

    \I__11402\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46858\
        );

    \I__11401\ : InMux
    port map (
            O => \N__46904\,
            I => \N__46855\
        );

    \I__11400\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46848\
        );

    \I__11399\ : InMux
    port map (
            O => \N__46902\,
            I => \N__46848\
        );

    \I__11398\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46848\
        );

    \I__11397\ : InMux
    port map (
            O => \N__46900\,
            I => \N__46845\
        );

    \I__11396\ : InMux
    port map (
            O => \N__46899\,
            I => \N__46842\
        );

    \I__11395\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46837\
        );

    \I__11394\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46837\
        );

    \I__11393\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46830\
        );

    \I__11392\ : InMux
    port map (
            O => \N__46895\,
            I => \N__46830\
        );

    \I__11391\ : InMux
    port map (
            O => \N__46894\,
            I => \N__46830\
        );

    \I__11390\ : InMux
    port map (
            O => \N__46893\,
            I => \N__46825\
        );

    \I__11389\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46825\
        );

    \I__11388\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46820\
        );

    \I__11387\ : InMux
    port map (
            O => \N__46890\,
            I => \N__46820\
        );

    \I__11386\ : InMux
    port map (
            O => \N__46889\,
            I => \N__46815\
        );

    \I__11385\ : InMux
    port map (
            O => \N__46888\,
            I => \N__46815\
        );

    \I__11384\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46812\
        );

    \I__11383\ : InMux
    port map (
            O => \N__46884\,
            I => \N__46805\
        );

    \I__11382\ : InMux
    port map (
            O => \N__46883\,
            I => \N__46805\
        );

    \I__11381\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46805\
        );

    \I__11380\ : CascadeMux
    port map (
            O => \N__46881\,
            I => \N__46801\
        );

    \I__11379\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46796\
        );

    \I__11378\ : CascadeMux
    port map (
            O => \N__46879\,
            I => \N__46790\
        );

    \I__11377\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46780\
        );

    \I__11376\ : InMux
    port map (
            O => \N__46877\,
            I => \N__46780\
        );

    \I__11375\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46773\
        );

    \I__11374\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46773\
        );

    \I__11373\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46773\
        );

    \I__11372\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46766\
        );

    \I__11371\ : InMux
    port map (
            O => \N__46870\,
            I => \N__46766\
        );

    \I__11370\ : InMux
    port map (
            O => \N__46869\,
            I => \N__46766\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__46866\,
            I => \N__46759\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__46863\,
            I => \N__46759\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__46858\,
            I => \N__46759\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__46855\,
            I => \N__46756\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46753\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46744\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__46842\,
            I => \N__46744\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__46837\,
            I => \N__46744\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__46830\,
            I => \N__46744\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46733\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__46820\,
            I => \N__46733\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__46815\,
            I => \N__46733\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__46812\,
            I => \N__46733\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__46805\,
            I => \N__46733\
        );

    \I__11355\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46730\
        );

    \I__11354\ : InMux
    port map (
            O => \N__46801\,
            I => \N__46725\
        );

    \I__11353\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46725\
        );

    \I__11352\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46720\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__46796\,
            I => \N__46717\
        );

    \I__11350\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46714\
        );

    \I__11349\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46711\
        );

    \I__11348\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46706\
        );

    \I__11347\ : InMux
    port map (
            O => \N__46790\,
            I => \N__46706\
        );

    \I__11346\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46703\
        );

    \I__11345\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46698\
        );

    \I__11344\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46698\
        );

    \I__11343\ : InMux
    port map (
            O => \N__46786\,
            I => \N__46691\
        );

    \I__11342\ : InMux
    port map (
            O => \N__46785\,
            I => \N__46688\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__46780\,
            I => \N__46673\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46673\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__46766\,
            I => \N__46673\
        );

    \I__11338\ : Span4Mux_s2_v
    port map (
            O => \N__46759\,
            I => \N__46673\
        );

    \I__11337\ : Span4Mux_h
    port map (
            O => \N__46756\,
            I => \N__46673\
        );

    \I__11336\ : Span4Mux_h
    port map (
            O => \N__46753\,
            I => \N__46673\
        );

    \I__11335\ : Span4Mux_s2_v
    port map (
            O => \N__46744\,
            I => \N__46673\
        );

    \I__11334\ : Span4Mux_s3_v
    port map (
            O => \N__46733\,
            I => \N__46667\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__46730\,
            I => \N__46662\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__46725\,
            I => \N__46662\
        );

    \I__11331\ : InMux
    port map (
            O => \N__46724\,
            I => \N__46657\
        );

    \I__11330\ : InMux
    port map (
            O => \N__46723\,
            I => \N__46657\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46654\
        );

    \I__11328\ : Span4Mux_v
    port map (
            O => \N__46717\,
            I => \N__46647\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46647\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__46711\,
            I => \N__46647\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__46706\,
            I => \N__46642\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__46703\,
            I => \N__46637\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__46698\,
            I => \N__46637\
        );

    \I__11322\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46628\
        );

    \I__11321\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46628\
        );

    \I__11320\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46628\
        );

    \I__11319\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46628\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46624\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__46688\,
            I => \N__46621\
        );

    \I__11316\ : Span4Mux_v
    port map (
            O => \N__46673\,
            I => \N__46618\
        );

    \I__11315\ : InMux
    port map (
            O => \N__46672\,
            I => \N__46611\
        );

    \I__11314\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46611\
        );

    \I__11313\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46611\
        );

    \I__11312\ : Span4Mux_h
    port map (
            O => \N__46667\,
            I => \N__46606\
        );

    \I__11311\ : Span4Mux_s3_v
    port map (
            O => \N__46662\,
            I => \N__46606\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__46657\,
            I => \N__46599\
        );

    \I__11309\ : Span4Mux_v
    port map (
            O => \N__46654\,
            I => \N__46599\
        );

    \I__11308\ : Span4Mux_h
    port map (
            O => \N__46647\,
            I => \N__46599\
        );

    \I__11307\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46594\
        );

    \I__11306\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46594\
        );

    \I__11305\ : Span4Mux_h
    port map (
            O => \N__46642\,
            I => \N__46587\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__46637\,
            I => \N__46587\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__46628\,
            I => \N__46587\
        );

    \I__11302\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46584\
        );

    \I__11301\ : Odrv12
    port map (
            O => \N__46624\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11300\ : Odrv12
    port map (
            O => \N__46621\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__46618\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__46611\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11297\ : Odrv4
    port map (
            O => \N__46606\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11296\ : Odrv4
    port map (
            O => \N__46599\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__46594\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11294\ : Odrv4
    port map (
            O => \N__46587\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__46584\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__11292\ : CEMux
    port map (
            O => \N__46565\,
            I => \N__46561\
        );

    \I__11291\ : CEMux
    port map (
            O => \N__46564\,
            I => \N__46558\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46554\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__46558\,
            I => \N__46551\
        );

    \I__11288\ : CEMux
    port map (
            O => \N__46557\,
            I => \N__46548\
        );

    \I__11287\ : Span4Mux_s1_v
    port map (
            O => \N__46554\,
            I => \N__46539\
        );

    \I__11286\ : Span4Mux_h
    port map (
            O => \N__46551\,
            I => \N__46539\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46539\
        );

    \I__11284\ : CEMux
    port map (
            O => \N__46547\,
            I => \N__46535\
        );

    \I__11283\ : CEMux
    port map (
            O => \N__46546\,
            I => \N__46532\
        );

    \I__11282\ : Span4Mux_h
    port map (
            O => \N__46539\,
            I => \N__46528\
        );

    \I__11281\ : CEMux
    port map (
            O => \N__46538\,
            I => \N__46525\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__46535\,
            I => \N__46520\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__46532\,
            I => \N__46517\
        );

    \I__11278\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46513\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__46528\,
            I => \N__46508\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__46525\,
            I => \N__46508\
        );

    \I__11275\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46503\
        );

    \I__11274\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46503\
        );

    \I__11273\ : Span4Mux_v
    port map (
            O => \N__46520\,
            I => \N__46499\
        );

    \I__11272\ : Span4Mux_v
    port map (
            O => \N__46517\,
            I => \N__46496\
        );

    \I__11271\ : CEMux
    port map (
            O => \N__46516\,
            I => \N__46493\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__46513\,
            I => \N__46490\
        );

    \I__11269\ : Span4Mux_h
    port map (
            O => \N__46508\,
            I => \N__46485\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46485\
        );

    \I__11267\ : CascadeMux
    port map (
            O => \N__46502\,
            I => \N__46481\
        );

    \I__11266\ : Span4Mux_h
    port map (
            O => \N__46499\,
            I => \N__46478\
        );

    \I__11265\ : Sp12to4
    port map (
            O => \N__46496\,
            I => \N__46475\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__46493\,
            I => \N__46472\
        );

    \I__11263\ : Span4Mux_h
    port map (
            O => \N__46490\,
            I => \N__46467\
        );

    \I__11262\ : Span4Mux_s1_v
    port map (
            O => \N__46485\,
            I => \N__46467\
        );

    \I__11261\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46462\
        );

    \I__11260\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46462\
        );

    \I__11259\ : Odrv4
    port map (
            O => \N__46478\,
            I => n9519
        );

    \I__11258\ : Odrv12
    port map (
            O => \N__46475\,
            I => n9519
        );

    \I__11257\ : Odrv4
    port map (
            O => \N__46472\,
            I => n9519
        );

    \I__11256\ : Odrv4
    port map (
            O => \N__46467\,
            I => n9519
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__46462\,
            I => n9519
        );

    \I__11254\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46442\
        );

    \I__11253\ : InMux
    port map (
            O => \N__46450\,
            I => \N__46442\
        );

    \I__11252\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46435\
        );

    \I__11251\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46435\
        );

    \I__11250\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46432\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__46442\,
            I => \N__46429\
        );

    \I__11248\ : InMux
    port map (
            O => \N__46441\,
            I => \N__46426\
        );

    \I__11247\ : InMux
    port map (
            O => \N__46440\,
            I => \N__46423\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__46435\,
            I => \N__46416\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__46432\,
            I => \N__46416\
        );

    \I__11244\ : Span4Mux_s2_v
    port map (
            O => \N__46429\,
            I => \N__46416\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46413\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__46423\,
            I => \N__46409\
        );

    \I__11241\ : Span4Mux_h
    port map (
            O => \N__46416\,
            I => \N__46406\
        );

    \I__11240\ : Span4Mux_h
    port map (
            O => \N__46413\,
            I => \N__46403\
        );

    \I__11239\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46400\
        );

    \I__11238\ : Span12Mux_h
    port map (
            O => \N__46409\,
            I => \N__46397\
        );

    \I__11237\ : Span4Mux_v
    port map (
            O => \N__46406\,
            I => \N__46394\
        );

    \I__11236\ : Span4Mux_v
    port map (
            O => \N__46403\,
            I => \N__46391\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__46400\,
            I => \data_out_5__7__N_931\
        );

    \I__11234\ : Odrv12
    port map (
            O => \N__46397\,
            I => \data_out_5__7__N_931\
        );

    \I__11233\ : Odrv4
    port map (
            O => \N__46394\,
            I => \data_out_5__7__N_931\
        );

    \I__11232\ : Odrv4
    port map (
            O => \N__46391\,
            I => \data_out_5__7__N_931\
        );

    \I__11231\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46379\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__46379\,
            I => \N__46375\
        );

    \I__11229\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46372\
        );

    \I__11228\ : Odrv4
    port map (
            O => \N__46375\,
            I => \c0.data_out_6__4__N_765\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__46372\,
            I => \c0.data_out_6__4__N_765\
        );

    \I__11226\ : InMux
    port map (
            O => \N__46367\,
            I => \N__46361\
        );

    \I__11225\ : InMux
    port map (
            O => \N__46366\,
            I => \N__46358\
        );

    \I__11224\ : CascadeMux
    port map (
            O => \N__46365\,
            I => \N__46355\
        );

    \I__11223\ : InMux
    port map (
            O => \N__46364\,
            I => \N__46352\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__46361\,
            I => \N__46349\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__46358\,
            I => \N__46346\
        );

    \I__11220\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46343\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__46352\,
            I => \N__46340\
        );

    \I__11218\ : Span4Mux_h
    port map (
            O => \N__46349\,
            I => \N__46335\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__46346\,
            I => \N__46335\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__46343\,
            I => \c0.data_out_7_2\
        );

    \I__11215\ : Odrv12
    port map (
            O => \N__46340\,
            I => \c0.data_out_7_2\
        );

    \I__11214\ : Odrv4
    port map (
            O => \N__46335\,
            I => \c0.data_out_7_2\
        );

    \I__11213\ : CascadeMux
    port map (
            O => \N__46328\,
            I => \N__46325\
        );

    \I__11212\ : InMux
    port map (
            O => \N__46325\,
            I => \N__46322\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__46322\,
            I => \N__46319\
        );

    \I__11210\ : Odrv12
    port map (
            O => \N__46319\,
            I => \c0.n17600\
        );

    \I__11209\ : InMux
    port map (
            O => \N__46316\,
            I => \N__46313\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__46313\,
            I => \c0.data_out_9_6\
        );

    \I__11207\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46306\
        );

    \I__11206\ : InMux
    port map (
            O => \N__46309\,
            I => \N__46303\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__46306\,
            I => \N__46297\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__46303\,
            I => \N__46297\
        );

    \I__11203\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46294\
        );

    \I__11202\ : Span4Mux_h
    port map (
            O => \N__46297\,
            I => \N__46291\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__46294\,
            I => \c0.data_out_7_1\
        );

    \I__11200\ : Odrv4
    port map (
            O => \N__46291\,
            I => \c0.data_out_7_1\
        );

    \I__11199\ : InMux
    port map (
            O => \N__46286\,
            I => \N__46283\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__46283\,
            I => \c0.n17454\
        );

    \I__11197\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46276\
        );

    \I__11196\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46272\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__46276\,
            I => \N__46269\
        );

    \I__11194\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46266\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__46272\,
            I => \N__46261\
        );

    \I__11192\ : Span4Mux_h
    port map (
            O => \N__46269\,
            I => \N__46261\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__46266\,
            I => \c0.data_out_6_5\
        );

    \I__11190\ : Odrv4
    port map (
            O => \N__46261\,
            I => \c0.data_out_6_5\
        );

    \I__11189\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46252\
        );

    \I__11188\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46249\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__46252\,
            I => \c0.data_out_6__5__N_752\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__46249\,
            I => \c0.data_out_6__5__N_752\
        );

    \I__11185\ : CascadeMux
    port map (
            O => \N__46244\,
            I => \c0.n17454_cascade_\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46241\,
            I => \N__46238\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__46238\,
            I => \c0.data_out_9_5\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46232\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__46232\,
            I => \N__46229\
        );

    \I__11180\ : Span4Mux_h
    port map (
            O => \N__46229\,
            I => \N__46226\
        );

    \I__11179\ : Odrv4
    port map (
            O => \N__46226\,
            I => \c0.n8_adj_2537\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46223\,
            I => \N__46220\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__46220\,
            I => \N__46216\
        );

    \I__11176\ : CascadeMux
    port map (
            O => \N__46219\,
            I => \N__46213\
        );

    \I__11175\ : Span4Mux_s3_v
    port map (
            O => \N__46216\,
            I => \N__46210\
        );

    \I__11174\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46207\
        );

    \I__11173\ : Span4Mux_h
    port map (
            O => \N__46210\,
            I => \N__46204\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__46207\,
            I => \c0.n17626\
        );

    \I__11171\ : Odrv4
    port map (
            O => \N__46204\,
            I => \c0.n17626\
        );

    \I__11170\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46195\
        );

    \I__11169\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46192\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46195\,
            I => \N__46189\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__46192\,
            I => \c0.n17608\
        );

    \I__11166\ : Odrv4
    port map (
            O => \N__46189\,
            I => \c0.n17608\
        );

    \I__11165\ : CascadeMux
    port map (
            O => \N__46184\,
            I => \N__46180\
        );

    \I__11164\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46177\
        );

    \I__11163\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46174\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__46177\,
            I => \N__46169\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__46174\,
            I => \N__46169\
        );

    \I__11160\ : Span4Mux_h
    port map (
            O => \N__46169\,
            I => \N__46166\
        );

    \I__11159\ : Odrv4
    port map (
            O => \N__46166\,
            I => \c0.n8970\
        );

    \I__11158\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46160\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__46160\,
            I => \N__46157\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__46157\,
            I => \N__46154\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__46154\,
            I => \c0.n17662\
        );

    \I__11154\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46143\
        );

    \I__11153\ : InMux
    port map (
            O => \N__46150\,
            I => \N__46143\
        );

    \I__11152\ : InMux
    port map (
            O => \N__46149\,
            I => \N__46138\
        );

    \I__11151\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46138\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46135\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__46138\,
            I => \N__46131\
        );

    \I__11148\ : Span4Mux_h
    port map (
            O => \N__46135\,
            I => \N__46128\
        );

    \I__11147\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46125\
        );

    \I__11146\ : Span4Mux_v
    port map (
            O => \N__46131\,
            I => \N__46122\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__46128\,
            I => \N__46119\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__46125\,
            I => data_out_8_6
        );

    \I__11143\ : Odrv4
    port map (
            O => \N__46122\,
            I => data_out_8_6
        );

    \I__11142\ : Odrv4
    port map (
            O => \N__46119\,
            I => data_out_8_6
        );

    \I__11141\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46109\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__46109\,
            I => \N__46106\
        );

    \I__11139\ : Span4Mux_v
    port map (
            O => \N__46106\,
            I => \N__46102\
        );

    \I__11138\ : InMux
    port map (
            O => \N__46105\,
            I => \N__46099\
        );

    \I__11137\ : Sp12to4
    port map (
            O => \N__46102\,
            I => \N__46094\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__46099\,
            I => \N__46094\
        );

    \I__11135\ : Odrv12
    port map (
            O => \N__46094\,
            I => \c0.n17665\
        );

    \I__11134\ : CascadeMux
    port map (
            O => \N__46091\,
            I => \c0.n12_adj_2482_cascade_\
        );

    \I__11133\ : InMux
    port map (
            O => \N__46088\,
            I => \N__46083\
        );

    \I__11132\ : InMux
    port map (
            O => \N__46087\,
            I => \N__46080\
        );

    \I__11131\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46076\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46073\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__46080\,
            I => \N__46070\
        );

    \I__11128\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46067\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__46076\,
            I => \N__46064\
        );

    \I__11126\ : Span4Mux_h
    port map (
            O => \N__46073\,
            I => \N__46057\
        );

    \I__11125\ : Span4Mux_v
    port map (
            O => \N__46070\,
            I => \N__46057\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__46067\,
            I => \N__46057\
        );

    \I__11123\ : Span4Mux_h
    port map (
            O => \N__46064\,
            I => \N__46054\
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__46057\,
            I => \c0.data_out_7_3\
        );

    \I__11121\ : Odrv4
    port map (
            O => \N__46054\,
            I => \c0.data_out_7_3\
        );

    \I__11120\ : InMux
    port map (
            O => \N__46049\,
            I => \N__46042\
        );

    \I__11119\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46042\
        );

    \I__11118\ : CEMux
    port map (
            O => \N__46047\,
            I => \N__46038\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__46042\,
            I => \N__46026\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46041\,
            I => \N__46023\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__46038\,
            I => \N__46019\
        );

    \I__11114\ : CEMux
    port map (
            O => \N__46037\,
            I => \N__46016\
        );

    \I__11113\ : CEMux
    port map (
            O => \N__46036\,
            I => \N__46012\
        );

    \I__11112\ : CEMux
    port map (
            O => \N__46035\,
            I => \N__46009\
        );

    \I__11111\ : CEMux
    port map (
            O => \N__46034\,
            I => \N__46005\
        );

    \I__11110\ : InMux
    port map (
            O => \N__46033\,
            I => \N__46002\
        );

    \I__11109\ : InMux
    port map (
            O => \N__46032\,
            I => \N__45995\
        );

    \I__11108\ : InMux
    port map (
            O => \N__46031\,
            I => \N__45995\
        );

    \I__11107\ : InMux
    port map (
            O => \N__46030\,
            I => \N__45995\
        );

    \I__11106\ : CEMux
    port map (
            O => \N__46029\,
            I => \N__45992\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__46026\,
            I => \N__45987\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__46023\,
            I => \N__45987\
        );

    \I__11103\ : InMux
    port map (
            O => \N__46022\,
            I => \N__45984\
        );

    \I__11102\ : Span4Mux_h
    port map (
            O => \N__46019\,
            I => \N__45981\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__46016\,
            I => \N__45978\
        );

    \I__11100\ : CEMux
    port map (
            O => \N__46015\,
            I => \N__45975\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__46012\,
            I => \N__45970\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__46009\,
            I => \N__45970\
        );

    \I__11097\ : CEMux
    port map (
            O => \N__46008\,
            I => \N__45967\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45964\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45959\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__45995\,
            I => \N__45959\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__45992\,
            I => \N__45952\
        );

    \I__11092\ : Span4Mux_h
    port map (
            O => \N__45987\,
            I => \N__45952\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__45984\,
            I => \N__45952\
        );

    \I__11090\ : Span4Mux_v
    port map (
            O => \N__45981\,
            I => \N__45949\
        );

    \I__11089\ : Span4Mux_v
    port map (
            O => \N__45978\,
            I => \N__45942\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__45975\,
            I => \N__45942\
        );

    \I__11087\ : Span4Mux_v
    port map (
            O => \N__45970\,
            I => \N__45942\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__45967\,
            I => \N__45939\
        );

    \I__11085\ : Span4Mux_h
    port map (
            O => \N__45964\,
            I => \N__45934\
        );

    \I__11084\ : Span4Mux_v
    port map (
            O => \N__45959\,
            I => \N__45934\
        );

    \I__11083\ : Span4Mux_v
    port map (
            O => \N__45952\,
            I => \N__45931\
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__45949\,
            I => \data_out_10__7__N_114\
        );

    \I__11081\ : Odrv4
    port map (
            O => \N__45942\,
            I => \data_out_10__7__N_114\
        );

    \I__11080\ : Odrv12
    port map (
            O => \N__45939\,
            I => \data_out_10__7__N_114\
        );

    \I__11079\ : Odrv4
    port map (
            O => \N__45934\,
            I => \data_out_10__7__N_114\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__45931\,
            I => \data_out_10__7__N_114\
        );

    \I__11077\ : InMux
    port map (
            O => \N__45920\,
            I => \N__45917\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__45917\,
            I => \c0.data_out_9_7\
        );

    \I__11075\ : InMux
    port map (
            O => \N__45914\,
            I => \N__45908\
        );

    \I__11074\ : InMux
    port map (
            O => \N__45913\,
            I => \N__45905\
        );

    \I__11073\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45900\
        );

    \I__11072\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45900\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__45908\,
            I => \N__45896\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__45905\,
            I => \N__45891\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__45900\,
            I => \N__45891\
        );

    \I__11068\ : InMux
    port map (
            O => \N__45899\,
            I => \N__45888\
        );

    \I__11067\ : Span4Mux_v
    port map (
            O => \N__45896\,
            I => \N__45883\
        );

    \I__11066\ : Span4Mux_v
    port map (
            O => \N__45891\,
            I => \N__45883\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45878\
        );

    \I__11064\ : Span4Mux_h
    port map (
            O => \N__45883\,
            I => \N__45878\
        );

    \I__11063\ : Odrv4
    port map (
            O => \N__45878\,
            I => data_out_8_7
        );

    \I__11062\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45872\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__45872\,
            I => \N__45869\
        );

    \I__11060\ : Span12Mux_v
    port map (
            O => \N__45869\,
            I => \N__45866\
        );

    \I__11059\ : Odrv12
    port map (
            O => \N__45866\,
            I => \c0.n8_adj_2538\
        );

    \I__11058\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45860\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__45860\,
            I => \c0.data_out_10_5\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__45857\,
            I => \N__45854\
        );

    \I__11055\ : InMux
    port map (
            O => \N__45854\,
            I => \N__45851\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__45851\,
            I => \N__45848\
        );

    \I__11053\ : Odrv4
    port map (
            O => \N__45848\,
            I => \c0.n18064\
        );

    \I__11052\ : InMux
    port map (
            O => \N__45845\,
            I => \N__45842\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__45842\,
            I => \c0.n17668\
        );

    \I__11050\ : CascadeMux
    port map (
            O => \N__45839\,
            I => \N__45835\
        );

    \I__11049\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45831\
        );

    \I__11048\ : InMux
    port map (
            O => \N__45835\,
            I => \N__45828\
        );

    \I__11047\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45825\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__45831\,
            I => \N__45820\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__45828\,
            I => \N__45820\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__45825\,
            I => \N__45817\
        );

    \I__11043\ : Span4Mux_v
    port map (
            O => \N__45820\,
            I => \N__45814\
        );

    \I__11042\ : Span4Mux_v
    port map (
            O => \N__45817\,
            I => \N__45811\
        );

    \I__11041\ : Span4Mux_h
    port map (
            O => \N__45814\,
            I => \N__45808\
        );

    \I__11040\ : Odrv4
    port map (
            O => \N__45811\,
            I => \c0.n9087\
        );

    \I__11039\ : Odrv4
    port map (
            O => \N__45808\,
            I => \c0.n9087\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__45803\,
            I => \c0.n8_adj_2528_cascade_\
        );

    \I__11037\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45797\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__45797\,
            I => \c0.data_out_10_1\
        );

    \I__11035\ : InMux
    port map (
            O => \N__45794\,
            I => \N__45791\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__45791\,
            I => \N__45788\
        );

    \I__11033\ : Span4Mux_v
    port map (
            O => \N__45788\,
            I => \N__45785\
        );

    \I__11032\ : Span4Mux_h
    port map (
            O => \N__45785\,
            I => \N__45782\
        );

    \I__11031\ : Odrv4
    port map (
            O => \N__45782\,
            I => \c0.n17556\
        );

    \I__11030\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45775\
        );

    \I__11029\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45772\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__45775\,
            I => \N__45769\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__45772\,
            I => \N__45766\
        );

    \I__11026\ : Span4Mux_s2_v
    port map (
            O => \N__45769\,
            I => \N__45763\
        );

    \I__11025\ : Odrv4
    port map (
            O => \N__45766\,
            I => \c0.data_out_6__7__N_675\
        );

    \I__11024\ : Odrv4
    port map (
            O => \N__45763\,
            I => \c0.data_out_6__7__N_675\
        );

    \I__11023\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45755\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__45755\,
            I => \N__45752\
        );

    \I__11021\ : Odrv12
    port map (
            O => \N__45752\,
            I => \c0.data_out_10_7\
        );

    \I__11020\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45746\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__45746\,
            I => \N__45742\
        );

    \I__11018\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45739\
        );

    \I__11017\ : Span4Mux_v
    port map (
            O => \N__45742\,
            I => \N__45736\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__45739\,
            I => \N__45733\
        );

    \I__11015\ : Sp12to4
    port map (
            O => \N__45736\,
            I => \N__45728\
        );

    \I__11014\ : Span12Mux_s5_v
    port map (
            O => \N__45733\,
            I => \N__45728\
        );

    \I__11013\ : Span12Mux_h
    port map (
            O => \N__45728\,
            I => \N__45725\
        );

    \I__11012\ : Odrv12
    port map (
            O => \N__45725\,
            I => \c0.n8600\
        );

    \I__11011\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45718\
        );

    \I__11010\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45714\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__45718\,
            I => \N__45710\
        );

    \I__11008\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45707\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__45714\,
            I => \N__45704\
        );

    \I__11006\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45701\
        );

    \I__11005\ : Span4Mux_v
    port map (
            O => \N__45710\,
            I => \N__45696\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__45707\,
            I => \N__45696\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__45704\,
            I => \N__45691\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__45701\,
            I => \N__45691\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__45696\,
            I => \N__45688\
        );

    \I__11000\ : Span4Mux_h
    port map (
            O => \N__45691\,
            I => \N__45685\
        );

    \I__10999\ : Odrv4
    port map (
            O => \N__45688\,
            I => \c0.data_out_5_3\
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__45685\,
            I => \c0.data_out_5_3\
        );

    \I__10997\ : CascadeMux
    port map (
            O => \N__45680\,
            I => \c0.n17635_cascade_\
        );

    \I__10996\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__45674\,
            I => \N__45671\
        );

    \I__10994\ : Span4Mux_s3_v
    port map (
            O => \N__45671\,
            I => \N__45668\
        );

    \I__10993\ : Span4Mux_h
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10992\ : Odrv4
    port map (
            O => \N__45665\,
            I => \c0.n17922\
        );

    \I__10991\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__45659\,
            I => \N__45650\
        );

    \I__10989\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45647\
        );

    \I__10988\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45640\
        );

    \I__10987\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45640\
        );

    \I__10986\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45640\
        );

    \I__10985\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45635\
        );

    \I__10984\ : InMux
    port map (
            O => \N__45653\,
            I => \N__45635\
        );

    \I__10983\ : Span4Mux_h
    port map (
            O => \N__45650\,
            I => \N__45632\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__45647\,
            I => \N__45629\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45626\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__45635\,
            I => \N__45622\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__45632\,
            I => \N__45619\
        );

    \I__10978\ : Span4Mux_h
    port map (
            O => \N__45629\,
            I => \N__45614\
        );

    \I__10977\ : Span4Mux_h
    port map (
            O => \N__45626\,
            I => \N__45614\
        );

    \I__10976\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45611\
        );

    \I__10975\ : Span4Mux_h
    port map (
            O => \N__45622\,
            I => \N__45606\
        );

    \I__10974\ : Span4Mux_v
    port map (
            O => \N__45619\,
            I => \N__45606\
        );

    \I__10973\ : Odrv4
    port map (
            O => \N__45614\,
            I => \c0.data_out_7__7__N_519\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__45611\,
            I => \c0.data_out_7__7__N_519\
        );

    \I__10971\ : Odrv4
    port map (
            O => \N__45606\,
            I => \c0.data_out_7__7__N_519\
        );

    \I__10970\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45591\
        );

    \I__10969\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45591\
        );

    \I__10968\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45587\
        );

    \I__10967\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45584\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__45591\,
            I => \N__45581\
        );

    \I__10965\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45578\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__45587\,
            I => \N__45575\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45572\
        );

    \I__10962\ : Span4Mux_v
    port map (
            O => \N__45581\,
            I => \N__45565\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45565\
        );

    \I__10960\ : Span4Mux_v
    port map (
            O => \N__45575\,
            I => \N__45565\
        );

    \I__10959\ : Span4Mux_h
    port map (
            O => \N__45572\,
            I => \N__45562\
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__45565\,
            I => \c0.data_out_7_5\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__45562\,
            I => \c0.data_out_7_5\
        );

    \I__10956\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45554\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__45554\,
            I => \c0.n17492\
        );

    \I__10954\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45548\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__45548\,
            I => \c0.n17635\
        );

    \I__10952\ : CascadeMux
    port map (
            O => \N__45545\,
            I => \c0.n17492_cascade_\
        );

    \I__10951\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45539\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__45539\,
            I => \N__45536\
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__45536\,
            I => \c0.data_out_10_3\
        );

    \I__10948\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45530\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__45530\,
            I => \c0.n8_adj_2531\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__45527\,
            I => \c0.n18069_cascade_\
        );

    \I__10945\ : InMux
    port map (
            O => \N__45524\,
            I => \N__45521\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__45521\,
            I => \N__45518\
        );

    \I__10943\ : Span4Mux_h
    port map (
            O => \N__45518\,
            I => \N__45515\
        );

    \I__10942\ : Odrv4
    port map (
            O => \N__45515\,
            I => \c0.n18070\
        );

    \I__10941\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45506\
        );

    \I__10940\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45506\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__45506\,
            I => \N__45498\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__45505\,
            I => \N__45490\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__45504\,
            I => \N__45478\
        );

    \I__10936\ : CascadeMux
    port map (
            O => \N__45503\,
            I => \N__45475\
        );

    \I__10935\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45469\
        );

    \I__10934\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45469\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__45498\,
            I => \N__45466\
        );

    \I__10932\ : InMux
    port map (
            O => \N__45497\,
            I => \N__45461\
        );

    \I__10931\ : InMux
    port map (
            O => \N__45496\,
            I => \N__45461\
        );

    \I__10930\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45457\
        );

    \I__10929\ : CascadeMux
    port map (
            O => \N__45494\,
            I => \N__45448\
        );

    \I__10928\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45434\
        );

    \I__10927\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45434\
        );

    \I__10926\ : InMux
    port map (
            O => \N__45489\,
            I => \N__45434\
        );

    \I__10925\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45434\
        );

    \I__10924\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45434\
        );

    \I__10923\ : CascadeMux
    port map (
            O => \N__45486\,
            I => \N__45426\
        );

    \I__10922\ : CascadeMux
    port map (
            O => \N__45485\,
            I => \N__45423\
        );

    \I__10921\ : CascadeMux
    port map (
            O => \N__45484\,
            I => \N__45420\
        );

    \I__10920\ : CascadeMux
    port map (
            O => \N__45483\,
            I => \N__45412\
        );

    \I__10919\ : InMux
    port map (
            O => \N__45482\,
            I => \N__45406\
        );

    \I__10918\ : InMux
    port map (
            O => \N__45481\,
            I => \N__45403\
        );

    \I__10917\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45396\
        );

    \I__10916\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45396\
        );

    \I__10915\ : InMux
    port map (
            O => \N__45474\,
            I => \N__45396\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__45469\,
            I => \N__45389\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__45466\,
            I => \N__45389\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__45461\,
            I => \N__45389\
        );

    \I__10911\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45386\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__45457\,
            I => \N__45382\
        );

    \I__10909\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45375\
        );

    \I__10908\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45375\
        );

    \I__10907\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45375\
        );

    \I__10906\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45360\
        );

    \I__10905\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45360\
        );

    \I__10904\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45360\
        );

    \I__10903\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45360\
        );

    \I__10902\ : InMux
    port map (
            O => \N__45447\,
            I => \N__45360\
        );

    \I__10901\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45360\
        );

    \I__10900\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45360\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__45434\,
            I => \N__45357\
        );

    \I__10898\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45354\
        );

    \I__10897\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45331\
        );

    \I__10896\ : InMux
    port map (
            O => \N__45431\,
            I => \N__45331\
        );

    \I__10895\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45331\
        );

    \I__10894\ : InMux
    port map (
            O => \N__45429\,
            I => \N__45331\
        );

    \I__10893\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45324\
        );

    \I__10892\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45324\
        );

    \I__10891\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45317\
        );

    \I__10890\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45317\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45317\
        );

    \I__10888\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45302\
        );

    \I__10887\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45302\
        );

    \I__10886\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45302\
        );

    \I__10885\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45302\
        );

    \I__10884\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45302\
        );

    \I__10883\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45302\
        );

    \I__10882\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45302\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__45406\,
            I => \N__45299\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__45403\,
            I => \N__45296\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__45396\,
            I => \N__45284\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__45389\,
            I => \N__45284\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__45386\,
            I => \N__45284\
        );

    \I__10876\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45281\
        );

    \I__10875\ : Span4Mux_v
    port map (
            O => \N__45382\,
            I => \N__45277\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__45375\,
            I => \N__45270\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__45360\,
            I => \N__45270\
        );

    \I__10872\ : Span4Mux_v
    port map (
            O => \N__45357\,
            I => \N__45270\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45267\
        );

    \I__10870\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45264\
        );

    \I__10869\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45255\
        );

    \I__10868\ : InMux
    port map (
            O => \N__45351\,
            I => \N__45255\
        );

    \I__10867\ : InMux
    port map (
            O => \N__45350\,
            I => \N__45255\
        );

    \I__10866\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45255\
        );

    \I__10865\ : CascadeMux
    port map (
            O => \N__45348\,
            I => \N__45242\
        );

    \I__10864\ : CascadeMux
    port map (
            O => \N__45347\,
            I => \N__45239\
        );

    \I__10863\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45235\
        );

    \I__10862\ : CascadeMux
    port map (
            O => \N__45345\,
            I => \N__45228\
        );

    \I__10861\ : InMux
    port map (
            O => \N__45344\,
            I => \N__45223\
        );

    \I__10860\ : CascadeMux
    port map (
            O => \N__45343\,
            I => \N__45220\
        );

    \I__10859\ : CascadeMux
    port map (
            O => \N__45342\,
            I => \N__45217\
        );

    \I__10858\ : CascadeMux
    port map (
            O => \N__45341\,
            I => \N__45214\
        );

    \I__10857\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45193\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__45331\,
            I => \N__45190\
        );

    \I__10855\ : InMux
    port map (
            O => \N__45330\,
            I => \N__45185\
        );

    \I__10854\ : InMux
    port map (
            O => \N__45329\,
            I => \N__45185\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45178\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__45317\,
            I => \N__45178\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__45302\,
            I => \N__45178\
        );

    \I__10850\ : Span4Mux_v
    port map (
            O => \N__45299\,
            I => \N__45173\
        );

    \I__10849\ : Span4Mux_s2_h
    port map (
            O => \N__45296\,
            I => \N__45173\
        );

    \I__10848\ : InMux
    port map (
            O => \N__45295\,
            I => \N__45168\
        );

    \I__10847\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45168\
        );

    \I__10846\ : InMux
    port map (
            O => \N__45293\,
            I => \N__45165\
        );

    \I__10845\ : InMux
    port map (
            O => \N__45292\,
            I => \N__45149\
        );

    \I__10844\ : InMux
    port map (
            O => \N__45291\,
            I => \N__45146\
        );

    \I__10843\ : Span4Mux_v
    port map (
            O => \N__45284\,
            I => \N__45143\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__45281\,
            I => \N__45137\
        );

    \I__10841\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45134\
        );

    \I__10840\ : Span4Mux_h
    port map (
            O => \N__45277\,
            I => \N__45123\
        );

    \I__10839\ : Span4Mux_h
    port map (
            O => \N__45270\,
            I => \N__45123\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__45267\,
            I => \N__45123\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45123\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__45255\,
            I => \N__45123\
        );

    \I__10835\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45118\
        );

    \I__10834\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45118\
        );

    \I__10833\ : CascadeMux
    port map (
            O => \N__45252\,
            I => \N__45107\
        );

    \I__10832\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45100\
        );

    \I__10831\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45100\
        );

    \I__10830\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45093\
        );

    \I__10829\ : InMux
    port map (
            O => \N__45248\,
            I => \N__45093\
        );

    \I__10828\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45093\
        );

    \I__10827\ : InMux
    port map (
            O => \N__45246\,
            I => \N__45088\
        );

    \I__10826\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45088\
        );

    \I__10825\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45081\
        );

    \I__10824\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45081\
        );

    \I__10823\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45081\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__45235\,
            I => \N__45078\
        );

    \I__10821\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45072\
        );

    \I__10820\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45072\
        );

    \I__10819\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45069\
        );

    \I__10818\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45057\
        );

    \I__10817\ : InMux
    port map (
            O => \N__45228\,
            I => \N__45057\
        );

    \I__10816\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45057\
        );

    \I__10815\ : InMux
    port map (
            O => \N__45226\,
            I => \N__45057\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__45223\,
            I => \N__45047\
        );

    \I__10813\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45032\
        );

    \I__10812\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45032\
        );

    \I__10811\ : InMux
    port map (
            O => \N__45214\,
            I => \N__45032\
        );

    \I__10810\ : InMux
    port map (
            O => \N__45213\,
            I => \N__45032\
        );

    \I__10809\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45032\
        );

    \I__10808\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45032\
        );

    \I__10807\ : InMux
    port map (
            O => \N__45210\,
            I => \N__45032\
        );

    \I__10806\ : InMux
    port map (
            O => \N__45209\,
            I => \N__45029\
        );

    \I__10805\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45020\
        );

    \I__10804\ : InMux
    port map (
            O => \N__45207\,
            I => \N__45020\
        );

    \I__10803\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45020\
        );

    \I__10802\ : InMux
    port map (
            O => \N__45205\,
            I => \N__45020\
        );

    \I__10801\ : InMux
    port map (
            O => \N__45204\,
            I => \N__45017\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45014\
        );

    \I__10799\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45007\
        );

    \I__10798\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45007\
        );

    \I__10797\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45007\
        );

    \I__10796\ : InMux
    port map (
            O => \N__45199\,
            I => \N__45000\
        );

    \I__10795\ : InMux
    port map (
            O => \N__45198\,
            I => \N__45000\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45197\,
            I => \N__45000\
        );

    \I__10793\ : InMux
    port map (
            O => \N__45196\,
            I => \N__44997\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__45193\,
            I => \N__44984\
        );

    \I__10791\ : Span4Mux_v
    port map (
            O => \N__45190\,
            I => \N__44984\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__45185\,
            I => \N__44984\
        );

    \I__10789\ : Span4Mux_v
    port map (
            O => \N__45178\,
            I => \N__44984\
        );

    \I__10788\ : Span4Mux_h
    port map (
            O => \N__45173\,
            I => \N__44984\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__45168\,
            I => \N__44984\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__45165\,
            I => \N__44981\
        );

    \I__10785\ : InMux
    port map (
            O => \N__45164\,
            I => \N__44978\
        );

    \I__10784\ : InMux
    port map (
            O => \N__45163\,
            I => \N__44969\
        );

    \I__10783\ : InMux
    port map (
            O => \N__45162\,
            I => \N__44969\
        );

    \I__10782\ : InMux
    port map (
            O => \N__45161\,
            I => \N__44969\
        );

    \I__10781\ : InMux
    port map (
            O => \N__45160\,
            I => \N__44969\
        );

    \I__10780\ : InMux
    port map (
            O => \N__45159\,
            I => \N__44963\
        );

    \I__10779\ : InMux
    port map (
            O => \N__45158\,
            I => \N__44963\
        );

    \I__10778\ : InMux
    port map (
            O => \N__45157\,
            I => \N__44960\
        );

    \I__10777\ : InMux
    port map (
            O => \N__45156\,
            I => \N__44953\
        );

    \I__10776\ : InMux
    port map (
            O => \N__45155\,
            I => \N__44953\
        );

    \I__10775\ : InMux
    port map (
            O => \N__45154\,
            I => \N__44953\
        );

    \I__10774\ : CascadeMux
    port map (
            O => \N__45153\,
            I => \N__44941\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__45152\,
            I => \N__44938\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__45149\,
            I => \N__44929\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__45146\,
            I => \N__44929\
        );

    \I__10770\ : Span4Mux_v
    port map (
            O => \N__45143\,
            I => \N__44926\
        );

    \I__10769\ : InMux
    port map (
            O => \N__45142\,
            I => \N__44923\
        );

    \I__10768\ : InMux
    port map (
            O => \N__45141\,
            I => \N__44918\
        );

    \I__10767\ : InMux
    port map (
            O => \N__45140\,
            I => \N__44918\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__45137\,
            I => \N__44913\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__45134\,
            I => \N__44913\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__45123\,
            I => \N__44908\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__45118\,
            I => \N__44908\
        );

    \I__10762\ : InMux
    port map (
            O => \N__45117\,
            I => \N__44903\
        );

    \I__10761\ : InMux
    port map (
            O => \N__45116\,
            I => \N__44903\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45115\,
            I => \N__44899\
        );

    \I__10759\ : InMux
    port map (
            O => \N__45114\,
            I => \N__44894\
        );

    \I__10758\ : InMux
    port map (
            O => \N__45113\,
            I => \N__44894\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__45112\,
            I => \N__44891\
        );

    \I__10756\ : InMux
    port map (
            O => \N__45111\,
            I => \N__44885\
        );

    \I__10755\ : InMux
    port map (
            O => \N__45110\,
            I => \N__44876\
        );

    \I__10754\ : InMux
    port map (
            O => \N__45107\,
            I => \N__44876\
        );

    \I__10753\ : InMux
    port map (
            O => \N__45106\,
            I => \N__44876\
        );

    \I__10752\ : InMux
    port map (
            O => \N__45105\,
            I => \N__44876\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__45100\,
            I => \N__44867\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__45093\,
            I => \N__44867\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__45088\,
            I => \N__44867\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__45081\,
            I => \N__44867\
        );

    \I__10747\ : Span4Mux_v
    port map (
            O => \N__45078\,
            I => \N__44862\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45077\,
            I => \N__44859\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__44854\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__45069\,
            I => \N__44854\
        );

    \I__10743\ : InMux
    port map (
            O => \N__45068\,
            I => \N__44847\
        );

    \I__10742\ : InMux
    port map (
            O => \N__45067\,
            I => \N__44847\
        );

    \I__10741\ : InMux
    port map (
            O => \N__45066\,
            I => \N__44847\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__45057\,
            I => \N__44844\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45056\,
            I => \N__44839\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45055\,
            I => \N__44839\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45054\,
            I => \N__44836\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45053\,
            I => \N__44827\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45052\,
            I => \N__44827\
        );

    \I__10734\ : InMux
    port map (
            O => \N__45051\,
            I => \N__44827\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45050\,
            I => \N__44827\
        );

    \I__10732\ : Span4Mux_h
    port map (
            O => \N__45047\,
            I => \N__44824\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45032\,
            I => \N__44817\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__45029\,
            I => \N__44817\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__45020\,
            I => \N__44817\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__45017\,
            I => \N__44812\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45014\,
            I => \N__44812\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45007\,
            I => \N__44801\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__45000\,
            I => \N__44801\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__44997\,
            I => \N__44801\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__44984\,
            I => \N__44801\
        );

    \I__10722\ : Span4Mux_h
    port map (
            O => \N__44981\,
            I => \N__44801\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__44978\,
            I => \N__44796\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__44969\,
            I => \N__44796\
        );

    \I__10719\ : CascadeMux
    port map (
            O => \N__44968\,
            I => \N__44793\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__44963\,
            I => \N__44786\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__44960\,
            I => \N__44786\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44783\
        );

    \I__10715\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44776\
        );

    \I__10714\ : InMux
    port map (
            O => \N__44951\,
            I => \N__44776\
        );

    \I__10713\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44776\
        );

    \I__10712\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44769\
        );

    \I__10711\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44769\
        );

    \I__10710\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44769\
        );

    \I__10709\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44762\
        );

    \I__10708\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44762\
        );

    \I__10707\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44759\
        );

    \I__10706\ : InMux
    port map (
            O => \N__44941\,
            I => \N__44746\
        );

    \I__10705\ : InMux
    port map (
            O => \N__44938\,
            I => \N__44746\
        );

    \I__10704\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44746\
        );

    \I__10703\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44746\
        );

    \I__10702\ : InMux
    port map (
            O => \N__44935\,
            I => \N__44746\
        );

    \I__10701\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44746\
        );

    \I__10700\ : Span4Mux_h
    port map (
            O => \N__44929\,
            I => \N__44741\
        );

    \I__10699\ : Span4Mux_v
    port map (
            O => \N__44926\,
            I => \N__44741\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__44923\,
            I => \N__44730\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__44918\,
            I => \N__44730\
        );

    \I__10696\ : Span4Mux_h
    port map (
            O => \N__44913\,
            I => \N__44730\
        );

    \I__10695\ : Span4Mux_v
    port map (
            O => \N__44908\,
            I => \N__44730\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44730\
        );

    \I__10693\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44727\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44722\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__44894\,
            I => \N__44722\
        );

    \I__10690\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44713\
        );

    \I__10689\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44713\
        );

    \I__10688\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44713\
        );

    \I__10687\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44713\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__44885\,
            I => \N__44710\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__44876\,
            I => \N__44705\
        );

    \I__10684\ : Span4Mux_v
    port map (
            O => \N__44867\,
            I => \N__44705\
        );

    \I__10683\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44700\
        );

    \I__10682\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44700\
        );

    \I__10681\ : Span4Mux_v
    port map (
            O => \N__44862\,
            I => \N__44689\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__44859\,
            I => \N__44689\
        );

    \I__10679\ : Span4Mux_v
    port map (
            O => \N__44854\,
            I => \N__44689\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__44847\,
            I => \N__44689\
        );

    \I__10677\ : Span4Mux_h
    port map (
            O => \N__44844\,
            I => \N__44689\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__44839\,
            I => \N__44672\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__44836\,
            I => \N__44672\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__44827\,
            I => \N__44672\
        );

    \I__10673\ : Span4Mux_h
    port map (
            O => \N__44824\,
            I => \N__44672\
        );

    \I__10672\ : Span4Mux_v
    port map (
            O => \N__44817\,
            I => \N__44672\
        );

    \I__10671\ : Span4Mux_h
    port map (
            O => \N__44812\,
            I => \N__44672\
        );

    \I__10670\ : Span4Mux_v
    port map (
            O => \N__44801\,
            I => \N__44672\
        );

    \I__10669\ : Span4Mux_h
    port map (
            O => \N__44796\,
            I => \N__44672\
        );

    \I__10668\ : InMux
    port map (
            O => \N__44793\,
            I => \N__44665\
        );

    \I__10667\ : InMux
    port map (
            O => \N__44792\,
            I => \N__44665\
        );

    \I__10666\ : InMux
    port map (
            O => \N__44791\,
            I => \N__44665\
        );

    \I__10665\ : Span4Mux_h
    port map (
            O => \N__44786\,
            I => \N__44656\
        );

    \I__10664\ : Span4Mux_h
    port map (
            O => \N__44783\,
            I => \N__44656\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44656\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__44769\,
            I => \N__44656\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__44768\,
            I => \N__44653\
        );

    \I__10660\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44645\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__44762\,
            I => \N__44640\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__44759\,
            I => \N__44640\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__44746\,
            I => \N__44637\
        );

    \I__10656\ : Span4Mux_h
    port map (
            O => \N__44741\,
            I => \N__44632\
        );

    \I__10655\ : Span4Mux_v
    port map (
            O => \N__44730\,
            I => \N__44632\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__44727\,
            I => \N__44625\
        );

    \I__10653\ : Span4Mux_v
    port map (
            O => \N__44722\,
            I => \N__44625\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__44713\,
            I => \N__44625\
        );

    \I__10651\ : Span4Mux_v
    port map (
            O => \N__44710\,
            I => \N__44614\
        );

    \I__10650\ : Span4Mux_h
    port map (
            O => \N__44705\,
            I => \N__44614\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__44700\,
            I => \N__44614\
        );

    \I__10648\ : Span4Mux_h
    port map (
            O => \N__44689\,
            I => \N__44614\
        );

    \I__10647\ : Span4Mux_v
    port map (
            O => \N__44672\,
            I => \N__44614\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__44665\,
            I => \N__44609\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__44656\,
            I => \N__44609\
        );

    \I__10644\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44606\
        );

    \I__10643\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44601\
        );

    \I__10642\ : InMux
    port map (
            O => \N__44651\,
            I => \N__44601\
        );

    \I__10641\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44594\
        );

    \I__10640\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44594\
        );

    \I__10639\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44594\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__44645\,
            I => \N__44589\
        );

    \I__10637\ : Span12Mux_h
    port map (
            O => \N__44640\,
            I => \N__44589\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__44637\,
            I => \N__44584\
        );

    \I__10635\ : Span4Mux_v
    port map (
            O => \N__44632\,
            I => \N__44584\
        );

    \I__10634\ : Span4Mux_v
    port map (
            O => \N__44625\,
            I => \N__44579\
        );

    \I__10633\ : Span4Mux_v
    port map (
            O => \N__44614\,
            I => \N__44579\
        );

    \I__10632\ : Span4Mux_v
    port map (
            O => \N__44609\,
            I => \N__44576\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__44606\,
            I => rx_data_ready
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__44601\,
            I => rx_data_ready
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__44594\,
            I => rx_data_ready
        );

    \I__10628\ : Odrv12
    port map (
            O => \N__44589\,
            I => rx_data_ready
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__44584\,
            I => rx_data_ready
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__44579\,
            I => rx_data_ready
        );

    \I__10625\ : Odrv4
    port map (
            O => \N__44576\,
            I => rx_data_ready
        );

    \I__10624\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44558\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__10622\ : Span4Mux_h
    port map (
            O => \N__44555\,
            I => \N__44552\
        );

    \I__10621\ : Span4Mux_h
    port map (
            O => \N__44552\,
            I => \N__44548\
        );

    \I__10620\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44545\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__44548\,
            I => data_in_14_6
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__44545\,
            I => data_in_14_6
        );

    \I__10617\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44537\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__44537\,
            I => \N__44534\
        );

    \I__10615\ : Span4Mux_h
    port map (
            O => \N__44534\,
            I => \N__44530\
        );

    \I__10614\ : InMux
    port map (
            O => \N__44533\,
            I => \N__44527\
        );

    \I__10613\ : Odrv4
    port map (
            O => \N__44530\,
            I => data_in_13_6
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__44527\,
            I => data_in_13_6
        );

    \I__10611\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44519\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__44519\,
            I => \N__44516\
        );

    \I__10609\ : Odrv12
    port map (
            O => \N__44516\,
            I => \c0.n17445\
        );

    \I__10608\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44509\
        );

    \I__10607\ : InMux
    port map (
            O => \N__44512\,
            I => \N__44506\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__44509\,
            I => \N__44503\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44500\
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__44503\,
            I => \c0.n17510\
        );

    \I__10603\ : Odrv4
    port map (
            O => \N__44500\,
            I => \c0.n17510\
        );

    \I__10602\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44492\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__44492\,
            I => \c0.data_out_9_1\
        );

    \I__10600\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44485\
        );

    \I__10599\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44482\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__44485\,
            I => \N__44478\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__44482\,
            I => \N__44475\
        );

    \I__10596\ : InMux
    port map (
            O => \N__44481\,
            I => \N__44471\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__44478\,
            I => \N__44468\
        );

    \I__10594\ : Span4Mux_v
    port map (
            O => \N__44475\,
            I => \N__44465\
        );

    \I__10593\ : InMux
    port map (
            O => \N__44474\,
            I => \N__44462\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__44471\,
            I => data_out_8_1
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__44468\,
            I => data_out_8_1
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__44465\,
            I => data_out_8_1
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__44462\,
            I => data_out_8_1
        );

    \I__10588\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44450\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__44450\,
            I => \c0.n8_adj_2519\
        );

    \I__10586\ : InMux
    port map (
            O => \N__44447\,
            I => \N__44444\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44441\
        );

    \I__10584\ : Span4Mux_h
    port map (
            O => \N__44441\,
            I => \N__44438\
        );

    \I__10583\ : Odrv4
    port map (
            O => \N__44438\,
            I => \c0.n8_adj_2535\
        );

    \I__10582\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44432\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44429\
        );

    \I__10580\ : Span4Mux_h
    port map (
            O => \N__44429\,
            I => \N__44426\
        );

    \I__10579\ : Odrv4
    port map (
            O => \N__44426\,
            I => \c0.n17398\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__10577\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44416\
        );

    \I__10576\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44413\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__44416\,
            I => \N__44410\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44407\
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__44410\,
            I => \c0.n9091\
        );

    \I__10572\ : Odrv12
    port map (
            O => \N__44407\,
            I => \c0.n9091\
        );

    \I__10571\ : InMux
    port map (
            O => \N__44402\,
            I => \N__44399\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__44399\,
            I => \c0.data_out_9_4\
        );

    \I__10569\ : InMux
    port map (
            O => \N__44396\,
            I => \N__44392\
        );

    \I__10568\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44389\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__44392\,
            I => \N__44383\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44383\
        );

    \I__10565\ : InMux
    port map (
            O => \N__44388\,
            I => \N__44380\
        );

    \I__10564\ : Odrv4
    port map (
            O => \N__44383\,
            I => \c0.data_out_6_1\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__44380\,
            I => \c0.data_out_6_1\
        );

    \I__10562\ : CascadeMux
    port map (
            O => \N__44375\,
            I => \N__44372\
        );

    \I__10561\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44369\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__44369\,
            I => \N__44365\
        );

    \I__10559\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44362\
        );

    \I__10558\ : Span4Mux_h
    port map (
            O => \N__44365\,
            I => \N__44359\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__44362\,
            I => \c0.n17499\
        );

    \I__10556\ : Odrv4
    port map (
            O => \N__44359\,
            I => \c0.n17499\
        );

    \I__10555\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__44351\,
            I => \N__44348\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__44345\,
            I => \c0.n6_adj_2451\
        );

    \I__10551\ : CascadeMux
    port map (
            O => \N__44342\,
            I => \c0.n18065_cascade_\
        );

    \I__10550\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44336\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__44336\,
            I => \N__44333\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__44333\,
            I => \tx_data_5_N_keep\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__44330\,
            I => \N__44327\
        );

    \I__10546\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44324\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__44324\,
            I => \N__44321\
        );

    \I__10544\ : Odrv4
    port map (
            O => \N__44321\,
            I => \c0.n18014\
        );

    \I__10543\ : InMux
    port map (
            O => \N__44318\,
            I => \N__44315\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__44315\,
            I => \tx_data_1_N_keep\
        );

    \I__10541\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44309\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__44306\,
            I => \c0.n17943\
        );

    \I__10538\ : CascadeMux
    port map (
            O => \N__44303\,
            I => \c0.n5_adj_2481_cascade_\
        );

    \I__10537\ : InMux
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__44297\,
            I => \c0.n18091\
        );

    \I__10535\ : CascadeMux
    port map (
            O => \N__44294\,
            I => \c0.n18402_cascade_\
        );

    \I__10534\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__10532\ : Span4Mux_h
    port map (
            O => \N__44285\,
            I => \N__44282\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__44282\,
            I => \c0.n2_adj_2476\
        );

    \I__10530\ : InMux
    port map (
            O => \N__44279\,
            I => \N__44276\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__44276\,
            I => \c0.n18405\
        );

    \I__10528\ : InMux
    port map (
            O => \N__44273\,
            I => \N__44269\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__44272\,
            I => \N__44265\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__44269\,
            I => \N__44261\
        );

    \I__10525\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44258\
        );

    \I__10524\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44255\
        );

    \I__10523\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44252\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__44261\,
            I => \N__44247\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__44258\,
            I => \N__44247\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__44255\,
            I => \c0.data_out_5_1\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__44252\,
            I => \c0.data_out_5_1\
        );

    \I__10518\ : Odrv4
    port map (
            O => \N__44247\,
            I => \c0.data_out_5_1\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__44240\,
            I => \c0.n45_adj_2518_cascade_\
        );

    \I__10516\ : InMux
    port map (
            O => \N__44237\,
            I => \N__44234\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__44234\,
            I => \N__44231\
        );

    \I__10514\ : Odrv4
    port map (
            O => \N__44231\,
            I => \c0.n1_adj_2522\
        );

    \I__10513\ : CascadeMux
    port map (
            O => \N__44228\,
            I => \c0.n46_cascade_\
        );

    \I__10512\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44222\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__44222\,
            I => \c0.n44_adj_2524\
        );

    \I__10510\ : CascadeMux
    port map (
            O => \N__44219\,
            I => \N__44216\
        );

    \I__10509\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44213\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__44213\,
            I => \N__44210\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__44210\,
            I => \N__44206\
        );

    \I__10506\ : CascadeMux
    port map (
            O => \N__44209\,
            I => \N__44203\
        );

    \I__10505\ : Span4Mux_h
    port map (
            O => \N__44206\,
            I => \N__44200\
        );

    \I__10504\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44197\
        );

    \I__10503\ : Odrv4
    port map (
            O => \N__44200\,
            I => rand_setpoint_9
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__44197\,
            I => rand_setpoint_9
        );

    \I__10501\ : CEMux
    port map (
            O => \N__44192\,
            I => \N__44189\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44183\
        );

    \I__10499\ : CEMux
    port map (
            O => \N__44188\,
            I => \N__44180\
        );

    \I__10498\ : CEMux
    port map (
            O => \N__44187\,
            I => \N__44177\
        );

    \I__10497\ : CEMux
    port map (
            O => \N__44186\,
            I => \N__44174\
        );

    \I__10496\ : Span4Mux_h
    port map (
            O => \N__44183\,
            I => \N__44168\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__44180\,
            I => \N__44168\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__44177\,
            I => \N__44165\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44162\
        );

    \I__10492\ : CEMux
    port map (
            O => \N__44173\,
            I => \N__44159\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__44168\,
            I => \N__44156\
        );

    \I__10490\ : Sp12to4
    port map (
            O => \N__44165\,
            I => \N__44153\
        );

    \I__10489\ : Span4Mux_h
    port map (
            O => \N__44162\,
            I => \N__44148\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__44159\,
            I => \N__44148\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__44156\,
            I => \c0.n9518\
        );

    \I__10486\ : Odrv12
    port map (
            O => \N__44153\,
            I => \c0.n9518\
        );

    \I__10485\ : Odrv4
    port map (
            O => \N__44148\,
            I => \c0.n9518\
        );

    \I__10484\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44135\
        );

    \I__10483\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44132\
        );

    \I__10482\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44129\
        );

    \I__10481\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44125\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44120\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44115\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__44129\,
            I => \N__44115\
        );

    \I__10477\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44112\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__44125\,
            I => \N__44109\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44106\
        );

    \I__10474\ : InMux
    port map (
            O => \N__44123\,
            I => \N__44103\
        );

    \I__10473\ : Span4Mux_h
    port map (
            O => \N__44120\,
            I => \N__44100\
        );

    \I__10472\ : Span4Mux_v
    port map (
            O => \N__44115\,
            I => \N__44095\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44112\,
            I => \N__44095\
        );

    \I__10470\ : Odrv12
    port map (
            O => \N__44109\,
            I => \data_out_6__2__N_804\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__44106\,
            I => \data_out_6__2__N_804\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__44103\,
            I => \data_out_6__2__N_804\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__44100\,
            I => \data_out_6__2__N_804\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__44095\,
            I => \data_out_6__2__N_804\
        );

    \I__10465\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44081\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__44081\,
            I => \N__44077\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44074\
        );

    \I__10462\ : Odrv4
    port map (
            O => \N__44077\,
            I => \c0.n17457\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__44074\,
            I => \c0.n17457\
        );

    \I__10460\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44066\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__44066\,
            I => \c0.n17654\
        );

    \I__10458\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44057\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__44057\,
            I => \N__44054\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__44054\,
            I => \c0.n18061\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44051\,
            I => \N__44047\
        );

    \I__10453\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44043\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44047\,
            I => \N__44040\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44037\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__44034\
        );

    \I__10449\ : Span4Mux_s3_v
    port map (
            O => \N__44040\,
            I => \N__44029\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__44037\,
            I => \N__44029\
        );

    \I__10447\ : Span4Mux_v
    port map (
            O => \N__44034\,
            I => \N__44026\
        );

    \I__10446\ : Span4Mux_h
    port map (
            O => \N__44029\,
            I => \N__44023\
        );

    \I__10445\ : Span4Mux_h
    port map (
            O => \N__44026\,
            I => \N__44020\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__44023\,
            I => \c0.data_out_7__5__N_543\
        );

    \I__10443\ : Odrv4
    port map (
            O => \N__44020\,
            I => \c0.data_out_7__5__N_543\
        );

    \I__10442\ : InMux
    port map (
            O => \N__44015\,
            I => \N__44010\
        );

    \I__10441\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44005\
        );

    \I__10440\ : InMux
    port map (
            O => \N__44013\,
            I => \N__44005\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__44010\,
            I => \N__44002\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__44005\,
            I => \N__43995\
        );

    \I__10437\ : Span4Mux_v
    port map (
            O => \N__44002\,
            I => \N__43995\
        );

    \I__10436\ : CascadeMux
    port map (
            O => \N__44001\,
            I => \N__43991\
        );

    \I__10435\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43988\
        );

    \I__10434\ : Span4Mux_h
    port map (
            O => \N__43995\,
            I => \N__43985\
        );

    \I__10433\ : InMux
    port map (
            O => \N__43994\,
            I => \N__43980\
        );

    \I__10432\ : InMux
    port map (
            O => \N__43991\,
            I => \N__43980\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__43988\,
            I => \data_out_6__1__N_850\
        );

    \I__10430\ : Odrv4
    port map (
            O => \N__43985\,
            I => \data_out_6__1__N_850\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__43980\,
            I => \data_out_6__1__N_850\
        );

    \I__10428\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43970\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__43970\,
            I => \N__43967\
        );

    \I__10426\ : Span4Mux_v
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__10425\ : Odrv4
    port map (
            O => \N__43964\,
            I => \c0.n2\
        );

    \I__10424\ : CascadeMux
    port map (
            O => \N__43961\,
            I => \N__43958\
        );

    \I__10423\ : InMux
    port map (
            O => \N__43958\,
            I => \N__43955\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__43955\,
            I => \N__43952\
        );

    \I__10421\ : Odrv12
    port map (
            O => \N__43952\,
            I => \c0.n18060\
        );

    \I__10420\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43941\
        );

    \I__10419\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43937\
        );

    \I__10418\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43934\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__43946\,
            I => \N__43931\
        );

    \I__10416\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43926\
        );

    \I__10415\ : InMux
    port map (
            O => \N__43944\,
            I => \N__43926\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__43941\,
            I => \N__43923\
        );

    \I__10413\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43920\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__43937\,
            I => \N__43917\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__43934\,
            I => \N__43914\
        );

    \I__10410\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43911\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__43926\,
            I => \N__43906\
        );

    \I__10408\ : Span4Mux_h
    port map (
            O => \N__43923\,
            I => \N__43906\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__43920\,
            I => \N__43901\
        );

    \I__10406\ : Span12Mux_h
    port map (
            O => \N__43917\,
            I => \N__43901\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__43914\,
            I => \N__43898\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__43911\,
            I => data_out_0_5
        );

    \I__10403\ : Odrv4
    port map (
            O => \N__43906\,
            I => data_out_0_5
        );

    \I__10402\ : Odrv12
    port map (
            O => \N__43901\,
            I => data_out_0_5
        );

    \I__10401\ : Odrv4
    port map (
            O => \N__43898\,
            I => data_out_0_5
        );

    \I__10400\ : InMux
    port map (
            O => \N__43889\,
            I => \N__43886\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__43886\,
            I => \N__43883\
        );

    \I__10398\ : Span4Mux_h
    port map (
            O => \N__43883\,
            I => \N__43880\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__43880\,
            I => \N__43876\
        );

    \I__10396\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43873\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__43876\,
            I => rand_setpoint_21
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__43873\,
            I => rand_setpoint_21
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__43868\,
            I => \c0.n9656_cascade_\
        );

    \I__10392\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43862\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__43862\,
            I => \N__43859\
        );

    \I__10390\ : Span4Mux_s3_v
    port map (
            O => \N__43859\,
            I => \N__43855\
        );

    \I__10389\ : CascadeMux
    port map (
            O => \N__43858\,
            I => \N__43852\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__43855\,
            I => \N__43849\
        );

    \I__10387\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43846\
        );

    \I__10386\ : Odrv4
    port map (
            O => \N__43849\,
            I => rand_setpoint_17
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__43846\,
            I => rand_setpoint_17
        );

    \I__10384\ : CascadeMux
    port map (
            O => \N__43841\,
            I => \c0.n2251_cascade_\
        );

    \I__10383\ : InMux
    port map (
            O => \N__43838\,
            I => \N__43835\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__43835\,
            I => \N__43832\
        );

    \I__10381\ : Odrv12
    port map (
            O => \N__43832\,
            I => \c0.n17962\
        );

    \I__10380\ : CascadeMux
    port map (
            O => \N__43829\,
            I => \N__43826\
        );

    \I__10379\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43820\
        );

    \I__10378\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43820\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__43820\,
            I => \N__43817\
        );

    \I__10376\ : Span4Mux_h
    port map (
            O => \N__43817\,
            I => \N__43814\
        );

    \I__10375\ : Odrv4
    port map (
            O => \N__43814\,
            I => \c0.data_out_6__1__N_849\
        );

    \I__10374\ : InMux
    port map (
            O => \N__43811\,
            I => \N__43807\
        );

    \I__10373\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43804\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43798\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43798\
        );

    \I__10370\ : InMux
    port map (
            O => \N__43803\,
            I => \N__43793\
        );

    \I__10369\ : Span4Mux_v
    port map (
            O => \N__43798\,
            I => \N__43790\
        );

    \I__10368\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43787\
        );

    \I__10367\ : InMux
    port map (
            O => \N__43796\,
            I => \N__43784\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__43793\,
            I => \N__43777\
        );

    \I__10365\ : Span4Mux_v
    port map (
            O => \N__43790\,
            I => \N__43777\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__43787\,
            I => \N__43777\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__43784\,
            I => \c0.data_out_1_1\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__43777\,
            I => \c0.data_out_1_1\
        );

    \I__10361\ : InMux
    port map (
            O => \N__43772\,
            I => \N__43766\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__43771\,
            I => \N__43763\
        );

    \I__10359\ : CascadeMux
    port map (
            O => \N__43770\,
            I => \N__43760\
        );

    \I__10358\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43757\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__43766\,
            I => \N__43754\
        );

    \I__10356\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43751\
        );

    \I__10355\ : InMux
    port map (
            O => \N__43760\,
            I => \N__43746\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__43757\,
            I => \N__43743\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__43754\,
            I => \N__43738\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__43751\,
            I => \N__43738\
        );

    \I__10351\ : InMux
    port map (
            O => \N__43750\,
            I => \N__43733\
        );

    \I__10350\ : InMux
    port map (
            O => \N__43749\,
            I => \N__43733\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__43746\,
            I => \N__43726\
        );

    \I__10348\ : Span4Mux_v
    port map (
            O => \N__43743\,
            I => \N__43726\
        );

    \I__10347\ : Span4Mux_v
    port map (
            O => \N__43738\,
            I => \N__43726\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__43733\,
            I => data_out_1_2
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__43726\,
            I => data_out_1_2
        );

    \I__10344\ : CascadeMux
    port map (
            O => \N__43721\,
            I => \c0.n8767_cascade_\
        );

    \I__10343\ : InMux
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43712\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__43712\,
            I => \c0.n17525\
        );

    \I__10340\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43705\
        );

    \I__10339\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43702\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__43705\,
            I => \N__43699\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__43702\,
            I => \N__43696\
        );

    \I__10336\ : Span4Mux_v
    port map (
            O => \N__43699\,
            I => \N__43693\
        );

    \I__10335\ : Span4Mux_h
    port map (
            O => \N__43696\,
            I => \N__43690\
        );

    \I__10334\ : Sp12to4
    port map (
            O => \N__43693\,
            I => \N__43687\
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__43690\,
            I => \c0.n17641\
        );

    \I__10332\ : Odrv12
    port map (
            O => \N__43687\,
            I => \c0.n17641\
        );

    \I__10331\ : CascadeMux
    port map (
            O => \N__43682\,
            I => \c0.n17457_cascade_\
        );

    \I__10330\ : InMux
    port map (
            O => \N__43679\,
            I => \N__43676\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__10328\ : Span4Mux_h
    port map (
            O => \N__43673\,
            I => \N__43669\
        );

    \I__10327\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43666\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__43669\,
            I => \c0.n8964\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__43666\,
            I => \c0.n8964\
        );

    \I__10324\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43658\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__43658\,
            I => \c0.n17415\
        );

    \I__10322\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__43652\,
            I => \N__43643\
        );

    \I__10320\ : InMux
    port map (
            O => \N__43651\,
            I => \N__43640\
        );

    \I__10319\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43637\
        );

    \I__10318\ : InMux
    port map (
            O => \N__43649\,
            I => \N__43634\
        );

    \I__10317\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43631\
        );

    \I__10316\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43628\
        );

    \I__10315\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43625\
        );

    \I__10314\ : Span4Mux_h
    port map (
            O => \N__43643\,
            I => \N__43620\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__43640\,
            I => \N__43620\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__43637\,
            I => \N__43617\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__43634\,
            I => \N__43614\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__43631\,
            I => \N__43607\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__43628\,
            I => \N__43607\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__43625\,
            I => \N__43607\
        );

    \I__10307\ : Span4Mux_h
    port map (
            O => \N__43620\,
            I => \N__43604\
        );

    \I__10306\ : Span4Mux_h
    port map (
            O => \N__43617\,
            I => \N__43601\
        );

    \I__10305\ : Odrv12
    port map (
            O => \N__43614\,
            I => \c0.data_out_6__3__N_788\
        );

    \I__10304\ : Odrv12
    port map (
            O => \N__43607\,
            I => \c0.data_out_6__3__N_788\
        );

    \I__10303\ : Odrv4
    port map (
            O => \N__43604\,
            I => \c0.data_out_6__3__N_788\
        );

    \I__10302\ : Odrv4
    port map (
            O => \N__43601\,
            I => \c0.data_out_6__3__N_788\
        );

    \I__10301\ : CascadeMux
    port map (
            O => \N__43592\,
            I => \c0.n17415_cascade_\
        );

    \I__10300\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43585\
        );

    \I__10299\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43581\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43577\
        );

    \I__10297\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43574\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__43581\,
            I => \N__43571\
        );

    \I__10295\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43568\
        );

    \I__10294\ : Span4Mux_v
    port map (
            O => \N__43577\,
            I => \N__43563\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__43574\,
            I => \N__43563\
        );

    \I__10292\ : Span4Mux_h
    port map (
            O => \N__43571\,
            I => \N__43558\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43555\
        );

    \I__10290\ : Span4Mux_h
    port map (
            O => \N__43563\,
            I => \N__43552\
        );

    \I__10289\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43549\
        );

    \I__10288\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43546\
        );

    \I__10287\ : Span4Mux_v
    port map (
            O => \N__43558\,
            I => \N__43543\
        );

    \I__10286\ : Odrv4
    port map (
            O => \N__43555\,
            I => \c0.data_out_5_2\
        );

    \I__10285\ : Odrv4
    port map (
            O => \N__43552\,
            I => \c0.data_out_5_2\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__43549\,
            I => \c0.data_out_5_2\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__43546\,
            I => \c0.data_out_5_2\
        );

    \I__10282\ : Odrv4
    port map (
            O => \N__43543\,
            I => \c0.data_out_5_2\
        );

    \I__10281\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43529\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__43529\,
            I => \N__43524\
        );

    \I__10279\ : InMux
    port map (
            O => \N__43528\,
            I => \N__43521\
        );

    \I__10278\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43518\
        );

    \I__10277\ : Span4Mux_h
    port map (
            O => \N__43524\,
            I => \N__43515\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43512\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__43518\,
            I => \N__43509\
        );

    \I__10274\ : Span4Mux_v
    port map (
            O => \N__43515\,
            I => \N__43502\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__43512\,
            I => \N__43502\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__43509\,
            I => \N__43502\
        );

    \I__10271\ : Odrv4
    port map (
            O => \N__43502\,
            I => \c0.data_out_6_7\
        );

    \I__10270\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43496\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__43496\,
            I => \c0.n9195\
        );

    \I__10268\ : CascadeMux
    port map (
            O => \N__43493\,
            I => \c0.n17668_cascade_\
        );

    \I__10267\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43487\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__43487\,
            I => \N__43483\
        );

    \I__10265\ : InMux
    port map (
            O => \N__43486\,
            I => \N__43480\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__43483\,
            I => \c0.n8812\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__43480\,
            I => \c0.n8812\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__43475\,
            I => \c0.n8_adj_2511_cascade_\
        );

    \I__10261\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43469\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__43469\,
            I => \c0.n17623\
        );

    \I__10259\ : InMux
    port map (
            O => \N__43466\,
            I => \N__43462\
        );

    \I__10258\ : InMux
    port map (
            O => \N__43465\,
            I => \N__43458\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43455\
        );

    \I__10256\ : InMux
    port map (
            O => \N__43461\,
            I => \N__43452\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__43458\,
            I => \N__43449\
        );

    \I__10254\ : Span4Mux_h
    port map (
            O => \N__43455\,
            I => \N__43446\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__43452\,
            I => \c0.n8950\
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__43449\,
            I => \c0.n8950\
        );

    \I__10251\ : Odrv4
    port map (
            O => \N__43446\,
            I => \c0.n8950\
        );

    \I__10250\ : InMux
    port map (
            O => \N__43439\,
            I => \N__43436\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__43436\,
            I => \c0.data_out_9_0\
        );

    \I__10248\ : InMux
    port map (
            O => \N__43433\,
            I => \N__43430\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__43430\,
            I => \c0.data_out_10_0\
        );

    \I__10246\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43424\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__43424\,
            I => \c0.n18016\
        );

    \I__10244\ : CascadeMux
    port map (
            O => \N__43421\,
            I => \N__43417\
        );

    \I__10243\ : InMux
    port map (
            O => \N__43420\,
            I => \N__43414\
        );

    \I__10242\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43410\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43404\
        );

    \I__10240\ : InMux
    port map (
            O => \N__43413\,
            I => \N__43401\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__43410\,
            I => \N__43398\
        );

    \I__10238\ : CascadeMux
    port map (
            O => \N__43409\,
            I => \N__43395\
        );

    \I__10237\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43391\
        );

    \I__10236\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43388\
        );

    \I__10235\ : Span4Mux_v
    port map (
            O => \N__43404\,
            I => \N__43385\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__43401\,
            I => \N__43380\
        );

    \I__10233\ : Span4Mux_h
    port map (
            O => \N__43398\,
            I => \N__43380\
        );

    \I__10232\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43375\
        );

    \I__10231\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43375\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__43391\,
            I => \N__43370\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43370\
        );

    \I__10228\ : Odrv4
    port map (
            O => \N__43385\,
            I => \c0.data_out_2_3\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__43380\,
            I => \c0.data_out_2_3\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__43375\,
            I => \c0.data_out_2_3\
        );

    \I__10225\ : Odrv12
    port map (
            O => \N__43370\,
            I => \c0.data_out_2_3\
        );

    \I__10224\ : CascadeMux
    port map (
            O => \N__43361\,
            I => \c0.n4_adj_2543_cascade_\
        );

    \I__10223\ : CascadeMux
    port map (
            O => \N__43358\,
            I => \c0.n18073_cascade_\
        );

    \I__10222\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43352\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__43352\,
            I => \N__43348\
        );

    \I__10220\ : CascadeMux
    port map (
            O => \N__43351\,
            I => \N__43345\
        );

    \I__10219\ : Span12Mux_h
    port map (
            O => \N__43348\,
            I => \N__43342\
        );

    \I__10218\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43339\
        );

    \I__10217\ : Odrv12
    port map (
            O => \N__43342\,
            I => rand_setpoint_3
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__43339\,
            I => rand_setpoint_3
        );

    \I__10215\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43329\
        );

    \I__10214\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43325\
        );

    \I__10213\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43322\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__43329\,
            I => \N__43319\
        );

    \I__10211\ : InMux
    port map (
            O => \N__43328\,
            I => \N__43316\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__43325\,
            I => \N__43313\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__43322\,
            I => \N__43308\
        );

    \I__10208\ : Span4Mux_h
    port map (
            O => \N__43319\,
            I => \N__43308\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__43316\,
            I => data_out_8_2
        );

    \I__10206\ : Odrv12
    port map (
            O => \N__43313\,
            I => data_out_8_2
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__43308\,
            I => data_out_8_2
        );

    \I__10204\ : InMux
    port map (
            O => \N__43301\,
            I => \N__43297\
        );

    \I__10203\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43294\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43291\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__43294\,
            I => \N__43288\
        );

    \I__10200\ : Span4Mux_h
    port map (
            O => \N__43291\,
            I => \N__43285\
        );

    \I__10199\ : Odrv12
    port map (
            O => \N__43288\,
            I => \c0.data_out_6_4\
        );

    \I__10198\ : Odrv4
    port map (
            O => \N__43285\,
            I => \c0.data_out_6_4\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__43280\,
            I => \c0.n9091_cascade_\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__43277\,
            I => \c0.n17566_cascade_\
        );

    \I__10195\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43271\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43266\
        );

    \I__10193\ : InMux
    port map (
            O => \N__43270\,
            I => \N__43263\
        );

    \I__10192\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43260\
        );

    \I__10191\ : Span4Mux_h
    port map (
            O => \N__43266\,
            I => \N__43257\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__43263\,
            I => \N__43254\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__43260\,
            I => \N__43251\
        );

    \I__10188\ : Span4Mux_v
    port map (
            O => \N__43257\,
            I => \N__43248\
        );

    \I__10187\ : Span4Mux_h
    port map (
            O => \N__43254\,
            I => \N__43245\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__43251\,
            I => \N__43242\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__43248\,
            I => \c0.data_out_6_3\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__43245\,
            I => \c0.data_out_6_3\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__43242\,
            I => \c0.data_out_6_3\
        );

    \I__10182\ : CascadeMux
    port map (
            O => \N__43235\,
            I => \c0.n9195_cascade_\
        );

    \I__10181\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43227\
        );

    \I__10180\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43223\
        );

    \I__10179\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43220\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__43227\,
            I => \N__43217\
        );

    \I__10177\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43214\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__43223\,
            I => \N__43211\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__43220\,
            I => \c0.data_out_7__4__N_556\
        );

    \I__10174\ : Odrv4
    port map (
            O => \N__43217\,
            I => \c0.data_out_7__4__N_556\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__43214\,
            I => \c0.data_out_7__4__N_556\
        );

    \I__10172\ : Odrv12
    port map (
            O => \N__43211\,
            I => \c0.data_out_7__4__N_556\
        );

    \I__10171\ : InMux
    port map (
            O => \N__43202\,
            I => \N__43199\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__43199\,
            I => \N__43196\
        );

    \I__10169\ : Span4Mux_h
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__43193\,
            I => \c0.n18015\
        );

    \I__10167\ : CascadeMux
    port map (
            O => \N__43190\,
            I => \N__43187\
        );

    \I__10166\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__43184\,
            I => \c0.n8_adj_2516\
        );

    \I__10164\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43177\
        );

    \I__10163\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43174\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__43177\,
            I => \N__43171\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__43174\,
            I => \r_Tx_Data_1\
        );

    \I__10160\ : Odrv12
    port map (
            O => \N__43171\,
            I => \r_Tx_Data_1\
        );

    \I__10159\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__43163\,
            I => \c0.n18071\
        );

    \I__10157\ : CascadeMux
    port map (
            O => \N__43160\,
            I => \c0.n8_adj_2526_cascade_\
        );

    \I__10156\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43151\
        );

    \I__10154\ : Span4Mux_h
    port map (
            O => \N__43151\,
            I => \N__43148\
        );

    \I__10153\ : Odrv4
    port map (
            O => \N__43148\,
            I => \c0.n18072\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__43145\,
            I => \N__43142\
        );

    \I__10151\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43139\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__43139\,
            I => \N__43136\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__43136\,
            I => \N__43133\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__43133\,
            I => \N__43129\
        );

    \I__10147\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43126\
        );

    \I__10146\ : Odrv4
    port map (
            O => \N__43129\,
            I => \c0.n17644\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__43126\,
            I => \c0.n17644\
        );

    \I__10144\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43118\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__43118\,
            I => \N__43115\
        );

    \I__10142\ : Span4Mux_v
    port map (
            O => \N__43115\,
            I => \N__43112\
        );

    \I__10141\ : Odrv4
    port map (
            O => \N__43112\,
            I => \c0.data_out_7__2__N_574\
        );

    \I__10140\ : CascadeMux
    port map (
            O => \N__43109\,
            I => \c0.data_out_7__2__N_574_cascade_\
        );

    \I__10139\ : InMux
    port map (
            O => \N__43106\,
            I => \N__43103\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__43103\,
            I => \c0.data_out_10_2\
        );

    \I__10137\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43097\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__43097\,
            I => \c0.data_out_9_2\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43094\,
            I => \N__43091\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__43091\,
            I => \N__43088\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__43088\,
            I => \N__43085\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__43085\,
            I => \N__43082\
        );

    \I__10131\ : Odrv4
    port map (
            O => \N__43082\,
            I => \c0.data_out_9_3\
        );

    \I__10130\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__43076\,
            I => \c0.n2650\
        );

    \I__10128\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43070\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__43070\,
            I => \N__43065\
        );

    \I__10126\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43062\
        );

    \I__10125\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43059\
        );

    \I__10124\ : Odrv4
    port map (
            O => \N__43065\,
            I => \c0.tx_transmit_N_2239_0\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__43062\,
            I => \c0.tx_transmit_N_2239_0\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43059\,
            I => \c0.tx_transmit_N_2239_0\
        );

    \I__10121\ : InMux
    port map (
            O => \N__43052\,
            I => \N__43047\
        );

    \I__10120\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43044\
        );

    \I__10119\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43041\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43047\,
            I => \c0.tx_transmit_N_2239_1\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__43044\,
            I => \c0.tx_transmit_N_2239_1\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__43041\,
            I => \c0.tx_transmit_N_2239_1\
        );

    \I__10115\ : InMux
    port map (
            O => \N__43034\,
            I => \N__43031\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__43031\,
            I => \N__43028\
        );

    \I__10113\ : Span4Mux_h
    port map (
            O => \N__43028\,
            I => \N__43023\
        );

    \I__10112\ : InMux
    port map (
            O => \N__43027\,
            I => \N__43020\
        );

    \I__10111\ : InMux
    port map (
            O => \N__43026\,
            I => \N__43017\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__43023\,
            I => \tx_transmit_N_2239_2\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__43020\,
            I => \tx_transmit_N_2239_2\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__43017\,
            I => \tx_transmit_N_2239_2\
        );

    \I__10107\ : InMux
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__43007\,
            I => \N__43003\
        );

    \I__10105\ : InMux
    port map (
            O => \N__43006\,
            I => \N__42999\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__43003\,
            I => \N__42996\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42993\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__42999\,
            I => \c0.n97\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__42996\,
            I => \c0.n97\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__42993\,
            I => \c0.n97\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__42986\,
            I => \N__42980\
        );

    \I__10098\ : CascadeMux
    port map (
            O => \N__42985\,
            I => \N__42976\
        );

    \I__10097\ : InMux
    port map (
            O => \N__42984\,
            I => \N__42971\
        );

    \I__10096\ : InMux
    port map (
            O => \N__42983\,
            I => \N__42971\
        );

    \I__10095\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42968\
        );

    \I__10094\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42965\
        );

    \I__10093\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42962\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__42971\,
            I => \N__42959\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__42968\,
            I => \N__42956\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42951\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42951\
        );

    \I__10088\ : Span4Mux_v
    port map (
            O => \N__42959\,
            I => \N__42947\
        );

    \I__10087\ : Span12Mux_h
    port map (
            O => \N__42956\,
            I => \N__42942\
        );

    \I__10086\ : Span12Mux_h
    port map (
            O => \N__42951\,
            I => \N__42942\
        );

    \I__10085\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42939\
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__42947\,
            I => \c0.tx_transmit\
        );

    \I__10083\ : Odrv12
    port map (
            O => \N__42942\,
            I => \c0.tx_transmit\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__42939\,
            I => \c0.tx_transmit\
        );

    \I__10081\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42927\
        );

    \I__10080\ : InMux
    port map (
            O => \N__42931\,
            I => \N__42924\
        );

    \I__10079\ : InMux
    port map (
            O => \N__42930\,
            I => \N__42921\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__42927\,
            I => \N__42916\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__42924\,
            I => \N__42916\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__42921\,
            I => \N__42910\
        );

    \I__10075\ : Span4Mux_v
    port map (
            O => \N__42916\,
            I => \N__42907\
        );

    \I__10074\ : InMux
    port map (
            O => \N__42915\,
            I => \N__42900\
        );

    \I__10073\ : InMux
    port map (
            O => \N__42914\,
            I => \N__42900\
        );

    \I__10072\ : InMux
    port map (
            O => \N__42913\,
            I => \N__42900\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__42910\,
            I => tx_active
        );

    \I__10070\ : Odrv4
    port map (
            O => \N__42907\,
            I => tx_active
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__42900\,
            I => tx_active
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__42893\,
            I => \N__42889\
        );

    \I__10067\ : CascadeMux
    port map (
            O => \N__42892\,
            I => \N__42885\
        );

    \I__10066\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42881\
        );

    \I__10065\ : InMux
    port map (
            O => \N__42888\,
            I => \N__42878\
        );

    \I__10064\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42875\
        );

    \I__10063\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42871\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42867\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__42878\,
            I => \N__42862\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42862\
        );

    \I__10059\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42859\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42856\
        );

    \I__10057\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42853\
        );

    \I__10056\ : Span4Mux_v
    port map (
            O => \N__42867\,
            I => \N__42848\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__42862\,
            I => \N__42848\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__42859\,
            I => n13415
        );

    \I__10053\ : Odrv4
    port map (
            O => \N__42856\,
            I => n13415
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__42853\,
            I => n13415
        );

    \I__10051\ : Odrv4
    port map (
            O => \N__42848\,
            I => n13415
        );

    \I__10050\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42833\
        );

    \I__10049\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42830\
        );

    \I__10048\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42824\
        );

    \I__10047\ : InMux
    port map (
            O => \N__42836\,
            I => \N__42821\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__42833\,
            I => \N__42818\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__42830\,
            I => \N__42815\
        );

    \I__10044\ : InMux
    port map (
            O => \N__42829\,
            I => \N__42808\
        );

    \I__10043\ : InMux
    port map (
            O => \N__42828\,
            I => \N__42808\
        );

    \I__10042\ : InMux
    port map (
            O => \N__42827\,
            I => \N__42808\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__42824\,
            I => \tx_transmit_N_2239_3\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__42821\,
            I => \tx_transmit_N_2239_3\
        );

    \I__10039\ : Odrv12
    port map (
            O => \N__42818\,
            I => \tx_transmit_N_2239_3\
        );

    \I__10038\ : Odrv4
    port map (
            O => \N__42815\,
            I => \tx_transmit_N_2239_3\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__42808\,
            I => \tx_transmit_N_2239_3\
        );

    \I__10036\ : CascadeMux
    port map (
            O => \N__42797\,
            I => \N__42794\
        );

    \I__10035\ : InMux
    port map (
            O => \N__42794\,
            I => \N__42790\
        );

    \I__10034\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42787\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__42790\,
            I => \N__42784\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__42787\,
            I => \r_Tx_Data_5\
        );

    \I__10031\ : Odrv12
    port map (
            O => \N__42784\,
            I => \r_Tx_Data_5\
        );

    \I__10030\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42775\
        );

    \I__10029\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42772\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__42775\,
            I => \N__42769\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__42772\,
            I => n16485
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__42769\,
            I => n16485
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__42764\,
            I => \N__42761\
        );

    \I__10024\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42758\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42755\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__42755\,
            I => \N__42752\
        );

    \I__10021\ : Odrv4
    port map (
            O => \N__42752\,
            I => \c0.n7428\
        );

    \I__10020\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42746\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__42746\,
            I => \N__42741\
        );

    \I__10018\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42736\
        );

    \I__10017\ : InMux
    port map (
            O => \N__42744\,
            I => \N__42736\
        );

    \I__10016\ : Sp12to4
    port map (
            O => \N__42741\,
            I => \N__42731\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__42736\,
            I => \N__42731\
        );

    \I__10014\ : Span12Mux_s7_v
    port map (
            O => \N__42731\,
            I => \N__42726\
        );

    \I__10013\ : InMux
    port map (
            O => \N__42730\,
            I => \N__42723\
        );

    \I__10012\ : InMux
    port map (
            O => \N__42729\,
            I => \N__42720\
        );

    \I__10011\ : Odrv12
    port map (
            O => \N__42726\,
            I => n14_adj_2615
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__42723\,
            I => n14_adj_2615
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__42720\,
            I => n14_adj_2615
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__42713\,
            I => \N__42709\
        );

    \I__10007\ : InMux
    port map (
            O => \N__42712\,
            I => \N__42701\
        );

    \I__10006\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42701\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__42708\,
            I => \N__42698\
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__42707\,
            I => \N__42693\
        );

    \I__10003\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42689\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__42701\,
            I => \N__42686\
        );

    \I__10001\ : InMux
    port map (
            O => \N__42698\,
            I => \N__42683\
        );

    \I__10000\ : InMux
    port map (
            O => \N__42697\,
            I => \N__42678\
        );

    \I__9999\ : InMux
    port map (
            O => \N__42696\,
            I => \N__42678\
        );

    \I__9998\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42675\
        );

    \I__9997\ : CascadeMux
    port map (
            O => \N__42692\,
            I => \N__42672\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__42689\,
            I => \N__42669\
        );

    \I__9995\ : Span4Mux_h
    port map (
            O => \N__42686\,
            I => \N__42660\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__42683\,
            I => \N__42660\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__42678\,
            I => \N__42660\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__42675\,
            I => \N__42660\
        );

    \I__9991\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42657\
        );

    \I__9990\ : Span4Mux_v
    port map (
            O => \N__42669\,
            I => \N__42653\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__42660\,
            I => \N__42650\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42647\
        );

    \I__9987\ : InMux
    port map (
            O => \N__42656\,
            I => \N__42644\
        );

    \I__9986\ : Odrv4
    port map (
            O => \N__42653\,
            I => n9631
        );

    \I__9985\ : Odrv4
    port map (
            O => \N__42650\,
            I => n9631
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__42647\,
            I => n9631
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__42644\,
            I => n9631
        );

    \I__9982\ : CascadeMux
    port map (
            O => \N__42635\,
            I => \N__42632\
        );

    \I__9981\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42629\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42625\
        );

    \I__9979\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42622\
        );

    \I__9978\ : Odrv4
    port map (
            O => \N__42625\,
            I => \tx_transmit_N_2239_6\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__42622\,
            I => \tx_transmit_N_2239_6\
        );

    \I__9976\ : CascadeMux
    port map (
            O => \N__42617\,
            I => \N__42613\
        );

    \I__9975\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9974\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__42610\,
            I => byte_transmit_counter_6
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__42607\,
            I => byte_transmit_counter_6
        );

    \I__9971\ : InMux
    port map (
            O => \N__42602\,
            I => \N__42598\
        );

    \I__9970\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42595\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__42598\,
            I => \c0.n149\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__42595\,
            I => \c0.n149\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__42590\,
            I => \N__42587\
        );

    \I__9966\ : InMux
    port map (
            O => \N__42587\,
            I => \N__42584\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__42584\,
            I => \c0.n17741\
        );

    \I__9964\ : CascadeMux
    port map (
            O => \N__42581\,
            I => \N__42576\
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__42580\,
            I => \N__42563\
        );

    \I__9962\ : InMux
    port map (
            O => \N__42579\,
            I => \N__42556\
        );

    \I__9961\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42556\
        );

    \I__9960\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42546\
        );

    \I__9959\ : InMux
    port map (
            O => \N__42574\,
            I => \N__42546\
        );

    \I__9958\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42541\
        );

    \I__9957\ : InMux
    port map (
            O => \N__42572\,
            I => \N__42541\
        );

    \I__9956\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42538\
        );

    \I__9955\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42535\
        );

    \I__9954\ : InMux
    port map (
            O => \N__42569\,
            I => \N__42532\
        );

    \I__9953\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42529\
        );

    \I__9952\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42526\
        );

    \I__9951\ : InMux
    port map (
            O => \N__42566\,
            I => \N__42521\
        );

    \I__9950\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42521\
        );

    \I__9949\ : InMux
    port map (
            O => \N__42562\,
            I => \N__42516\
        );

    \I__9948\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42516\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__42556\,
            I => \N__42513\
        );

    \I__9946\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42510\
        );

    \I__9945\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42507\
        );

    \I__9944\ : InMux
    port map (
            O => \N__42553\,
            I => \N__42504\
        );

    \I__9943\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42499\
        );

    \I__9942\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42499\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__42546\,
            I => \N__42496\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__42541\,
            I => \N__42493\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__42538\,
            I => \N__42488\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__42535\,
            I => \N__42488\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__42532\,
            I => n29
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__42529\,
            I => n29
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__42526\,
            I => n29
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__42521\,
            I => n29
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__42516\,
            I => n29
        );

    \I__9932\ : Odrv4
    port map (
            O => \N__42513\,
            I => n29
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__42510\,
            I => n29
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__42507\,
            I => n29
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__42504\,
            I => n29
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__42499\,
            I => n29
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__42496\,
            I => n29
        );

    \I__9926\ : Odrv4
    port map (
            O => \N__42493\,
            I => n29
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__42488\,
            I => n29
        );

    \I__9924\ : CascadeMux
    port map (
            O => \N__42461\,
            I => \N__42458\
        );

    \I__9923\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42455\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__42455\,
            I => \N__42452\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__42452\,
            I => \c0.n7268\
        );

    \I__9920\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42445\
        );

    \I__9919\ : InMux
    port map (
            O => \N__42448\,
            I => \N__42442\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__42445\,
            I => \N__42439\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__42442\,
            I => \N__42424\
        );

    \I__9916\ : Span4Mux_h
    port map (
            O => \N__42439\,
            I => \N__42421\
        );

    \I__9915\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42416\
        );

    \I__9914\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42416\
        );

    \I__9913\ : InMux
    port map (
            O => \N__42436\,
            I => \N__42407\
        );

    \I__9912\ : InMux
    port map (
            O => \N__42435\,
            I => \N__42407\
        );

    \I__9911\ : InMux
    port map (
            O => \N__42434\,
            I => \N__42407\
        );

    \I__9910\ : InMux
    port map (
            O => \N__42433\,
            I => \N__42407\
        );

    \I__9909\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42400\
        );

    \I__9908\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42400\
        );

    \I__9907\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42400\
        );

    \I__9906\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42393\
        );

    \I__9905\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42393\
        );

    \I__9904\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42393\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__42424\,
            I => \c0.n1314\
        );

    \I__9902\ : Odrv4
    port map (
            O => \N__42421\,
            I => \c0.n1314\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__42416\,
            I => \c0.n1314\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__42407\,
            I => \c0.n1314\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__42400\,
            I => \c0.n1314\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__42393\,
            I => \c0.n1314\
        );

    \I__9897\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42376\
        );

    \I__9896\ : InMux
    port map (
            O => \N__42379\,
            I => \N__42371\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__42376\,
            I => \N__42368\
        );

    \I__9894\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42363\
        );

    \I__9893\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42363\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__42371\,
            I => \c0.delay_counter_7\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__42368\,
            I => \c0.delay_counter_7\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__42363\,
            I => \c0.delay_counter_7\
        );

    \I__9889\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42350\
        );

    \I__9888\ : InMux
    port map (
            O => \N__42355\,
            I => \N__42347\
        );

    \I__9887\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42342\
        );

    \I__9886\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42342\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__42350\,
            I => \c0.delay_counter_11\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__42347\,
            I => \c0.delay_counter_11\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__42342\,
            I => \c0.delay_counter_11\
        );

    \I__9882\ : InMux
    port map (
            O => \N__42335\,
            I => \N__42330\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__42334\,
            I => \N__42326\
        );

    \I__9880\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42323\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__42330\,
            I => \N__42320\
        );

    \I__9878\ : InMux
    port map (
            O => \N__42329\,
            I => \N__42315\
        );

    \I__9877\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42315\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__42323\,
            I => \N__42312\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__42320\,
            I => \N__42309\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__42315\,
            I => \c0.delay_counter_8\
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__42312\,
            I => \c0.delay_counter_8\
        );

    \I__9872\ : Odrv4
    port map (
            O => \N__42309\,
            I => \c0.delay_counter_8\
        );

    \I__9871\ : CascadeMux
    port map (
            O => \N__42302\,
            I => \N__42297\
        );

    \I__9870\ : InMux
    port map (
            O => \N__42301\,
            I => \N__42293\
        );

    \I__9869\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42290\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42287\
        );

    \I__9867\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42284\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__42293\,
            I => \c0.delay_counter_5\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__42290\,
            I => \c0.delay_counter_5\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__42287\,
            I => \c0.delay_counter_5\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__42284\,
            I => \c0.delay_counter_5\
        );

    \I__9862\ : CascadeMux
    port map (
            O => \N__42275\,
            I => \c0.n10_adj_2532_cascade_\
        );

    \I__9861\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42269\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__42269\,
            I => \N__42266\
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__42266\,
            I => \c0.n14_adj_2533\
        );

    \I__9858\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42260\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__42260\,
            I => \N__42257\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__42257\,
            I => \N__42254\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__42254\,
            I => n17306
        );

    \I__9854\ : CascadeMux
    port map (
            O => \N__42251\,
            I => \n17306_cascade_\
        );

    \I__9853\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42245\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__42245\,
            I => \N__42242\
        );

    \I__9851\ : Span12Mux_s4_v
    port map (
            O => \N__42242\,
            I => \N__42237\
        );

    \I__9850\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42234\
        );

    \I__9849\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42231\
        );

    \I__9848\ : Odrv12
    port map (
            O => \N__42237\,
            I => \c0.n17387\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__42234\,
            I => \c0.n17387\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__42231\,
            I => \c0.n17387\
        );

    \I__9845\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42221\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__42221\,
            I => \c0.n6_adj_2534\
        );

    \I__9843\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42215\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__42215\,
            I => \N__42212\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__42212\,
            I => \N__42209\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__42209\,
            I => \tx_data_4_N_keep\
        );

    \I__9839\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42202\
        );

    \I__9838\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42199\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__42202\,
            I => \N__42196\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__42199\,
            I => \r_Tx_Data_4\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__42196\,
            I => \r_Tx_Data_4\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__42191\,
            I => \c0.n16_adj_2445_cascade_\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__42188\,
            I => \c0.n19_adj_2446_cascade_\
        );

    \I__9832\ : InMux
    port map (
            O => \N__42185\,
            I => \N__42180\
        );

    \I__9831\ : InMux
    port map (
            O => \N__42184\,
            I => \N__42177\
        );

    \I__9830\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42172\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__42180\,
            I => \N__42167\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__42177\,
            I => \N__42167\
        );

    \I__9827\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42162\
        );

    \I__9826\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42162\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__42172\,
            I => \c0.n8550\
        );

    \I__9824\ : Odrv4
    port map (
            O => \N__42167\,
            I => \c0.n8550\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__42162\,
            I => \c0.n8550\
        );

    \I__9822\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42151\
        );

    \I__9821\ : InMux
    port map (
            O => \N__42154\,
            I => \N__42148\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__42151\,
            I => n96
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__42148\,
            I => n96
        );

    \I__9818\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42139\
        );

    \I__9817\ : InMux
    port map (
            O => \N__42142\,
            I => \N__42136\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__42139\,
            I => n6878
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__42136\,
            I => n6878
        );

    \I__9814\ : CascadeMux
    port map (
            O => \N__42131\,
            I => \n17672_cascade_\
        );

    \I__9813\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42123\
        );

    \I__9812\ : InMux
    port map (
            O => \N__42127\,
            I => \N__42120\
        );

    \I__9811\ : InMux
    port map (
            O => \N__42126\,
            I => \N__42117\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__42123\,
            I => \c0.n113\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__42120\,
            I => \c0.n113\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__42117\,
            I => \c0.n113\
        );

    \I__9807\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42103\
        );

    \I__9806\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42103\
        );

    \I__9805\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42100\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__42103\,
            I => n17364
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__42100\,
            I => n17364
        );

    \I__9802\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42092\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__42092\,
            I => \N__42089\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__42089\,
            I => \N__42086\
        );

    \I__9799\ : Odrv4
    port map (
            O => \N__42086\,
            I => \c0.n18009\
        );

    \I__9798\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42078\
        );

    \I__9797\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42075\
        );

    \I__9796\ : InMux
    port map (
            O => \N__42081\,
            I => \N__42072\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__42078\,
            I => \N__42069\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__42075\,
            I => \N__42066\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__42072\,
            I => \N__42058\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__42069\,
            I => \N__42058\
        );

    \I__9791\ : Span4Mux_v
    port map (
            O => \N__42066\,
            I => \N__42058\
        );

    \I__9790\ : InMux
    port map (
            O => \N__42065\,
            I => \N__42055\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__42058\,
            I => \c0.delay_counter_12\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__42055\,
            I => \c0.delay_counter_12\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42050\,
            I => \N__42044\
        );

    \I__9786\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42041\
        );

    \I__9785\ : InMux
    port map (
            O => \N__42048\,
            I => \N__42038\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42047\,
            I => \N__42035\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__42044\,
            I => \N__42032\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__42041\,
            I => \N__42029\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__42038\,
            I => \N__42026\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__42035\,
            I => \N__42023\
        );

    \I__9779\ : Odrv12
    port map (
            O => \N__42032\,
            I => n119
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__42029\,
            I => n119
        );

    \I__9777\ : Odrv4
    port map (
            O => \N__42026\,
            I => n119
        );

    \I__9776\ : Odrv12
    port map (
            O => \N__42023\,
            I => n119
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__42014\,
            I => \UART_TRANSMITTER_state_7_N_1749_2_cascade_\
        );

    \I__9774\ : InMux
    port map (
            O => \N__42011\,
            I => \N__42008\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__42008\,
            I => n18032
        );

    \I__9772\ : InMux
    port map (
            O => \N__42005\,
            I => \N__42000\
        );

    \I__9771\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41995\
        );

    \I__9770\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41995\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__42000\,
            I => n8488
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__41995\,
            I => n8488
        );

    \I__9767\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41985\
        );

    \I__9766\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41980\
        );

    \I__9765\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41980\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__41985\,
            I => n17709
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__41980\,
            I => n17709
        );

    \I__9762\ : CascadeMux
    port map (
            O => \N__41975\,
            I => \N__41971\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__41974\,
            I => \N__41968\
        );

    \I__9760\ : InMux
    port map (
            O => \N__41971\,
            I => \N__41965\
        );

    \I__9759\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41961\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__41965\,
            I => \N__41957\
        );

    \I__9757\ : InMux
    port map (
            O => \N__41964\,
            I => \N__41954\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41951\
        );

    \I__9755\ : InMux
    port map (
            O => \N__41960\,
            I => \N__41948\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__41957\,
            I => \N__41945\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__41954\,
            I => \c0.delay_counter_6\
        );

    \I__9752\ : Odrv12
    port map (
            O => \N__41951\,
            I => \c0.delay_counter_6\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__41948\,
            I => \c0.delay_counter_6\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__41945\,
            I => \c0.delay_counter_6\
        );

    \I__9749\ : CascadeMux
    port map (
            O => \N__41936\,
            I => \N__41932\
        );

    \I__9748\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41928\
        );

    \I__9747\ : InMux
    port map (
            O => \N__41932\,
            I => \N__41924\
        );

    \I__9746\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41921\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41918\
        );

    \I__9744\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41915\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__41924\,
            I => \N__41910\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__41921\,
            I => \N__41910\
        );

    \I__9741\ : Span4Mux_h
    port map (
            O => \N__41918\,
            I => \N__41907\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__41915\,
            I => \c0.delay_counter_9\
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__41910\,
            I => \c0.delay_counter_9\
        );

    \I__9738\ : Odrv4
    port map (
            O => \N__41907\,
            I => \c0.delay_counter_9\
        );

    \I__9737\ : InMux
    port map (
            O => \N__41900\,
            I => \N__41897\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__41897\,
            I => \N__41894\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9734\ : Odrv4
    port map (
            O => \N__41891\,
            I => \c0.n17753\
        );

    \I__9733\ : CascadeMux
    port map (
            O => \N__41888\,
            I => \c0.n17662_cascade_\
        );

    \I__9732\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__41882\,
            I => \N__41878\
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__41881\,
            I => \N__41875\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__41878\,
            I => \N__41872\
        );

    \I__9728\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41869\
        );

    \I__9727\ : Odrv4
    port map (
            O => \N__41872\,
            I => rand_setpoint_23
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__41869\,
            I => rand_setpoint_23
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__41864\,
            I => \c0.n2041_cascade_\
        );

    \I__9724\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41858\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41855\
        );

    \I__9722\ : Span4Mux_s2_v
    port map (
            O => \N__41855\,
            I => \N__41852\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__41852\,
            I => \c0.n17974\
        );

    \I__9720\ : InMux
    port map (
            O => \N__41849\,
            I => \N__41846\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__41846\,
            I => \N__41842\
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__41845\,
            I => \N__41839\
        );

    \I__9717\ : Span4Mux_s1_v
    port map (
            O => \N__41842\,
            I => \N__41836\
        );

    \I__9716\ : InMux
    port map (
            O => \N__41839\,
            I => \N__41833\
        );

    \I__9715\ : Odrv4
    port map (
            O => \N__41836\,
            I => rand_setpoint_16
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__41833\,
            I => rand_setpoint_16
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__41828\,
            I => \c0.n17693_cascade_\
        );

    \I__9712\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41822\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__41822\,
            I => \N__41818\
        );

    \I__9710\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41815\
        );

    \I__9709\ : Span4Mux_h
    port map (
            O => \N__41818\,
            I => \N__41810\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__41815\,
            I => \N__41810\
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__41810\,
            I => \c0.data_out_6_0\
        );

    \I__9706\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41804\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__41804\,
            I => \N__41801\
        );

    \I__9704\ : Span4Mux_v
    port map (
            O => \N__41801\,
            I => \N__41798\
        );

    \I__9703\ : Span4Mux_h
    port map (
            O => \N__41798\,
            I => \N__41794\
        );

    \I__9702\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41789\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__41794\,
            I => \N__41786\
        );

    \I__9700\ : CascadeMux
    port map (
            O => \N__41793\,
            I => \N__41783\
        );

    \I__9699\ : InMux
    port map (
            O => \N__41792\,
            I => \N__41780\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__41789\,
            I => \N__41775\
        );

    \I__9697\ : Sp12to4
    port map (
            O => \N__41786\,
            I => \N__41775\
        );

    \I__9696\ : InMux
    port map (
            O => \N__41783\,
            I => \N__41772\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__41780\,
            I => \N__41769\
        );

    \I__9694\ : Span12Mux_v
    port map (
            O => \N__41775\,
            I => \N__41766\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__41772\,
            I => data_out_1_7
        );

    \I__9692\ : Odrv4
    port map (
            O => \N__41769\,
            I => data_out_1_7
        );

    \I__9691\ : Odrv12
    port map (
            O => \N__41766\,
            I => data_out_1_7
        );

    \I__9690\ : InMux
    port map (
            O => \N__41759\,
            I => \N__41756\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__41756\,
            I => \N__41752\
        );

    \I__9688\ : InMux
    port map (
            O => \N__41755\,
            I => \N__41749\
        );

    \I__9687\ : Odrv12
    port map (
            O => \N__41752\,
            I => \c0.n17578\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__41749\,
            I => \c0.n17578\
        );

    \I__9685\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41740\
        );

    \I__9684\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41735\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41732\
        );

    \I__9682\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41727\
        );

    \I__9681\ : InMux
    port map (
            O => \N__41738\,
            I => \N__41727\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__41735\,
            I => \N__41722\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__41732\,
            I => \N__41722\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__41727\,
            I => \c0.delay_counter_10\
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__41722\,
            I => \c0.delay_counter_10\
        );

    \I__9676\ : InMux
    port map (
            O => \N__41717\,
            I => \N__41713\
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__41716\,
            I => \N__41710\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__41713\,
            I => \N__41707\
        );

    \I__9673\ : InMux
    port map (
            O => \N__41710\,
            I => \N__41704\
        );

    \I__9672\ : Odrv12
    port map (
            O => \N__41707\,
            I => rand_setpoint_12
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__41704\,
            I => rand_setpoint_12
        );

    \I__9670\ : CascadeMux
    port map (
            O => \N__41699\,
            I => \c0.n17931_cascade_\
        );

    \I__9669\ : CascadeMux
    port map (
            O => \N__41696\,
            I => \N__41693\
        );

    \I__9668\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41690\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__41690\,
            I => \N__41686\
        );

    \I__9666\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41683\
        );

    \I__9665\ : Span4Mux_h
    port map (
            O => \N__41686\,
            I => \N__41678\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__41683\,
            I => \N__41678\
        );

    \I__9663\ : Span4Mux_s2_v
    port map (
            O => \N__41678\,
            I => \N__41675\
        );

    \I__9662\ : Odrv4
    port map (
            O => \N__41675\,
            I => \c0.n17400\
        );

    \I__9661\ : InMux
    port map (
            O => \N__41672\,
            I => \N__41669\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__41669\,
            I => \N__41665\
        );

    \I__9659\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41662\
        );

    \I__9658\ : Odrv12
    port map (
            O => \N__41665\,
            I => \c0.data_out_7__4__N_550\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__41662\,
            I => \c0.data_out_7__4__N_550\
        );

    \I__9656\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41653\
        );

    \I__9655\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41650\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__41653\,
            I => \N__41645\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__41650\,
            I => \N__41642\
        );

    \I__9652\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41637\
        );

    \I__9651\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41637\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__41645\,
            I => \N__41634\
        );

    \I__9649\ : Span4Mux_h
    port map (
            O => \N__41642\,
            I => \N__41631\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__41637\,
            I => \c0.data_out_7_4\
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__41634\,
            I => \c0.data_out_7_4\
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__41631\,
            I => \c0.data_out_7_4\
        );

    \I__9645\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41616\
        );

    \I__9644\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41616\
        );

    \I__9643\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41611\
        );

    \I__9642\ : InMux
    port map (
            O => \N__41621\,
            I => \N__41608\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__41616\,
            I => \N__41605\
        );

    \I__9640\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41600\
        );

    \I__9639\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41600\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__41611\,
            I => \data_out_5__4__N_959\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__41608\,
            I => \data_out_5__4__N_959\
        );

    \I__9636\ : Odrv4
    port map (
            O => \N__41605\,
            I => \data_out_5__4__N_959\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__41600\,
            I => \data_out_5__4__N_959\
        );

    \I__9634\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41588\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__41588\,
            I => \N__41584\
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__41587\,
            I => \N__41581\
        );

    \I__9631\ : Span4Mux_h
    port map (
            O => \N__41584\,
            I => \N__41578\
        );

    \I__9630\ : InMux
    port map (
            O => \N__41581\,
            I => \N__41575\
        );

    \I__9629\ : Odrv4
    port map (
            O => \N__41578\,
            I => rand_setpoint_28
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__41575\,
            I => rand_setpoint_28
        );

    \I__9627\ : CascadeMux
    port map (
            O => \N__41570\,
            I => \c0.n17967_cascade_\
        );

    \I__9626\ : CascadeMux
    port map (
            O => \N__41567\,
            I => \N__41564\
        );

    \I__9625\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41561\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__41561\,
            I => \N__41558\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__41558\,
            I => \c0.n6_adj_2467\
        );

    \I__9622\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41552\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__41552\,
            I => \N__41549\
        );

    \I__9620\ : Odrv4
    port map (
            O => \N__41549\,
            I => \c0.n9276\
        );

    \I__9619\ : CascadeMux
    port map (
            O => \N__41546\,
            I => \N__41542\
        );

    \I__9618\ : InMux
    port map (
            O => \N__41545\,
            I => \N__41538\
        );

    \I__9617\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41535\
        );

    \I__9616\ : InMux
    port map (
            O => \N__41541\,
            I => \N__41532\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__41538\,
            I => \c0.n8634\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__41535\,
            I => \c0.n8634\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__41532\,
            I => \c0.n8634\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__41525\,
            I => \c0.n9276_cascade_\
        );

    \I__9611\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41519\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__41519\,
            I => \N__41516\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__41516\,
            I => \N__41513\
        );

    \I__9608\ : Odrv4
    port map (
            O => \N__41513\,
            I => \c0.data_out_7__1__N_626\
        );

    \I__9607\ : CascadeMux
    port map (
            O => \N__41510\,
            I => \c0.n17623_cascade_\
        );

    \I__9606\ : InMux
    port map (
            O => \N__41507\,
            I => \N__41504\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__41504\,
            I => \N__41501\
        );

    \I__9604\ : Span4Mux_v
    port map (
            O => \N__41501\,
            I => \N__41497\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__41500\,
            I => \N__41494\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__41497\,
            I => \N__41491\
        );

    \I__9601\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41488\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__41491\,
            I => rand_setpoint_8
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__41488\,
            I => rand_setpoint_8
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__41483\,
            I => \c0.n17916_cascade_\
        );

    \I__9597\ : InMux
    port map (
            O => \N__41480\,
            I => \N__41477\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__41477\,
            I => \N__41473\
        );

    \I__9595\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41470\
        );

    \I__9594\ : Span4Mux_h
    port map (
            O => \N__41473\,
            I => \N__41467\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__41470\,
            I => \N__41464\
        );

    \I__9592\ : Span4Mux_v
    port map (
            O => \N__41467\,
            I => \N__41461\
        );

    \I__9591\ : Span4Mux_h
    port map (
            O => \N__41464\,
            I => \N__41458\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__41461\,
            I => \c0.data_out_7_0\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__41458\,
            I => \c0.data_out_7_0\
        );

    \I__9588\ : CascadeMux
    port map (
            O => \N__41453\,
            I => \N__41450\
        );

    \I__9587\ : InMux
    port map (
            O => \N__41450\,
            I => \N__41447\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__41447\,
            I => \N__41444\
        );

    \I__9585\ : Span4Mux_v
    port map (
            O => \N__41444\,
            I => \N__41441\
        );

    \I__9584\ : Span4Mux_v
    port map (
            O => \N__41441\,
            I => \N__41438\
        );

    \I__9583\ : Odrv4
    port map (
            O => \N__41438\,
            I => \c0.n8486\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__41435\,
            I => \c0.n8486_cascade_\
        );

    \I__9581\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41429\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41426\
        );

    \I__9579\ : Odrv12
    port map (
            O => \N__41426\,
            I => \c0.n16450\
        );

    \I__9578\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41420\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41417\
        );

    \I__9576\ : Span4Mux_v
    port map (
            O => \N__41417\,
            I => \N__41414\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__41414\,
            I => n4_adj_2612
        );

    \I__9574\ : InMux
    port map (
            O => \N__41411\,
            I => \N__41407\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__41410\,
            I => \N__41404\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__41407\,
            I => \N__41401\
        );

    \I__9571\ : InMux
    port map (
            O => \N__41404\,
            I => \N__41398\
        );

    \I__9570\ : Odrv12
    port map (
            O => \N__41401\,
            I => rand_setpoint_13
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__41398\,
            I => rand_setpoint_13
        );

    \I__9568\ : CascadeMux
    port map (
            O => \N__41393\,
            I => \c0.n17925_cascade_\
        );

    \I__9567\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41387\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__41387\,
            I => \c0.n18068\
        );

    \I__9565\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41381\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__41381\,
            I => \c0.n5_adj_2490\
        );

    \I__9563\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41375\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__41375\,
            I => \c0.data_out_10_4\
        );

    \I__9561\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41369\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__41369\,
            I => \c0.n18067\
        );

    \I__9559\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41363\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__41363\,
            I => \c0.n18092\
        );

    \I__9557\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41357\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__41354\,
            I => \c0.n18094\
        );

    \I__9554\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41348\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__41348\,
            I => \N__41345\
        );

    \I__9552\ : Span4Mux_h
    port map (
            O => \N__41345\,
            I => \N__41342\
        );

    \I__9551\ : Span4Mux_v
    port map (
            O => \N__41342\,
            I => \N__41339\
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__41339\,
            I => \c0.n18096\
        );

    \I__9549\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__9547\ : Span4Mux_h
    port map (
            O => \N__41330\,
            I => \N__41327\
        );

    \I__9546\ : Odrv4
    port map (
            O => \N__41327\,
            I => \c0.n18088\
        );

    \I__9545\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41317\
        );

    \I__9543\ : InMux
    port map (
            O => \N__41320\,
            I => \N__41314\
        );

    \I__9542\ : Span4Mux_h
    port map (
            O => \N__41317\,
            I => \N__41311\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__41314\,
            I => byte_transmit_counter_5
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__41311\,
            I => byte_transmit_counter_5
        );

    \I__9539\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41303\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__41303\,
            I => \N__41300\
        );

    \I__9537\ : Span4Mux_h
    port map (
            O => \N__41300\,
            I => \N__41296\
        );

    \I__9536\ : InMux
    port map (
            O => \N__41299\,
            I => \N__41293\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__41296\,
            I => \tx_transmit_N_2239_5\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41293\,
            I => \tx_transmit_N_2239_5\
        );

    \I__9533\ : InMux
    port map (
            O => \N__41288\,
            I => \c0.n16354\
        );

    \I__9532\ : InMux
    port map (
            O => \N__41285\,
            I => \c0.n16355\
        );

    \I__9531\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41278\
        );

    \I__9530\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41275\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__41278\,
            I => byte_transmit_counter_7
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__41275\,
            I => byte_transmit_counter_7
        );

    \I__9527\ : InMux
    port map (
            O => \N__41270\,
            I => \c0.n16356\
        );

    \I__9526\ : InMux
    port map (
            O => \N__41267\,
            I => \N__41263\
        );

    \I__9525\ : InMux
    port map (
            O => \N__41266\,
            I => \N__41260\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__41263\,
            I => \tx_transmit_N_2239_7\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__41260\,
            I => \tx_transmit_N_2239_7\
        );

    \I__9522\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41251\
        );

    \I__9521\ : CascadeMux
    port map (
            O => \N__41254\,
            I => \N__41248\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__41251\,
            I => \N__41245\
        );

    \I__9519\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41241\
        );

    \I__9518\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41238\
        );

    \I__9517\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41234\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__41241\,
            I => \N__41231\
        );

    \I__9515\ : Span4Mux_v
    port map (
            O => \N__41238\,
            I => \N__41228\
        );

    \I__9514\ : InMux
    port map (
            O => \N__41237\,
            I => \N__41225\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__41234\,
            I => data_out_3_4
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__41231\,
            I => data_out_3_4
        );

    \I__9511\ : Odrv4
    port map (
            O => \N__41228\,
            I => data_out_3_4
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__41225\,
            I => data_out_3_4
        );

    \I__9509\ : CascadeMux
    port map (
            O => \N__41216\,
            I => \c0.n18093_cascade_\
        );

    \I__9508\ : CascadeMux
    port map (
            O => \N__41213\,
            I => \c0.n18399_cascade_\
        );

    \I__9507\ : CascadeMux
    port map (
            O => \N__41210\,
            I => \N__41206\
        );

    \I__9506\ : InMux
    port map (
            O => \N__41209\,
            I => \N__41203\
        );

    \I__9505\ : InMux
    port map (
            O => \N__41206\,
            I => \N__41200\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__41203\,
            I => \tx_transmit_N_2239_4\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__41200\,
            I => \tx_transmit_N_2239_4\
        );

    \I__9502\ : InMux
    port map (
            O => \N__41195\,
            I => \N__41192\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__41192\,
            I => \c0.n5_adj_2447\
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__41189\,
            I => \c0.n17941_cascade_\
        );

    \I__9499\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__41183\,
            I => \c0.n18396\
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__41180\,
            I => \n8529_cascade_\
        );

    \I__9496\ : CascadeMux
    port map (
            O => \N__41177\,
            I => \c0.n8550_cascade_\
        );

    \I__9495\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__41171\,
            I => n121_adj_2606
        );

    \I__9493\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41165\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__41165\,
            I => n8529
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__41162\,
            I => \n121_adj_2606_cascade_\
        );

    \I__9490\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41156\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__41156\,
            I => \N__41153\
        );

    \I__9488\ : Odrv4
    port map (
            O => \N__41153\,
            I => n13_adj_2652
        );

    \I__9487\ : InMux
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__41147\,
            I => \c0.n251\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41144\,
            I => \c0.n16350\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41141\,
            I => \c0.n16351\
        );

    \I__9483\ : InMux
    port map (
            O => \N__41138\,
            I => \c0.n16352\
        );

    \I__9482\ : InMux
    port map (
            O => \N__41135\,
            I => \c0.n16353\
        );

    \I__9481\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41129\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__41126\,
            I => \c0.n18008\
        );

    \I__9478\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41118\
        );

    \I__9477\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41115\
        );

    \I__9476\ : InMux
    port map (
            O => \N__41121\,
            I => \N__41112\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__41118\,
            I => \N__41107\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41107\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__41112\,
            I => \c0.delay_counter_3\
        );

    \I__9472\ : Odrv4
    port map (
            O => \N__41107\,
            I => \c0.delay_counter_3\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41097\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41092\
        );

    \I__9469\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41092\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__41097\,
            I => \c0.delay_counter_1\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__41092\,
            I => \c0.delay_counter_1\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__41087\,
            I => \N__41082\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41086\,
            I => \N__41079\
        );

    \I__9464\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41076\
        );

    \I__9463\ : InMux
    port map (
            O => \N__41082\,
            I => \N__41073\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__41079\,
            I => \c0.delay_counter_2\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__41076\,
            I => \c0.delay_counter_2\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__41073\,
            I => \c0.delay_counter_2\
        );

    \I__9459\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41061\
        );

    \I__9458\ : InMux
    port map (
            O => \N__41065\,
            I => \N__41058\
        );

    \I__9457\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41055\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__41061\,
            I => \c0.delay_counter_4\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__41058\,
            I => \c0.delay_counter_4\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__41055\,
            I => \c0.delay_counter_4\
        );

    \I__9453\ : InMux
    port map (
            O => \N__41048\,
            I => \N__41044\
        );

    \I__9452\ : InMux
    port map (
            O => \N__41047\,
            I => \N__41040\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__41044\,
            I => \N__41037\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41043\,
            I => \N__41033\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__41040\,
            I => \N__41028\
        );

    \I__9448\ : Span4Mux_v
    port map (
            O => \N__41037\,
            I => \N__41028\
        );

    \I__9447\ : InMux
    port map (
            O => \N__41036\,
            I => \N__41025\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__41033\,
            I => delay_counter_0
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__41028\,
            I => delay_counter_0
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41025\,
            I => delay_counter_0
        );

    \I__9443\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41012\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__41012\,
            I => \N__41006\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__41011\,
            I => \N__41003\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__41010\,
            I => \N__41000\
        );

    \I__9438\ : InMux
    port map (
            O => \N__41009\,
            I => \N__40997\
        );

    \I__9437\ : Sp12to4
    port map (
            O => \N__41006\,
            I => \N__40994\
        );

    \I__9436\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40989\
        );

    \I__9435\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40989\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__40997\,
            I => delay_counter_13
        );

    \I__9433\ : Odrv12
    port map (
            O => \N__40994\,
            I => delay_counter_13
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__40989\,
            I => delay_counter_13
        );

    \I__9431\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40978\
        );

    \I__9430\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40975\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__40978\,
            I => \N__40969\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__40975\,
            I => \N__40969\
        );

    \I__9427\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40965\
        );

    \I__9426\ : Span4Mux_v
    port map (
            O => \N__40969\,
            I => \N__40962\
        );

    \I__9425\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40959\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__40965\,
            I => delay_counter_14
        );

    \I__9423\ : Odrv4
    port map (
            O => \N__40962\,
            I => delay_counter_14
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__40959\,
            I => delay_counter_14
        );

    \I__9421\ : InMux
    port map (
            O => \N__40952\,
            I => \N__40949\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__40949\,
            I => \c0.n7264\
        );

    \I__9419\ : CascadeMux
    port map (
            O => \N__40946\,
            I => \n29_cascade_\
        );

    \I__9418\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40939\
        );

    \I__9417\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40936\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__40939\,
            I => data_in_12_6
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__40936\,
            I => data_in_12_6
        );

    \I__9414\ : CascadeMux
    port map (
            O => \N__40931\,
            I => \c0.n149_cascade_\
        );

    \I__9413\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40925\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__40925\,
            I => \N__40922\
        );

    \I__9411\ : Span4Mux_h
    port map (
            O => \N__40922\,
            I => \N__40919\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__40919\,
            I => \c0.n93\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__40916\,
            I => \N__40913\
        );

    \I__9408\ : InMux
    port map (
            O => \N__40913\,
            I => \N__40910\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__40910\,
            I => n17958
        );

    \I__9406\ : InMux
    port map (
            O => \N__40907\,
            I => \N__40904\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__40904\,
            I => n43
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__40901\,
            I => \N__40898\
        );

    \I__9403\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40895\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__40895\,
            I => \c0.n7271\
        );

    \I__9401\ : CascadeMux
    port map (
            O => \N__40892\,
            I => \N__40889\
        );

    \I__9400\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40886\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__40886\,
            I => \N__40883\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__40883\,
            I => \c0.n18105\
        );

    \I__9397\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40877\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__40877\,
            I => \c0.n18012\
        );

    \I__9395\ : InMux
    port map (
            O => \N__40874\,
            I => \N__40871\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__40871\,
            I => \N__40868\
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__40868\,
            I => \c0.n17936\
        );

    \I__9392\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40862\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__40862\,
            I => \c0.n7275\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__40859\,
            I => \N__40856\
        );

    \I__9389\ : InMux
    port map (
            O => \N__40856\,
            I => \N__40853\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__40853\,
            I => \c0.n7274\
        );

    \I__9387\ : InMux
    port map (
            O => \N__40850\,
            I => \N__40843\
        );

    \I__9386\ : InMux
    port map (
            O => \N__40849\,
            I => \N__40838\
        );

    \I__9385\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40838\
        );

    \I__9384\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40835\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__40846\,
            I => \N__40832\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__40843\,
            I => \N__40824\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__40838\,
            I => \N__40824\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__40835\,
            I => \N__40824\
        );

    \I__9379\ : InMux
    port map (
            O => \N__40832\,
            I => \N__40819\
        );

    \I__9378\ : InMux
    port map (
            O => \N__40831\,
            I => \N__40819\
        );

    \I__9377\ : Odrv12
    port map (
            O => \N__40824\,
            I => \data_out_6__7__N_678\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__40819\,
            I => \data_out_6__7__N_678\
        );

    \I__9375\ : CascadeMux
    port map (
            O => \N__40814\,
            I => \n96_cascade_\
        );

    \I__9374\ : CascadeMux
    port map (
            O => \N__40811\,
            I => \n47_cascade_\
        );

    \I__9373\ : InMux
    port map (
            O => \N__40808\,
            I => \N__40804\
        );

    \I__9372\ : InMux
    port map (
            O => \N__40807\,
            I => \N__40801\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__40804\,
            I => n2615
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__40801\,
            I => n2615
        );

    \I__9369\ : CascadeMux
    port map (
            O => \N__40796\,
            I => \n41_cascade_\
        );

    \I__9368\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40789\
        );

    \I__9367\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40786\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__40789\,
            I => \N__40783\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__40786\,
            I => \N__40780\
        );

    \I__9364\ : Span4Mux_h
    port map (
            O => \N__40783\,
            I => \N__40777\
        );

    \I__9363\ : Odrv4
    port map (
            O => \N__40780\,
            I => \c0.data_out_5__3__N_964\
        );

    \I__9362\ : Odrv4
    port map (
            O => \N__40777\,
            I => \c0.data_out_5__3__N_964\
        );

    \I__9361\ : CascadeMux
    port map (
            O => \N__40772\,
            I => \c0.data_out_5__3__N_964_cascade_\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__40769\,
            I => \c0.data_out_6__3__N_785_cascade_\
        );

    \I__9359\ : InMux
    port map (
            O => \N__40766\,
            I => \N__40762\
        );

    \I__9358\ : CascadeMux
    port map (
            O => \N__40765\,
            I => \N__40759\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__40762\,
            I => \N__40756\
        );

    \I__9356\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40753\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__40756\,
            I => rand_setpoint_19
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__40753\,
            I => rand_setpoint_19
        );

    \I__9353\ : CascadeMux
    port map (
            O => \N__40748\,
            I => \c0.n2181_cascade_\
        );

    \I__9352\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40733\
        );

    \I__9351\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40733\
        );

    \I__9350\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40733\
        );

    \I__9349\ : InMux
    port map (
            O => \N__40742\,
            I => \N__40730\
        );

    \I__9348\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40725\
        );

    \I__9347\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40722\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__40733\,
            I => \N__40717\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__40730\,
            I => \N__40717\
        );

    \I__9344\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40712\
        );

    \I__9343\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40712\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__40725\,
            I => \data_out_6__6__N_729\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__40722\,
            I => \data_out_6__6__N_729\
        );

    \I__9340\ : Odrv12
    port map (
            O => \N__40717\,
            I => \data_out_6__6__N_729\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__40712\,
            I => \data_out_6__6__N_729\
        );

    \I__9338\ : CascadeMux
    port map (
            O => \N__40703\,
            I => \N__40698\
        );

    \I__9337\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40694\
        );

    \I__9336\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40690\
        );

    \I__9335\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40687\
        );

    \I__9334\ : CascadeMux
    port map (
            O => \N__40697\,
            I => \N__40683\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40680\
        );

    \I__9332\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40677\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__40690\,
            I => \N__40674\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__40687\,
            I => \N__40671\
        );

    \I__9329\ : InMux
    port map (
            O => \N__40686\,
            I => \N__40666\
        );

    \I__9328\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40666\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__40680\,
            I => data_out_2_0
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__40677\,
            I => data_out_2_0
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__40674\,
            I => data_out_2_0
        );

    \I__9324\ : Odrv12
    port map (
            O => \N__40671\,
            I => data_out_2_0
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__40666\,
            I => data_out_2_0
        );

    \I__9322\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__40652\,
            I => \N__40649\
        );

    \I__9320\ : Span4Mux_v
    port map (
            O => \N__40649\,
            I => \N__40646\
        );

    \I__9319\ : Odrv4
    port map (
            O => \N__40646\,
            I => \c0.n2_adj_2483\
        );

    \I__9318\ : InMux
    port map (
            O => \N__40643\,
            I => \N__40640\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__40640\,
            I => \c0.n17389\
        );

    \I__9316\ : CascadeMux
    port map (
            O => \N__40637\,
            I => \c0.n17389_cascade_\
        );

    \I__9315\ : CascadeMux
    port map (
            O => \N__40634\,
            I => \c0.n17600_cascade_\
        );

    \I__9314\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40628\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__40628\,
            I => \N__40625\
        );

    \I__9312\ : Span4Mux_h
    port map (
            O => \N__40625\,
            I => \N__40622\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__40622\,
            I => \c0.n9658\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__40619\,
            I => \c0.n17398_cascade_\
        );

    \I__9309\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40612\
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__40615\,
            I => \N__40609\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__40612\,
            I => \N__40606\
        );

    \I__9306\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40603\
        );

    \I__9305\ : Odrv4
    port map (
            O => \N__40606\,
            I => rand_setpoint_20
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__40603\,
            I => rand_setpoint_20
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__40598\,
            I => \c0.n2146_cascade_\
        );

    \I__9302\ : CascadeMux
    port map (
            O => \N__40595\,
            I => \c0.data_out_6__7__N_675_cascade_\
        );

    \I__9301\ : InMux
    port map (
            O => \N__40592\,
            I => \N__40589\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40585\
        );

    \I__9299\ : CascadeMux
    port map (
            O => \N__40588\,
            I => \N__40582\
        );

    \I__9298\ : Span4Mux_h
    port map (
            O => \N__40585\,
            I => \N__40579\
        );

    \I__9297\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40576\
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__40579\,
            I => rand_setpoint_15
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__40576\,
            I => rand_setpoint_15
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__40571\,
            I => \c0.n17928_cascade_\
        );

    \I__9293\ : InMux
    port map (
            O => \N__40568\,
            I => \N__40565\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__40565\,
            I => \N__40562\
        );

    \I__9291\ : Span4Mux_h
    port map (
            O => \N__40562\,
            I => \N__40558\
        );

    \I__9290\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40555\
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__40558\,
            I => rand_setpoint_14
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__40555\,
            I => rand_setpoint_14
        );

    \I__9287\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40547\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__40547\,
            I => \N__40544\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__40544\,
            I => \c0.n17465\
        );

    \I__9284\ : CascadeMux
    port map (
            O => \N__40541\,
            I => \c0.n17906_cascade_\
        );

    \I__9283\ : InMux
    port map (
            O => \N__40538\,
            I => \N__40535\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__40535\,
            I => \N__40532\
        );

    \I__9281\ : Span4Mux_h
    port map (
            O => \N__40532\,
            I => \N__40529\
        );

    \I__9280\ : Odrv4
    port map (
            O => \N__40529\,
            I => \c0.n17921\
        );

    \I__9279\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40523\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__40523\,
            I => \N__40520\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__40520\,
            I => \c0.data_out_10_6\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__40517\,
            I => \c0.n18393_cascade_\
        );

    \I__9275\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40511\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__40511\,
            I => \tx_data_3_N_keep\
        );

    \I__9273\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40505\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__40505\,
            I => \c0.n18095\
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__40502\,
            I => \N__40498\
        );

    \I__9270\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40493\
        );

    \I__9269\ : InMux
    port map (
            O => \N__40498\,
            I => \N__40490\
        );

    \I__9268\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40485\
        );

    \I__9267\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40485\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40482\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__40490\,
            I => \N__40477\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__40485\,
            I => \N__40477\
        );

    \I__9263\ : Odrv4
    port map (
            O => \N__40482\,
            I => n9646
        );

    \I__9262\ : Odrv4
    port map (
            O => \N__40477\,
            I => n9646
        );

    \I__9261\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40468\
        );

    \I__9260\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40465\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__40468\,
            I => n9920
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40465\,
            I => n9920
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__40460\,
            I => \N__40456\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__40459\,
            I => \N__40453\
        );

    \I__9255\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40446\
        );

    \I__9254\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40446\
        );

    \I__9253\ : InMux
    port map (
            O => \N__40452\,
            I => \N__40441\
        );

    \I__9252\ : InMux
    port map (
            O => \N__40451\,
            I => \N__40438\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__40446\,
            I => \N__40435\
        );

    \I__9250\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40430\
        );

    \I__9249\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40430\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__40441\,
            I => \N__40427\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40418\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__40435\,
            I => \N__40418\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40418\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__40427\,
            I => \N__40418\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__40418\,
            I => \r_Bit_Index_0_adj_2627\
        );

    \I__9242\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40408\
        );

    \I__9241\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40408\
        );

    \I__9240\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40405\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__40408\,
            I => \N__40397\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__40405\,
            I => \N__40397\
        );

    \I__9237\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40394\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40389\
        );

    \I__9235\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40389\
        );

    \I__9234\ : Span4Mux_h
    port map (
            O => \N__40397\,
            I => \N__40386\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__40394\,
            I => \r_SM_Main_2_N_2323_1\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__40389\,
            I => \r_SM_Main_2_N_2323_1\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__40386\,
            I => \r_SM_Main_2_N_2323_1\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__40379\,
            I => \n4_adj_2653_cascade_\
        );

    \I__9229\ : CascadeMux
    port map (
            O => \N__40376\,
            I => \N__40366\
        );

    \I__9228\ : InMux
    port map (
            O => \N__40375\,
            I => \N__40363\
        );

    \I__9227\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40354\
        );

    \I__9226\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40354\
        );

    \I__9225\ : InMux
    port map (
            O => \N__40372\,
            I => \N__40354\
        );

    \I__9224\ : InMux
    port map (
            O => \N__40371\,
            I => \N__40354\
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__40370\,
            I => \N__40351\
        );

    \I__9222\ : CascadeMux
    port map (
            O => \N__40369\,
            I => \N__40347\
        );

    \I__9221\ : InMux
    port map (
            O => \N__40366\,
            I => \N__40343\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40363\,
            I => \N__40340\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__40354\,
            I => \N__40334\
        );

    \I__9218\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40329\
        );

    \I__9217\ : InMux
    port map (
            O => \N__40350\,
            I => \N__40329\
        );

    \I__9216\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40326\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40346\,
            I => \N__40321\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__40343\,
            I => \N__40316\
        );

    \I__9213\ : Span4Mux_h
    port map (
            O => \N__40340\,
            I => \N__40316\
        );

    \I__9212\ : InMux
    port map (
            O => \N__40339\,
            I => \N__40313\
        );

    \I__9211\ : InMux
    port map (
            O => \N__40338\,
            I => \N__40308\
        );

    \I__9210\ : InMux
    port map (
            O => \N__40337\,
            I => \N__40308\
        );

    \I__9209\ : Span4Mux_h
    port map (
            O => \N__40334\,
            I => \N__40305\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__40329\,
            I => \N__40302\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__40326\,
            I => \N__40299\
        );

    \I__9206\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40294\
        );

    \I__9205\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40294\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40281\
        );

    \I__9203\ : Span4Mux_v
    port map (
            O => \N__40316\,
            I => \N__40281\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__40313\,
            I => \N__40281\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__40308\,
            I => \N__40278\
        );

    \I__9200\ : Span4Mux_h
    port map (
            O => \N__40305\,
            I => \N__40273\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__40302\,
            I => \N__40273\
        );

    \I__9198\ : Span4Mux_v
    port map (
            O => \N__40299\,
            I => \N__40268\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__40294\,
            I => \N__40268\
        );

    \I__9196\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40259\
        );

    \I__9195\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40259\
        );

    \I__9194\ : InMux
    port map (
            O => \N__40291\,
            I => \N__40259\
        );

    \I__9193\ : InMux
    port map (
            O => \N__40290\,
            I => \N__40259\
        );

    \I__9192\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40254\
        );

    \I__9191\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40254\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__40281\,
            I => \r_SM_Main_2\
        );

    \I__9189\ : Odrv12
    port map (
            O => \N__40278\,
            I => \r_SM_Main_2\
        );

    \I__9188\ : Odrv4
    port map (
            O => \N__40273\,
            I => \r_SM_Main_2\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__40268\,
            I => \r_SM_Main_2\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__40259\,
            I => \r_SM_Main_2\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__40254\,
            I => \r_SM_Main_2\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__40241\,
            I => \N__40234\
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__40240\,
            I => \N__40231\
        );

    \I__9182\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40226\
        );

    \I__9181\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40226\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__40237\,
            I => \N__40223\
        );

    \I__9179\ : InMux
    port map (
            O => \N__40234\,
            I => \N__40216\
        );

    \I__9178\ : InMux
    port map (
            O => \N__40231\,
            I => \N__40216\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__40226\,
            I => \N__40210\
        );

    \I__9176\ : InMux
    port map (
            O => \N__40223\,
            I => \N__40207\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__40222\,
            I => \N__40203\
        );

    \I__9174\ : InMux
    port map (
            O => \N__40221\,
            I => \N__40200\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40197\
        );

    \I__9172\ : InMux
    port map (
            O => \N__40215\,
            I => \N__40194\
        );

    \I__9171\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40191\
        );

    \I__9170\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40188\
        );

    \I__9169\ : Span4Mux_h
    port map (
            O => \N__40210\,
            I => \N__40183\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__40207\,
            I => \N__40183\
        );

    \I__9167\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40178\
        );

    \I__9166\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40178\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__40200\,
            I => \r_SM_Main_0\
        );

    \I__9164\ : Odrv12
    port map (
            O => \N__40197\,
            I => \r_SM_Main_0\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__40194\,
            I => \r_SM_Main_0\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__40191\,
            I => \r_SM_Main_0\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__40188\,
            I => \r_SM_Main_0\
        );

    \I__9160\ : Odrv4
    port map (
            O => \N__40183\,
            I => \r_SM_Main_0\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__40178\,
            I => \r_SM_Main_0\
        );

    \I__9158\ : CascadeMux
    port map (
            O => \N__40163\,
            I => \N__40156\
        );

    \I__9157\ : CascadeMux
    port map (
            O => \N__40162\,
            I => \N__40150\
        );

    \I__9156\ : CascadeMux
    port map (
            O => \N__40161\,
            I => \N__40147\
        );

    \I__9155\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40142\
        );

    \I__9154\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40137\
        );

    \I__9153\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40137\
        );

    \I__9152\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40134\
        );

    \I__9151\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40130\
        );

    \I__9150\ : InMux
    port map (
            O => \N__40153\,
            I => \N__40123\
        );

    \I__9149\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40123\
        );

    \I__9148\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40123\
        );

    \I__9147\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40120\
        );

    \I__9146\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40117\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__40142\,
            I => \N__40112\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__40137\,
            I => \N__40112\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__40134\,
            I => \N__40109\
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__40133\,
            I => \N__40104\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40096\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__40123\,
            I => \N__40096\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__40120\,
            I => \N__40091\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__40117\,
            I => \N__40091\
        );

    \I__9137\ : Span4Mux_v
    port map (
            O => \N__40112\,
            I => \N__40086\
        );

    \I__9136\ : Span4Mux_h
    port map (
            O => \N__40109\,
            I => \N__40086\
        );

    \I__9135\ : InMux
    port map (
            O => \N__40108\,
            I => \N__40077\
        );

    \I__9134\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40077\
        );

    \I__9133\ : InMux
    port map (
            O => \N__40104\,
            I => \N__40077\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40077\
        );

    \I__9131\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40072\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40072\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__40096\,
            I => \r_SM_Main_1\
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__40091\,
            I => \r_SM_Main_1\
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__40086\,
            I => \r_SM_Main_1\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__40077\,
            I => \r_SM_Main_1\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__40072\,
            I => \r_SM_Main_1\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40061\,
            I => \N__40058\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__40058\,
            I => \c0.tx_active_prev\
        );

    \I__9122\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40051\
        );

    \I__9121\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40048\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__40051\,
            I => \c0.n17349\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__40048\,
            I => \c0.n17349\
        );

    \I__9118\ : InMux
    port map (
            O => \N__40043\,
            I => \N__40040\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__40040\,
            I => \c0.n17937\
        );

    \I__9116\ : CascadeMux
    port map (
            O => \N__40037\,
            I => \c0.n18390_cascade_\
        );

    \I__9115\ : InMux
    port map (
            O => \N__40034\,
            I => \c0.n16311\
        );

    \I__9114\ : InMux
    port map (
            O => \N__40031\,
            I => \N__40028\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__9112\ : Odrv4
    port map (
            O => \N__40025\,
            I => \c0.n18011\
        );

    \I__9111\ : InMux
    port map (
            O => \N__40022\,
            I => \bfn_12_25_0_\
        );

    \I__9110\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40016\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__40016\,
            I => \c0.n7266\
        );

    \I__9108\ : InMux
    port map (
            O => \N__40013\,
            I => \c0.n16313\
        );

    \I__9107\ : CascadeMux
    port map (
            O => \N__40010\,
            I => \N__40007\
        );

    \I__9106\ : InMux
    port map (
            O => \N__40007\,
            I => \N__40004\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__40004\,
            I => \N__40001\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__40001\,
            I => \c0.n7265\
        );

    \I__9103\ : InMux
    port map (
            O => \N__39998\,
            I => \c0.n16314\
        );

    \I__9102\ : InMux
    port map (
            O => \N__39995\,
            I => \c0.n16315\
        );

    \I__9101\ : InMux
    port map (
            O => \N__39992\,
            I => \c0.n16316\
        );

    \I__9100\ : InMux
    port map (
            O => \N__39989\,
            I => \c0.n16317\
        );

    \I__9099\ : InMux
    port map (
            O => \N__39986\,
            I => \c0.n16318\
        );

    \I__9098\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39980\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__39980\,
            I => \c0.n25_adj_2517\
        );

    \I__9096\ : CascadeMux
    port map (
            O => \N__39977\,
            I => \c0.n1314_cascade_\
        );

    \I__9095\ : InMux
    port map (
            O => \N__39974\,
            I => \bfn_12_24_0_\
        );

    \I__9094\ : InMux
    port map (
            O => \N__39971\,
            I => \c0.n16305\
        );

    \I__9093\ : InMux
    port map (
            O => \N__39968\,
            I => \N__39965\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__39965\,
            I => \c0.n7273\
        );

    \I__9091\ : InMux
    port map (
            O => \N__39962\,
            I => \c0.n16306\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__39959\,
            I => \N__39956\
        );

    \I__9089\ : InMux
    port map (
            O => \N__39956\,
            I => \N__39953\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__39953\,
            I => \c0.n7272\
        );

    \I__9087\ : InMux
    port map (
            O => \N__39950\,
            I => \c0.n16307\
        );

    \I__9086\ : InMux
    port map (
            O => \N__39947\,
            I => \c0.n16308\
        );

    \I__9085\ : InMux
    port map (
            O => \N__39944\,
            I => \c0.n16309\
        );

    \I__9084\ : InMux
    port map (
            O => \N__39941\,
            I => \N__39938\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__39938\,
            I => \c0.n7269\
        );

    \I__9082\ : InMux
    port map (
            O => \N__39935\,
            I => \c0.n16310\
        );

    \I__9081\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39928\
        );

    \I__9080\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39925\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__39928\,
            I => \N__39922\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__39925\,
            I => \N__39919\
        );

    \I__9077\ : Span4Mux_h
    port map (
            O => \N__39922\,
            I => \N__39915\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__39919\,
            I => \N__39912\
        );

    \I__9075\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39909\
        );

    \I__9074\ : Span4Mux_h
    port map (
            O => \N__39915\,
            I => \N__39906\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__39912\,
            I => \c0.data_in_6_1\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__39909\,
            I => \c0.data_in_6_1\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__39906\,
            I => \c0.data_in_6_1\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__39899\,
            I => \N__39896\
        );

    \I__9069\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39893\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__39893\,
            I => \N__39889\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__39892\,
            I => \N__39886\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__39889\,
            I => \N__39882\
        );

    \I__9065\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39879\
        );

    \I__9064\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39875\
        );

    \I__9063\ : Span4Mux_s1_h
    port map (
            O => \N__39882\,
            I => \N__39872\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__39879\,
            I => \N__39869\
        );

    \I__9061\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39866\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39863\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__39872\,
            I => \N__39858\
        );

    \I__9058\ : Span4Mux_v
    port map (
            O => \N__39869\,
            I => \N__39858\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__39866\,
            I => \N__39853\
        );

    \I__9056\ : Span4Mux_v
    port map (
            O => \N__39863\,
            I => \N__39853\
        );

    \I__9055\ : Span4Mux_h
    port map (
            O => \N__39858\,
            I => \N__39850\
        );

    \I__9054\ : Odrv4
    port map (
            O => \N__39853\,
            I => data_in_5_1
        );

    \I__9053\ : Odrv4
    port map (
            O => \N__39850\,
            I => data_in_5_1
        );

    \I__9052\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39841\
        );

    \I__9051\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39838\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__39841\,
            I => \N__39835\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39831\
        );

    \I__9048\ : Span4Mux_h
    port map (
            O => \N__39835\,
            I => \N__39828\
        );

    \I__9047\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39825\
        );

    \I__9046\ : Span4Mux_h
    port map (
            O => \N__39831\,
            I => \N__39822\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__39828\,
            I => \N__39819\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__39825\,
            I => data_in_10_6
        );

    \I__9043\ : Odrv4
    port map (
            O => \N__39822\,
            I => data_in_10_6
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__39819\,
            I => data_in_10_6
        );

    \I__9041\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39808\
        );

    \I__9040\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__39808\,
            I => data_in_11_6
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__39805\,
            I => data_in_11_6
        );

    \I__9037\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39797\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__39797\,
            I => \N__39794\
        );

    \I__9035\ : Odrv4
    port map (
            O => \N__39794\,
            I => \c0.n17755\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__39791\,
            I => \c0.n17525_cascade_\
        );

    \I__9033\ : InMux
    port map (
            O => \N__39788\,
            I => \N__39785\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__39785\,
            I => \N__39782\
        );

    \I__9031\ : Odrv4
    port map (
            O => \N__39782\,
            I => \c0.rx.n9553\
        );

    \I__9030\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39775\
        );

    \I__9029\ : InMux
    port map (
            O => \N__39778\,
            I => \N__39768\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__39775\,
            I => \N__39765\
        );

    \I__9027\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39758\
        );

    \I__9026\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39758\
        );

    \I__9025\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39758\
        );

    \I__9024\ : CascadeMux
    port map (
            O => \N__39771\,
            I => \N__39755\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__39768\,
            I => \N__39749\
        );

    \I__9022\ : Span4Mux_s2_v
    port map (
            O => \N__39765\,
            I => \N__39744\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39744\
        );

    \I__9020\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39735\
        );

    \I__9019\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39735\
        );

    \I__9018\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39735\
        );

    \I__9017\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39735\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__39749\,
            I => \N__39732\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__39744\,
            I => \N__39729\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__39735\,
            I => \N__39726\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__39732\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__9012\ : Odrv4
    port map (
            O => \N__39729\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__39726\,
            I => \c0.rx.r_SM_Main_2\
        );

    \I__9010\ : CascadeMux
    port map (
            O => \N__39719\,
            I => \N__39714\
        );

    \I__9009\ : InMux
    port map (
            O => \N__39718\,
            I => \N__39707\
        );

    \I__9008\ : InMux
    port map (
            O => \N__39717\,
            I => \N__39704\
        );

    \I__9007\ : InMux
    port map (
            O => \N__39714\,
            I => \N__39697\
        );

    \I__9006\ : InMux
    port map (
            O => \N__39713\,
            I => \N__39697\
        );

    \I__9005\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39697\
        );

    \I__9004\ : InMux
    port map (
            O => \N__39711\,
            I => \N__39694\
        );

    \I__9003\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39691\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__39707\,
            I => \N__39684\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39675\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__39697\,
            I => \N__39675\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__39694\,
            I => \N__39675\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__39691\,
            I => \N__39675\
        );

    \I__8997\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39666\
        );

    \I__8996\ : InMux
    port map (
            O => \N__39689\,
            I => \N__39666\
        );

    \I__8995\ : InMux
    port map (
            O => \N__39688\,
            I => \N__39666\
        );

    \I__8994\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39666\
        );

    \I__8993\ : Span4Mux_v
    port map (
            O => \N__39684\,
            I => \N__39661\
        );

    \I__8992\ : Span4Mux_s3_v
    port map (
            O => \N__39675\,
            I => \N__39661\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__39666\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__39661\,
            I => \c0.rx.r_SM_Main_1\
        );

    \I__8989\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39651\
        );

    \I__8988\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39645\
        );

    \I__8987\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39645\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__39651\,
            I => \N__39642\
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__39650\,
            I => \N__39638\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39635\
        );

    \I__8983\ : Span4Mux_s2_v
    port map (
            O => \N__39642\,
            I => \N__39632\
        );

    \I__8982\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39626\
        );

    \I__8981\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39626\
        );

    \I__8980\ : Span4Mux_h
    port map (
            O => \N__39635\,
            I => \N__39623\
        );

    \I__8979\ : Sp12to4
    port map (
            O => \N__39632\,
            I => \N__39620\
        );

    \I__8978\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39617\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__39626\,
            I => \c0.rx.r_SM_Main_2_N_2380_2\
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__39623\,
            I => \c0.rx.r_SM_Main_2_N_2380_2\
        );

    \I__8975\ : Odrv12
    port map (
            O => \N__39620\,
            I => \c0.rx.r_SM_Main_2_N_2380_2\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__39617\,
            I => \c0.rx.r_SM_Main_2_N_2380_2\
        );

    \I__8973\ : SRMux
    port map (
            O => \N__39608\,
            I => \N__39605\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8971\ : Span4Mux_s2_v
    port map (
            O => \N__39602\,
            I => \N__39599\
        );

    \I__8970\ : Span4Mux_h
    port map (
            O => \N__39599\,
            I => \N__39596\
        );

    \I__8969\ : Span4Mux_s2_v
    port map (
            O => \N__39596\,
            I => \N__39593\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__39593\,
            I => \c0.rx.n17351\
        );

    \I__8967\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39581\
        );

    \I__8966\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39572\
        );

    \I__8965\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39572\
        );

    \I__8964\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39572\
        );

    \I__8963\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39572\
        );

    \I__8962\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39566\
        );

    \I__8961\ : InMux
    port map (
            O => \N__39584\,
            I => \N__39566\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__39581\,
            I => \N__39560\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__39572\,
            I => \N__39560\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39557\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__39566\,
            I => \N__39553\
        );

    \I__8956\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39550\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__39560\,
            I => \N__39547\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__39557\,
            I => \N__39544\
        );

    \I__8953\ : InMux
    port map (
            O => \N__39556\,
            I => \N__39541\
        );

    \I__8952\ : Span4Mux_h
    port map (
            O => \N__39553\,
            I => \N__39536\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__39550\,
            I => \N__39536\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__39547\,
            I => \N__39533\
        );

    \I__8949\ : Span12Mux_v
    port map (
            O => \N__39544\,
            I => \N__39528\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__39541\,
            I => \N__39528\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__39536\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__8946\ : Odrv4
    port map (
            O => \N__39533\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__8945\ : Odrv12
    port map (
            O => \N__39528\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__8944\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39518\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__39518\,
            I => \N__39515\
        );

    \I__8942\ : Span4Mux_h
    port map (
            O => \N__39515\,
            I => \N__39512\
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__39512\,
            I => \c0.rx.n17376\
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__39509\,
            I => \c0.data_out_6__2__N_803_cascade_\
        );

    \I__8939\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39502\
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__39505\,
            I => \N__39499\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__39502\,
            I => \N__39496\
        );

    \I__8936\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39493\
        );

    \I__8935\ : Odrv4
    port map (
            O => \N__39496\,
            I => rand_setpoint_18
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__39493\,
            I => rand_setpoint_18
        );

    \I__8933\ : CascadeMux
    port map (
            O => \N__39488\,
            I => \c0.n2216_cascade_\
        );

    \I__8932\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39481\
        );

    \I__8931\ : InMux
    port map (
            O => \N__39484\,
            I => \N__39478\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__39481\,
            I => \N__39475\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__39478\,
            I => \N__39470\
        );

    \I__8928\ : Span4Mux_v
    port map (
            O => \N__39475\,
            I => \N__39470\
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__39470\,
            I => \c0.data_out_6_2\
        );

    \I__8926\ : InMux
    port map (
            O => \N__39467\,
            I => \N__39464\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39464\,
            I => \N__39460\
        );

    \I__8924\ : CascadeMux
    port map (
            O => \N__39463\,
            I => \N__39457\
        );

    \I__8923\ : Span4Mux_h
    port map (
            O => \N__39460\,
            I => \N__39454\
        );

    \I__8922\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39451\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__39454\,
            I => rand_setpoint_26
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__39451\,
            I => rand_setpoint_26
        );

    \I__8919\ : InMux
    port map (
            O => \N__39446\,
            I => \N__39443\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__39443\,
            I => \c0.data_out_6__2__N_803\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__39440\,
            I => \c0.n17964_cascade_\
        );

    \I__8916\ : InMux
    port map (
            O => \N__39437\,
            I => \N__39433\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__39436\,
            I => \N__39430\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__39433\,
            I => \N__39427\
        );

    \I__8913\ : InMux
    port map (
            O => \N__39430\,
            I => \N__39424\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__39427\,
            I => rand_setpoint_0
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__39424\,
            I => rand_setpoint_0
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__39419\,
            I => \c0.n8953_cascade_\
        );

    \I__8909\ : InMux
    port map (
            O => \N__39416\,
            I => \N__39413\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__39413\,
            I => \N__39409\
        );

    \I__8907\ : CascadeMux
    port map (
            O => \N__39412\,
            I => \N__39406\
        );

    \I__8906\ : Span4Mux_h
    port map (
            O => \N__39409\,
            I => \N__39403\
        );

    \I__8905\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39400\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__39403\,
            I => rand_setpoint_5
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__39400\,
            I => rand_setpoint_5
        );

    \I__8902\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39392\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__39392\,
            I => \N__39389\
        );

    \I__8900\ : Sp12to4
    port map (
            O => \N__39389\,
            I => \N__39386\
        );

    \I__8899\ : Odrv12
    port map (
            O => \N__39386\,
            I => \c0.n5\
        );

    \I__8898\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39380\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__39380\,
            I => \c0.n17972\
        );

    \I__8896\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39374\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__39374\,
            I => \c0.n18501\
        );

    \I__8894\ : CascadeMux
    port map (
            O => \N__39371\,
            I => \tx_data_0_N_keep_cascade_\
        );

    \I__8893\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39364\
        );

    \I__8892\ : InMux
    port map (
            O => \N__39367\,
            I => \N__39361\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__39364\,
            I => \N__39358\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__39361\,
            I => \r_Tx_Data_0\
        );

    \I__8889\ : Odrv12
    port map (
            O => \N__39358\,
            I => \r_Tx_Data_0\
        );

    \I__8888\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39350\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__39350\,
            I => \N__39346\
        );

    \I__8886\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39343\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__39346\,
            I => \N__39340\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__39343\,
            I => data_in_15_5
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__39340\,
            I => data_in_15_5
        );

    \I__8882\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39332\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__39332\,
            I => \N__39328\
        );

    \I__8880\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39325\
        );

    \I__8879\ : Odrv12
    port map (
            O => \N__39328\,
            I => data_in_14_5
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__39325\,
            I => data_in_14_5
        );

    \I__8877\ : InMux
    port map (
            O => \N__39320\,
            I => \N__39317\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__39317\,
            I => n4958
        );

    \I__8875\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39308\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39308\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39304\
        );

    \I__8872\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39301\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__39304\,
            I => \N__39297\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__39301\,
            I => \N__39294\
        );

    \I__8869\ : InMux
    port map (
            O => \N__39300\,
            I => \N__39291\
        );

    \I__8868\ : Span4Mux_h
    port map (
            O => \N__39297\,
            I => \N__39287\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__39294\,
            I => \N__39282\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__39291\,
            I => \N__39279\
        );

    \I__8865\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39276\
        );

    \I__8864\ : Sp12to4
    port map (
            O => \N__39287\,
            I => \N__39273\
        );

    \I__8863\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39270\
        );

    \I__8862\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39267\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__39282\,
            I => \N__39262\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__39279\,
            I => \N__39262\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__39276\,
            I => \r_Bit_Index_2_adj_2625\
        );

    \I__8858\ : Odrv12
    port map (
            O => \N__39273\,
            I => \r_Bit_Index_2_adj_2625\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__39270\,
            I => \r_Bit_Index_2_adj_2625\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__39267\,
            I => \r_Bit_Index_2_adj_2625\
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__39262\,
            I => \r_Bit_Index_2_adj_2625\
        );

    \I__8854\ : CascadeMux
    port map (
            O => \N__39251\,
            I => \n4958_cascade_\
        );

    \I__8853\ : CascadeMux
    port map (
            O => \N__39248\,
            I => \n9920_cascade_\
        );

    \I__8852\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39242\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__39242\,
            I => \N__39237\
        );

    \I__8850\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39231\
        );

    \I__8849\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39231\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__39237\,
            I => \N__39225\
        );

    \I__8847\ : InMux
    port map (
            O => \N__39236\,
            I => \N__39222\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__39231\,
            I => \N__39219\
        );

    \I__8845\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39216\
        );

    \I__8844\ : InMux
    port map (
            O => \N__39229\,
            I => \N__39211\
        );

    \I__8843\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39211\
        );

    \I__8842\ : Span4Mux_h
    port map (
            O => \N__39225\,
            I => \N__39206\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39206\
        );

    \I__8840\ : Span12Mux_v
    port map (
            O => \N__39219\,
            I => \N__39203\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__39216\,
            I => \r_Bit_Index_1_adj_2626\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__39211\,
            I => \r_Bit_Index_1_adj_2626\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__39206\,
            I => \r_Bit_Index_1_adj_2626\
        );

    \I__8836\ : Odrv12
    port map (
            O => \N__39203\,
            I => \r_Bit_Index_1_adj_2626\
        );

    \I__8835\ : InMux
    port map (
            O => \N__39194\,
            I => \N__39191\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__39191\,
            I => \N__39187\
        );

    \I__8833\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39184\
        );

    \I__8832\ : Odrv4
    port map (
            O => \N__39187\,
            I => data_in_15_0
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__39184\,
            I => data_in_15_0
        );

    \I__8830\ : InMux
    port map (
            O => \N__39179\,
            I => \N__39176\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__39176\,
            I => \N__39172\
        );

    \I__8828\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39169\
        );

    \I__8827\ : Odrv4
    port map (
            O => \N__39172\,
            I => data_in_14_0
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__39169\,
            I => data_in_14_0
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__39164\,
            I => \N__39161\
        );

    \I__8824\ : InMux
    port map (
            O => \N__39161\,
            I => \N__39157\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__39160\,
            I => \N__39154\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__39157\,
            I => \N__39151\
        );

    \I__8821\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39148\
        );

    \I__8820\ : Odrv12
    port map (
            O => \N__39151\,
            I => rand_setpoint_1
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__39148\,
            I => rand_setpoint_1
        );

    \I__8818\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39140\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__39140\,
            I => n18438
        );

    \I__8816\ : CascadeMux
    port map (
            O => \N__39137\,
            I => \N__39134\
        );

    \I__8815\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39131\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__39131\,
            I => \N__39127\
        );

    \I__8813\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39119\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__39127\,
            I => \N__39116\
        );

    \I__8811\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39113\
        );

    \I__8810\ : InMux
    port map (
            O => \N__39125\,
            I => \N__39108\
        );

    \I__8809\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39108\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__39123\,
            I => \N__39104\
        );

    \I__8807\ : InMux
    port map (
            O => \N__39122\,
            I => \N__39101\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__39119\,
            I => \N__39096\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__39116\,
            I => \N__39096\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__39113\,
            I => \N__39091\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__39108\,
            I => \N__39091\
        );

    \I__8802\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39086\
        );

    \I__8801\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39086\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__39101\,
            I => \r_Bit_Index_1\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__39096\,
            I => \r_Bit_Index_1\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__39091\,
            I => \r_Bit_Index_1\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__39086\,
            I => \r_Bit_Index_1\
        );

    \I__8796\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39074\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__39074\,
            I => \N__39071\
        );

    \I__8794\ : Odrv4
    port map (
            O => \N__39071\,
            I => n18441
        );

    \I__8793\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39065\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__39065\,
            I => \N__39061\
        );

    \I__8791\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39058\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__39061\,
            I => data_in_13_0
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__39058\,
            I => data_in_13_0
        );

    \I__8788\ : InMux
    port map (
            O => \N__39053\,
            I => \N__39049\
        );

    \I__8787\ : InMux
    port map (
            O => \N__39052\,
            I => \N__39046\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__39049\,
            I => \r_Tx_Data_3\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__39046\,
            I => \r_Tx_Data_3\
        );

    \I__8784\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39037\
        );

    \I__8783\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39034\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39037\,
            I => data_in_20_1
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__39034\,
            I => data_in_20_1
        );

    \I__8780\ : InMux
    port map (
            O => \N__39029\,
            I => \N__39023\
        );

    \I__8779\ : InMux
    port map (
            O => \N__39028\,
            I => \N__39023\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__39023\,
            I => data_in_19_1
        );

    \I__8777\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39016\
        );

    \I__8776\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39013\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__39016\,
            I => data_in_17_0
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__39013\,
            I => data_in_17_0
        );

    \I__8773\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39002\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39007\,
            I => \N__39002\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__39002\,
            I => data_in_16_0
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__38999\,
            I => \n17737_cascade_\
        );

    \I__8769\ : InMux
    port map (
            O => \N__38996\,
            I => \N__38993\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__38993\,
            I => n17312
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__38990\,
            I => \n17312_cascade_\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \n14_adj_2615_cascade_\
        );

    \I__8765\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38980\
        );

    \I__8764\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38977\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__38980\,
            I => data_in_17_1
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__38977\,
            I => data_in_17_1
        );

    \I__8761\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38969\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__38969\,
            I => \N__38966\
        );

    \I__8759\ : Span4Mux_h
    port map (
            O => \N__38966\,
            I => \N__38962\
        );

    \I__8758\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38959\
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__38962\,
            I => data_in_16_1
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__38959\,
            I => data_in_16_1
        );

    \I__8755\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38951\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__38951\,
            I => \N__38947\
        );

    \I__8753\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38944\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__38947\,
            I => \N__38940\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__38944\,
            I => \N__38937\
        );

    \I__8750\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38934\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__38940\,
            I => n17757
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__38937\,
            I => n17757
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__38934\,
            I => n17757
        );

    \I__8746\ : CascadeMux
    port map (
            O => \N__38927\,
            I => \N__38922\
        );

    \I__8745\ : CascadeMux
    port map (
            O => \N__38926\,
            I => \N__38919\
        );

    \I__8744\ : CascadeMux
    port map (
            O => \N__38925\,
            I => \N__38915\
        );

    \I__8743\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38912\
        );

    \I__8742\ : InMux
    port map (
            O => \N__38919\,
            I => \N__38907\
        );

    \I__8741\ : InMux
    port map (
            O => \N__38918\,
            I => \N__38907\
        );

    \I__8740\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38902\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__38912\,
            I => \N__38899\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38896\
        );

    \I__8737\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38893\
        );

    \I__8736\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38890\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38887\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__38899\,
            I => \N__38880\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__38896\,
            I => \N__38880\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38880\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__38890\,
            I => \r_Bit_Index_0\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__38887\,
            I => \r_Bit_Index_0\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__38880\,
            I => \r_Bit_Index_0\
        );

    \I__8728\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38869\
        );

    \I__8727\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38866\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__38869\,
            I => data_in_18_1
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__38866\,
            I => data_in_18_1
        );

    \I__8724\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38855\
        );

    \I__8723\ : InMux
    port map (
            O => \N__38860\,
            I => \N__38855\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__38855\,
            I => data_in_19_3
        );

    \I__8721\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38846\
        );

    \I__8720\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38846\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__38846\,
            I => data_in_18_3
        );

    \I__8718\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38839\
        );

    \I__8717\ : InMux
    port map (
            O => \N__38842\,
            I => \N__38836\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__38839\,
            I => \N__38833\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__38836\,
            I => data_in_12_0
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__38833\,
            I => data_in_12_0
        );

    \I__8713\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38825\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__38825\,
            I => \N__38821\
        );

    \I__8711\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38818\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__38821\,
            I => data_in_12_3
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__38818\,
            I => data_in_12_3
        );

    \I__8708\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38810\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__38810\,
            I => n18462
        );

    \I__8706\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38804\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__38804\,
            I => n18465
        );

    \I__8704\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38797\
        );

    \I__8703\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38794\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__38797\,
            I => \N__38791\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__38794\,
            I => \N__38787\
        );

    \I__8700\ : Span4Mux_v
    port map (
            O => \N__38791\,
            I => \N__38784\
        );

    \I__8699\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38781\
        );

    \I__8698\ : Span4Mux_h
    port map (
            O => \N__38787\,
            I => \N__38778\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__38784\,
            I => \N__38775\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__38781\,
            I => data_in_9_6
        );

    \I__8695\ : Odrv4
    port map (
            O => \N__38778\,
            I => data_in_9_6
        );

    \I__8694\ : Odrv4
    port map (
            O => \N__38775\,
            I => data_in_9_6
        );

    \I__8693\ : CascadeMux
    port map (
            O => \N__38768\,
            I => \N__38765\
        );

    \I__8692\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__38762\,
            I => \N__38758\
        );

    \I__8690\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38755\
        );

    \I__8689\ : Span4Mux_v
    port map (
            O => \N__38758\,
            I => \N__38752\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__38755\,
            I => \N__38749\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__38752\,
            I => \N__38744\
        );

    \I__8686\ : Span4Mux_h
    port map (
            O => \N__38749\,
            I => \N__38744\
        );

    \I__8685\ : Span4Mux_h
    port map (
            O => \N__38744\,
            I => \N__38740\
        );

    \I__8684\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38737\
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__38740\,
            I => data_in_8_6
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__38737\,
            I => data_in_8_6
        );

    \I__8681\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__38729\,
            I => \N__38726\
        );

    \I__8679\ : Span4Mux_h
    port map (
            O => \N__38726\,
            I => \N__38722\
        );

    \I__8678\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38719\
        );

    \I__8677\ : Odrv4
    port map (
            O => \N__38722\,
            I => data_in_16_5
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__38719\,
            I => data_in_16_5
        );

    \I__8675\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38710\
        );

    \I__8674\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38707\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__38710\,
            I => data_in_14_3
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__38707\,
            I => data_in_14_3
        );

    \I__8671\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38696\
        );

    \I__8670\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38696\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__38696\,
            I => data_in_13_3
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__38693\,
            I => \c0.n18429_cascade_\
        );

    \I__8667\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38687\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38684\
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__38684\,
            I => \tx_data_7_N_keep\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__38681\,
            I => \c0.n18017_cascade_\
        );

    \I__8663\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__38675\,
            I => \c0.n18426\
        );

    \I__8661\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38668\
        );

    \I__8660\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38665\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__38668\,
            I => data_in_17_3
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__38665\,
            I => data_in_17_3
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__38660\,
            I => \N__38657\
        );

    \I__8656\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38651\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__38651\,
            I => \N__38648\
        );

    \I__8653\ : Odrv4
    port map (
            O => \N__38648\,
            I => \c0.n5_adj_2499\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__38645\,
            I => \c0.n18378_cascade_\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__38642\,
            I => \c0.n18381_cascade_\
        );

    \I__8650\ : InMux
    port map (
            O => \N__38639\,
            I => \N__38636\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__38636\,
            I => \tx_data_2_N_keep\
        );

    \I__8648\ : InMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8646\ : Span4Mux_h
    port map (
            O => \N__38627\,
            I => \N__38623\
        );

    \I__8645\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38620\
        );

    \I__8644\ : Odrv4
    port map (
            O => \N__38623\,
            I => data_in_20_3
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__38620\,
            I => data_in_20_3
        );

    \I__8642\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38612\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__38612\,
            I => \N__38609\
        );

    \I__8640\ : Span4Mux_v
    port map (
            O => \N__38609\,
            I => \N__38605\
        );

    \I__8639\ : InMux
    port map (
            O => \N__38608\,
            I => \N__38602\
        );

    \I__8638\ : Odrv4
    port map (
            O => \N__38605\,
            I => data_in_13_5
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__38602\,
            I => data_in_13_5
        );

    \I__8636\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38591\
        );

    \I__8635\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38591\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__38591\,
            I => data_in_12_4
        );

    \I__8633\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38582\
        );

    \I__8632\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38582\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__38582\,
            I => data_in_13_4
        );

    \I__8630\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38573\
        );

    \I__8629\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38573\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__38573\,
            I => data_in_14_4
        );

    \I__8627\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38566\
        );

    \I__8626\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38563\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__38566\,
            I => data_in_11_3
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__38563\,
            I => data_in_11_3
        );

    \I__8623\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38554\
        );

    \I__8622\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38551\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__38554\,
            I => data_in_15_4
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__38551\,
            I => data_in_15_4
        );

    \I__8619\ : InMux
    port map (
            O => \N__38546\,
            I => \N__38543\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__38543\,
            I => \N__38540\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__38540\,
            I => \N__38537\
        );

    \I__8616\ : Span4Mux_v
    port map (
            O => \N__38537\,
            I => \N__38533\
        );

    \I__8615\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38530\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__38533\,
            I => data_in_17_4
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__38530\,
            I => data_in_17_4
        );

    \I__8612\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38521\
        );

    \I__8611\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38518\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__38521\,
            I => data_in_16_4
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__38518\,
            I => data_in_16_4
        );

    \I__8608\ : CascadeMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__8607\ : InMux
    port map (
            O => \N__38510\,
            I => \N__38507\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__38507\,
            I => \N__38503\
        );

    \I__8605\ : InMux
    port map (
            O => \N__38506\,
            I => \N__38500\
        );

    \I__8604\ : Span4Mux_h
    port map (
            O => \N__38503\,
            I => \N__38497\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__38500\,
            I => \N__38494\
        );

    \I__8602\ : Span4Mux_h
    port map (
            O => \N__38497\,
            I => \N__38490\
        );

    \I__8601\ : Span4Mux_h
    port map (
            O => \N__38494\,
            I => \N__38487\
        );

    \I__8600\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38484\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__38490\,
            I => data_in_4_1
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__38487\,
            I => data_in_4_1
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__38484\,
            I => data_in_4_1
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__38477\,
            I => \c0.n18089_cascade_\
        );

    \I__8595\ : InMux
    port map (
            O => \N__38474\,
            I => \N__38471\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8593\ : Span4Mux_s2_v
    port map (
            O => \N__38468\,
            I => \N__38465\
        );

    \I__8592\ : Span4Mux_h
    port map (
            O => \N__38465\,
            I => \N__38461\
        );

    \I__8591\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38458\
        );

    \I__8590\ : Odrv4
    port map (
            O => \N__38461\,
            I => data_in_19_2
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__38458\,
            I => data_in_19_2
        );

    \I__8588\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38450\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38447\
        );

    \I__8586\ : Span4Mux_s3_v
    port map (
            O => \N__38447\,
            I => \N__38444\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__38444\,
            I => \N__38440\
        );

    \I__8584\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38437\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__38440\,
            I => data_in_20_4
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__38437\,
            I => data_in_20_4
        );

    \I__8581\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38426\
        );

    \I__8580\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38426\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__38426\,
            I => data_in_19_4
        );

    \I__8578\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38417\
        );

    \I__8577\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38417\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__38417\,
            I => data_in_18_4
        );

    \I__8575\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38408\
        );

    \I__8574\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38408\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__38408\,
            I => data_in_18_2
        );

    \I__8572\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38402\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__38402\,
            I => \N__38399\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__38399\,
            I => \N__38395\
        );

    \I__8569\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__38395\,
            I => \N__38389\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__38392\,
            I => data_in_17_2
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__38389\,
            I => data_in_17_2
        );

    \I__8565\ : InMux
    port map (
            O => \N__38384\,
            I => \N__38381\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__8563\ : Span4Mux_v
    port map (
            O => \N__38378\,
            I => \N__38374\
        );

    \I__8562\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38371\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__38374\,
            I => \N__38368\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38365\
        );

    \I__8559\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38361\
        );

    \I__8558\ : Span12Mux_v
    port map (
            O => \N__38365\,
            I => \N__38358\
        );

    \I__8557\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38355\
        );

    \I__8556\ : Odrv4
    port map (
            O => \N__38361\,
            I => data_in_8_4
        );

    \I__8555\ : Odrv12
    port map (
            O => \N__38358\,
            I => data_in_8_4
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__38355\,
            I => data_in_8_4
        );

    \I__8553\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38343\
        );

    \I__8552\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38338\
        );

    \I__8551\ : InMux
    port map (
            O => \N__38346\,
            I => \N__38338\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__38343\,
            I => \N__38335\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__38338\,
            I => data_in_9_4
        );

    \I__8548\ : Odrv12
    port map (
            O => \N__38335\,
            I => data_in_9_4
        );

    \I__8547\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__38327\,
            I => \N__38322\
        );

    \I__8545\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38317\
        );

    \I__8544\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38317\
        );

    \I__8543\ : Span4Mux_h
    port map (
            O => \N__38322\,
            I => \N__38314\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__38317\,
            I => data_in_10_4
        );

    \I__8541\ : Odrv4
    port map (
            O => \N__38314\,
            I => data_in_10_4
        );

    \I__8540\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38303\
        );

    \I__8539\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38303\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__38303\,
            I => data_in_11_4
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__38300\,
            I => \c0.rx.n18000_cascade_\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__38297\,
            I => \N__38294\
        );

    \I__8535\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__8533\ : Span4Mux_h
    port map (
            O => \N__38288\,
            I => \N__38285\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__38285\,
            I => \c0.rx.n18594\
        );

    \I__8531\ : CascadeMux
    port map (
            O => \N__38282\,
            I => \N__38278\
        );

    \I__8530\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38275\
        );

    \I__8529\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38272\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__38275\,
            I => rand_setpoint_27
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__38272\,
            I => rand_setpoint_27
        );

    \I__8526\ : CascadeMux
    port map (
            O => \N__38267\,
            I => \c0.n17966_cascade_\
        );

    \I__8525\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38260\
        );

    \I__8524\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38257\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__38260\,
            I => rand_setpoint_29
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__38257\,
            I => rand_setpoint_29
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__38252\,
            I => \c0.n17970_cascade_\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__38249\,
            I => \N__38245\
        );

    \I__8519\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38242\
        );

    \I__8518\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38239\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__38242\,
            I => rand_setpoint_24
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__38239\,
            I => rand_setpoint_24
        );

    \I__8515\ : CascadeMux
    port map (
            O => \N__38234\,
            I => \c0.n17957_cascade_\
        );

    \I__8514\ : CascadeMux
    port map (
            O => \N__38231\,
            I => \N__38228\
        );

    \I__8513\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38224\
        );

    \I__8512\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38221\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__38224\,
            I => rand_setpoint_22
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__38221\,
            I => rand_setpoint_22
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__38216\,
            I => \N__38212\
        );

    \I__8508\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38209\
        );

    \I__8507\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38206\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__38209\,
            I => rand_setpoint_4
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__38206\,
            I => rand_setpoint_4
        );

    \I__8504\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38195\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38195\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__38195\,
            I => data_in_15_6
        );

    \I__8501\ : CascadeMux
    port map (
            O => \N__38192\,
            I => \N__38188\
        );

    \I__8500\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8499\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38182\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__38185\,
            I => rand_setpoint_11
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__38182\,
            I => rand_setpoint_11
        );

    \I__8496\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38173\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__38176\,
            I => \N__38170\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__38173\,
            I => \N__38167\
        );

    \I__8493\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38164\
        );

    \I__8492\ : Odrv4
    port map (
            O => \N__38167\,
            I => rand_setpoint_25
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__38164\,
            I => rand_setpoint_25
        );

    \I__8490\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38156\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__38156\,
            I => \N__38152\
        );

    \I__8488\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38149\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__38152\,
            I => \N__38146\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__38149\,
            I => rand_setpoint_30
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__38146\,
            I => rand_setpoint_30
        );

    \I__8484\ : InMux
    port map (
            O => \N__38141\,
            I => \N__38137\
        );

    \I__8483\ : InMux
    port map (
            O => \N__38140\,
            I => \N__38134\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__38137\,
            I => \N__38131\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__38134\,
            I => rand_setpoint_31
        );

    \I__8480\ : Odrv4
    port map (
            O => \N__38131\,
            I => rand_setpoint_31
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__38126\,
            I => \N__38122\
        );

    \I__8478\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38119\
        );

    \I__8477\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38116\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__38119\,
            I => rand_setpoint_10
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38116\,
            I => rand_setpoint_10
        );

    \I__8474\ : InMux
    port map (
            O => \N__38111\,
            I => \N__38107\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__38110\,
            I => \N__38103\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__38107\,
            I => \N__38097\
        );

    \I__8471\ : CascadeMux
    port map (
            O => \N__38106\,
            I => \N__38093\
        );

    \I__8470\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38090\
        );

    \I__8469\ : InMux
    port map (
            O => \N__38102\,
            I => \N__38087\
        );

    \I__8468\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38084\
        );

    \I__8467\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38081\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__38097\,
            I => \N__38078\
        );

    \I__8465\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38073\
        );

    \I__8464\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38073\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__38090\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38087\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__38084\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__38081\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8459\ : Odrv4
    port map (
            O => \N__38078\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__38073\,
            I => \r_Clock_Count_5_adj_2619\
        );

    \I__8457\ : InMux
    port map (
            O => \N__38060\,
            I => \N__38057\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__38057\,
            I => \N__38051\
        );

    \I__8455\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38046\
        );

    \I__8454\ : InMux
    port map (
            O => \N__38055\,
            I => \N__38043\
        );

    \I__8453\ : InMux
    port map (
            O => \N__38054\,
            I => \N__38040\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__38051\,
            I => \N__38037\
        );

    \I__8451\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38032\
        );

    \I__8450\ : InMux
    port map (
            O => \N__38049\,
            I => \N__38032\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__38046\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__38043\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__38040\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__38037\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__38032\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__38021\,
            I => \N__38017\
        );

    \I__8443\ : CascadeMux
    port map (
            O => \N__38020\,
            I => \N__38014\
        );

    \I__8442\ : InMux
    port map (
            O => \N__38017\,
            I => \N__38011\
        );

    \I__8441\ : InMux
    port map (
            O => \N__38014\,
            I => \N__38008\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__38011\,
            I => \N__38005\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__38008\,
            I => \c0.rx.n97\
        );

    \I__8438\ : Odrv12
    port map (
            O => \N__38005\,
            I => \c0.rx.n97\
        );

    \I__8437\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37994\
        );

    \I__8436\ : InMux
    port map (
            O => \N__37999\,
            I => \N__37989\
        );

    \I__8435\ : InMux
    port map (
            O => \N__37998\,
            I => \N__37986\
        );

    \I__8434\ : InMux
    port map (
            O => \N__37997\,
            I => \N__37983\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__37994\,
            I => \N__37980\
        );

    \I__8432\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37975\
        );

    \I__8431\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37975\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__37989\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__37986\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__37983\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__8427\ : Odrv12
    port map (
            O => \N__37980\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__37975\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__8425\ : CascadeMux
    port map (
            O => \N__37964\,
            I => \c0.rx.r_SM_Main_2_N_2380_2_cascade_\
        );

    \I__8424\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37958\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__37958\,
            I => \c0.n18498\
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__37955\,
            I => \c0.n2_adj_2487_cascade_\
        );

    \I__8421\ : InMux
    port map (
            O => \N__37952\,
            I => \N__37949\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__37949\,
            I => n4_adj_2649
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__37946\,
            I => \N__37942\
        );

    \I__8418\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37938\
        );

    \I__8417\ : InMux
    port map (
            O => \N__37942\,
            I => \N__37933\
        );

    \I__8416\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37933\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37930\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__37933\,
            I => \N__37927\
        );

    \I__8413\ : Odrv12
    port map (
            O => \N__37930\,
            I => n8562
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__37927\,
            I => n8562
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__37922\,
            I => \n4_adj_2649_cascade_\
        );

    \I__8410\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37911\
        );

    \I__8409\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37902\
        );

    \I__8408\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37902\
        );

    \I__8407\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37902\
        );

    \I__8406\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37899\
        );

    \I__8405\ : InMux
    port map (
            O => \N__37914\,
            I => \N__37896\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__37911\,
            I => \N__37891\
        );

    \I__8403\ : InMux
    port map (
            O => \N__37910\,
            I => \N__37888\
        );

    \I__8402\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37885\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37882\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__37899\,
            I => \N__37877\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__37896\,
            I => \N__37877\
        );

    \I__8398\ : CascadeMux
    port map (
            O => \N__37895\,
            I => \N__37873\
        );

    \I__8397\ : InMux
    port map (
            O => \N__37894\,
            I => \N__37870\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__37891\,
            I => \N__37867\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37862\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37862\
        );

    \I__8393\ : Span4Mux_h
    port map (
            O => \N__37882\,
            I => \N__37859\
        );

    \I__8392\ : Span4Mux_h
    port map (
            O => \N__37877\,
            I => \N__37856\
        );

    \I__8391\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37851\
        );

    \I__8390\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37851\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__37870\,
            I => \r_Rx_Data\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__37867\,
            I => \r_Rx_Data\
        );

    \I__8387\ : Odrv12
    port map (
            O => \N__37862\,
            I => \r_Rx_Data\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__37859\,
            I => \r_Rx_Data\
        );

    \I__8385\ : Odrv4
    port map (
            O => \N__37856\,
            I => \r_Rx_Data\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__37851\,
            I => \r_Rx_Data\
        );

    \I__8383\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__37835\,
            I => \N__37831\
        );

    \I__8381\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37828\
        );

    \I__8380\ : Odrv4
    port map (
            O => \N__37831\,
            I => rx_data_0
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__37828\,
            I => rx_data_0
        );

    \I__8378\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37820\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__37820\,
            I => \N__37816\
        );

    \I__8376\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37813\
        );

    \I__8375\ : Odrv12
    port map (
            O => \N__37816\,
            I => data_in_20_0
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__37813\,
            I => data_in_20_0
        );

    \I__8373\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37805\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__37805\,
            I => \N__37801\
        );

    \I__8371\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37798\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__37801\,
            I => data_in_17_6
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__37798\,
            I => data_in_17_6
        );

    \I__8368\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37787\
        );

    \I__8367\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37787\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__37787\,
            I => data_in_16_6
        );

    \I__8365\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37781\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__37781\,
            I => \N__37778\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__37778\,
            I => \c0.n6_adj_2448\
        );

    \I__8362\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37771\
        );

    \I__8361\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37768\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__37771\,
            I => data_in_19_6
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__37768\,
            I => data_in_19_6
        );

    \I__8358\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37757\
        );

    \I__8357\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37757\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__37757\,
            I => data_in_18_6
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__37754\,
            I => \N__37750\
        );

    \I__8354\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37747\
        );

    \I__8353\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37744\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__37747\,
            I => rx_data_1
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__37744\,
            I => rx_data_1
        );

    \I__8350\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37735\
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__37738\,
            I => \N__37732\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__37735\,
            I => \N__37729\
        );

    \I__8347\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37726\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__37729\,
            I => rand_setpoint_2
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__37726\,
            I => rand_setpoint_2
        );

    \I__8344\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37718\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__37718\,
            I => \N__37714\
        );

    \I__8342\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37711\
        );

    \I__8341\ : Odrv12
    port map (
            O => \N__37714\,
            I => data_in_19_5
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__37711\,
            I => data_in_19_5
        );

    \I__8339\ : InMux
    port map (
            O => \N__37706\,
            I => \N__37703\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__37703\,
            I => \N__37699\
        );

    \I__8337\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37696\
        );

    \I__8336\ : Odrv4
    port map (
            O => \N__37699\,
            I => rx_data_5
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__37696\,
            I => rx_data_5
        );

    \I__8334\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37685\
        );

    \I__8333\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37685\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__37685\,
            I => data_in_20_5
        );

    \I__8331\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37679\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__37679\,
            I => \N__37676\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__37676\,
            I => \c0.n17911\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__8327\ : InMux
    port map (
            O => \N__37670\,
            I => \N__37667\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__37667\,
            I => \c0.n5_adj_2488\
        );

    \I__8325\ : CascadeMux
    port map (
            O => \N__37664\,
            I => \c0.n17556_cascade_\
        );

    \I__8324\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37657\
        );

    \I__8323\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37653\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__37657\,
            I => \N__37649\
        );

    \I__8321\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37645\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__37653\,
            I => \N__37642\
        );

    \I__8319\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37639\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__37649\,
            I => \N__37636\
        );

    \I__8317\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37633\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__37645\,
            I => \N__37630\
        );

    \I__8315\ : Sp12to4
    port map (
            O => \N__37642\,
            I => \N__37625\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__37639\,
            I => \N__37625\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__37636\,
            I => data_in_1_4
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__37633\,
            I => data_in_1_4
        );

    \I__8311\ : Odrv12
    port map (
            O => \N__37630\,
            I => data_in_1_4
        );

    \I__8310\ : Odrv12
    port map (
            O => \N__37625\,
            I => data_in_1_4
        );

    \I__8309\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37613\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__37613\,
            I => \N__37609\
        );

    \I__8307\ : CascadeMux
    port map (
            O => \N__37612\,
            I => \N__37605\
        );

    \I__8306\ : Span4Mux_v
    port map (
            O => \N__37609\,
            I => \N__37601\
        );

    \I__8305\ : InMux
    port map (
            O => \N__37608\,
            I => \N__37598\
        );

    \I__8304\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37595\
        );

    \I__8303\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37592\
        );

    \I__8302\ : Span4Mux_h
    port map (
            O => \N__37601\,
            I => \N__37589\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__37598\,
            I => \N__37586\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37595\,
            I => \N__37583\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__37592\,
            I => data_in_0_5
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__37589\,
            I => data_in_0_5
        );

    \I__8297\ : Odrv12
    port map (
            O => \N__37586\,
            I => data_in_0_5
        );

    \I__8296\ : Odrv12
    port map (
            O => \N__37583\,
            I => data_in_0_5
        );

    \I__8295\ : CascadeMux
    port map (
            O => \N__37574\,
            I => \N__37570\
        );

    \I__8294\ : InMux
    port map (
            O => \N__37573\,
            I => \N__37567\
        );

    \I__8293\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37563\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37560\
        );

    \I__8291\ : InMux
    port map (
            O => \N__37566\,
            I => \N__37557\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__37563\,
            I => \N__37554\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__37560\,
            I => \N__37547\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37547\
        );

    \I__8287\ : Span4Mux_h
    port map (
            O => \N__37554\,
            I => \N__37544\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__37553\,
            I => \N__37541\
        );

    \I__8285\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37538\
        );

    \I__8284\ : Span4Mux_h
    port map (
            O => \N__37547\,
            I => \N__37533\
        );

    \I__8283\ : Span4Mux_v
    port map (
            O => \N__37544\,
            I => \N__37533\
        );

    \I__8282\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37530\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__37538\,
            I => data_in_2_3
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__37533\,
            I => data_in_2_3
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__37530\,
            I => data_in_2_3
        );

    \I__8278\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__37520\,
            I => \N__37515\
        );

    \I__8276\ : InMux
    port map (
            O => \N__37519\,
            I => \N__37512\
        );

    \I__8275\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37509\
        );

    \I__8274\ : Span4Mux_v
    port map (
            O => \N__37515\,
            I => \N__37504\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__37512\,
            I => \N__37501\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__37509\,
            I => \N__37498\
        );

    \I__8271\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37495\
        );

    \I__8270\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37492\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__37504\,
            I => \N__37489\
        );

    \I__8268\ : Span4Mux_v
    port map (
            O => \N__37501\,
            I => \N__37486\
        );

    \I__8267\ : Span12Mux_s6_h
    port map (
            O => \N__37498\,
            I => \N__37481\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__37495\,
            I => \N__37481\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__37492\,
            I => data_in_3_2
        );

    \I__8264\ : Odrv4
    port map (
            O => \N__37489\,
            I => data_in_3_2
        );

    \I__8263\ : Odrv4
    port map (
            O => \N__37486\,
            I => data_in_3_2
        );

    \I__8262\ : Odrv12
    port map (
            O => \N__37481\,
            I => data_in_3_2
        );

    \I__8261\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__8259\ : Span4Mux_h
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__8258\ : Span4Mux_h
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__37460\,
            I => \c0.n16_adj_2513\
        );

    \I__8256\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37450\
        );

    \I__8254\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37447\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__37450\,
            I => data_in_18_0
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__37447\,
            I => data_in_18_0
        );

    \I__8251\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37437\
        );

    \I__8250\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37434\
        );

    \I__8249\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37431\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37428\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37425\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37431\,
            I => n9796
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__37428\,
            I => n9796
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__37425\,
            I => n9796
        );

    \I__8243\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37414\
        );

    \I__8242\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37411\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__37414\,
            I => \N__37408\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__37411\,
            I => \r_Tx_Data_7\
        );

    \I__8239\ : Odrv12
    port map (
            O => \N__37408\,
            I => \r_Tx_Data_7\
        );

    \I__8238\ : CascadeMux
    port map (
            O => \N__37403\,
            I => \N__37399\
        );

    \I__8237\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37390\
        );

    \I__8236\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37390\
        );

    \I__8235\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37385\
        );

    \I__8234\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37385\
        );

    \I__8233\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37382\
        );

    \I__8232\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37379\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__37390\,
            I => \N__37376\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__37385\,
            I => \N__37373\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__37382\,
            I => \r_Bit_Index_2\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__37379\,
            I => \r_Bit_Index_2\
        );

    \I__8227\ : Odrv12
    port map (
            O => \N__37376\,
            I => \r_Bit_Index_2\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__37373\,
            I => \r_Bit_Index_2\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37364\,
            I => \N__37359\
        );

    \I__8224\ : InMux
    port map (
            O => \N__37363\,
            I => \N__37354\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37354\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__37359\,
            I => \N__37351\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37354\,
            I => n12_adj_2618
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__37351\,
            I => n12_adj_2618
        );

    \I__8219\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__37343\,
            I => \N__37340\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__37337\,
            I => n22
        );

    \I__8215\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__8213\ : Odrv12
    port map (
            O => \N__37328\,
            I => n17950
        );

    \I__8212\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37322\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__37322\,
            I => \N__37316\
        );

    \I__8210\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37312\
        );

    \I__8209\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37309\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37306\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__37316\,
            I => \N__37303\
        );

    \I__8206\ : InMux
    port map (
            O => \N__37315\,
            I => \N__37300\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__37312\,
            I => \N__37295\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__37309\,
            I => \N__37295\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__37306\,
            I => \r_Clock_Count_8\
        );

    \I__8202\ : Odrv4
    port map (
            O => \N__37303\,
            I => \r_Clock_Count_8\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__37300\,
            I => \r_Clock_Count_8\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__37295\,
            I => \r_Clock_Count_8\
        );

    \I__8199\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__37283\,
            I => n17767
        );

    \I__8197\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37277\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__37277\,
            I => \c0.tx.n17\
        );

    \I__8195\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37268\
        );

    \I__8194\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37268\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__37268\,
            I => \r_Tx_Data_2\
        );

    \I__8192\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37262\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__37262\,
            I => \N__37258\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__37261\,
            I => \N__37255\
        );

    \I__8189\ : Span4Mux_h
    port map (
            O => \N__37258\,
            I => \N__37249\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37246\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37241\
        );

    \I__8186\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37241\
        );

    \I__8185\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37238\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__37249\,
            I => \r_Clock_Count_6\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__37246\,
            I => \r_Clock_Count_6\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__37241\,
            I => \r_Clock_Count_6\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__37238\,
            I => \r_Clock_Count_6\
        );

    \I__8180\ : InMux
    port map (
            O => \N__37229\,
            I => \N__37226\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__37226\,
            I => \N__37223\
        );

    \I__8178\ : Span4Mux_v
    port map (
            O => \N__37223\,
            I => \N__37219\
        );

    \I__8177\ : InMux
    port map (
            O => \N__37222\,
            I => \N__37216\
        );

    \I__8176\ : Span4Mux_h
    port map (
            O => \N__37219\,
            I => \N__37210\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__37216\,
            I => \N__37210\
        );

    \I__8174\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37206\
        );

    \I__8173\ : Span4Mux_v
    port map (
            O => \N__37210\,
            I => \N__37203\
        );

    \I__8172\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37200\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__37206\,
            I => \N__37192\
        );

    \I__8170\ : Sp12to4
    port map (
            O => \N__37203\,
            I => \N__37192\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37192\
        );

    \I__8168\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37189\
        );

    \I__8167\ : Span12Mux_h
    port map (
            O => \N__37192\,
            I => \N__37186\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__37189\,
            I => \r_Clock_Count_7\
        );

    \I__8165\ : Odrv12
    port map (
            O => \N__37186\,
            I => \r_Clock_Count_7\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__37181\,
            I => \n1_cascade_\
        );

    \I__8163\ : CascadeMux
    port map (
            O => \N__37178\,
            I => \n3_adj_2650_cascade_\
        );

    \I__8162\ : IoInMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__8160\ : IoSpan4Mux
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__8159\ : Span4Mux_s0_v
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__8158\ : Span4Mux_h
    port map (
            O => \N__37163\,
            I => \N__37159\
        );

    \I__8157\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37156\
        );

    \I__8156\ : Span4Mux_s0_v
    port map (
            O => \N__37159\,
            I => \N__37151\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__37156\,
            I => \N__37151\
        );

    \I__8154\ : Span4Mux_v
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__8152\ : Span4Mux_h
    port map (
            O => \N__37145\,
            I => \N__37141\
        );

    \I__8151\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37138\
        );

    \I__8150\ : Odrv4
    port map (
            O => \N__37141\,
            I => tx_o_adj_2584
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__37138\,
            I => tx_o_adj_2584
        );

    \I__8148\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37129\
        );

    \I__8147\ : InMux
    port map (
            O => \N__37132\,
            I => \N__37126\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__37129\,
            I => data_in_18_7
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__37126\,
            I => data_in_18_7
        );

    \I__8144\ : InMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__37118\,
            I => \N__37114\
        );

    \I__8142\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37111\
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__37114\,
            I => rx_data_7
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__37111\,
            I => rx_data_7
        );

    \I__8139\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37099\
        );

    \I__8137\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37096\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__37099\,
            I => data_in_16_3
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__37096\,
            I => data_in_16_3
        );

    \I__8134\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37084\
        );

    \I__8132\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37081\
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__37084\,
            I => data_in_15_3
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__37081\,
            I => data_in_15_3
        );

    \I__8129\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37070\
        );

    \I__8128\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37070\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__37070\,
            I => data_in_20_7
        );

    \I__8126\ : InMux
    port map (
            O => \N__37067\,
            I => \N__37063\
        );

    \I__8125\ : InMux
    port map (
            O => \N__37066\,
            I => \N__37060\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__37063\,
            I => data_in_19_7
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__37060\,
            I => data_in_19_7
        );

    \I__8122\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__37052\,
            I => n12123
        );

    \I__8120\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__37046\,
            I => n7080
        );

    \I__8118\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37039\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37036\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__37039\,
            I => \N__37033\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37036\,
            I => \N__37029\
        );

    \I__8114\ : Span4Mux_h
    port map (
            O => \N__37033\,
            I => \N__37026\
        );

    \I__8113\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37023\
        );

    \I__8112\ : Odrv12
    port map (
            O => \N__37029\,
            I => data_in_8_1
        );

    \I__8111\ : Odrv4
    port map (
            O => \N__37026\,
            I => data_in_8_1
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__37023\,
            I => data_in_8_1
        );

    \I__8109\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37012\
        );

    \I__8108\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37009\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__37012\,
            I => \N__37005\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__37009\,
            I => \N__37002\
        );

    \I__8105\ : InMux
    port map (
            O => \N__37008\,
            I => \N__36999\
        );

    \I__8104\ : Span4Mux_h
    port map (
            O => \N__37005\,
            I => \N__36996\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__37002\,
            I => \c0.data_in_7_1\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__36999\,
            I => \c0.data_in_7_1\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__36996\,
            I => \c0.data_in_7_1\
        );

    \I__8100\ : CascadeMux
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__8099\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36979\
        );

    \I__8097\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36975\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__36979\,
            I => \N__36972\
        );

    \I__8095\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36969\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__36975\,
            I => data_in_10_3
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__36972\,
            I => data_in_10_3
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__36969\,
            I => data_in_10_3
        );

    \I__8091\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36958\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__36961\,
            I => \N__36955\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__36958\,
            I => \N__36952\
        );

    \I__8088\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36949\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__36952\,
            I => \N__36944\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__36949\,
            I => \N__36941\
        );

    \I__8085\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36938\
        );

    \I__8084\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36935\
        );

    \I__8083\ : Span4Mux_h
    port map (
            O => \N__36944\,
            I => \N__36930\
        );

    \I__8082\ : Span4Mux_v
    port map (
            O => \N__36941\,
            I => \N__36930\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__36938\,
            I => data_in_6_7
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__36935\,
            I => data_in_6_7
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__36930\,
            I => data_in_6_7
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__36923\,
            I => \N__36920\
        );

    \I__8077\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36917\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__36917\,
            I => \N__36913\
        );

    \I__8075\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36909\
        );

    \I__8074\ : Span4Mux_v
    port map (
            O => \N__36913\,
            I => \N__36906\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__36912\,
            I => \N__36903\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__36909\,
            I => \N__36899\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__36906\,
            I => \N__36896\
        );

    \I__8070\ : InMux
    port map (
            O => \N__36903\,
            I => \N__36893\
        );

    \I__8069\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36890\
        );

    \I__8068\ : Span4Mux_h
    port map (
            O => \N__36899\,
            I => \N__36887\
        );

    \I__8067\ : Span4Mux_h
    port map (
            O => \N__36896\,
            I => \N__36884\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__36893\,
            I => \N__36881\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__36890\,
            I => data_in_5_7
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__36887\,
            I => data_in_5_7
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__36884\,
            I => data_in_5_7
        );

    \I__8062\ : Odrv12
    port map (
            O => \N__36881\,
            I => data_in_5_7
        );

    \I__8061\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36868\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__36871\,
            I => \N__36865\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36862\
        );

    \I__8058\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36859\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__36862\,
            I => \N__36852\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__36859\,
            I => \N__36852\
        );

    \I__8055\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36849\
        );

    \I__8054\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36846\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__36852\,
            I => \N__36843\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__36849\,
            I => \c0.data_in_frame_10_1\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__36846\,
            I => \c0.data_in_frame_10_1\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__36843\,
            I => \c0.data_in_frame_10_1\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__36836\,
            I => \N__36833\
        );

    \I__8048\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36828\
        );

    \I__8047\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36825\
        );

    \I__8046\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36822\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36819\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__36825\,
            I => \N__36814\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__36822\,
            I => \N__36814\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__36819\,
            I => \N__36811\
        );

    \I__8041\ : Odrv12
    port map (
            O => \N__36814\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__36811\,
            I => \c0.data_in_frame_10_3\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__8038\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36800\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__8036\ : Span4Mux_h
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__8035\ : Span4Mux_h
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__8033\ : Odrv4
    port map (
            O => \N__36788\,
            I => \c0.n6\
        );

    \I__8032\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__36779\,
            I => \N__36775\
        );

    \I__8029\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36772\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__36775\,
            I => data_in_11_0
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__36772\,
            I => data_in_11_0
        );

    \I__8026\ : InMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__36764\,
            I => n7086
        );

    \I__8024\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__8022\ : Span4Mux_h
    port map (
            O => \N__36755\,
            I => \N__36751\
        );

    \I__8021\ : InMux
    port map (
            O => \N__36754\,
            I => \N__36748\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__36751\,
            I => data_in_15_1
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__36748\,
            I => data_in_15_1
        );

    \I__8018\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36736\
        );

    \I__8017\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36736\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__36741\,
            I => \N__36733\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__36736\,
            I => \N__36730\
        );

    \I__8014\ : InMux
    port map (
            O => \N__36733\,
            I => \N__36726\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__36730\,
            I => \N__36723\
        );

    \I__8012\ : InMux
    port map (
            O => \N__36729\,
            I => \N__36720\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__36726\,
            I => \N__36717\
        );

    \I__8010\ : IoSpan4Mux
    port map (
            O => \N__36723\,
            I => \N__36714\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36711\
        );

    \I__8008\ : Span4Mux_h
    port map (
            O => \N__36717\,
            I => \N__36708\
        );

    \I__8007\ : IoSpan4Mux
    port map (
            O => \N__36714\,
            I => \N__36705\
        );

    \I__8006\ : Span12Mux_h
    port map (
            O => \N__36711\,
            I => \N__36702\
        );

    \I__8005\ : Span4Mux_s2_h
    port map (
            O => \N__36708\,
            I => \N__36699\
        );

    \I__8004\ : Odrv4
    port map (
            O => \N__36705\,
            I => \c0.data_in_frame_9_1\
        );

    \I__8003\ : Odrv12
    port map (
            O => \N__36702\,
            I => \c0.data_in_frame_9_1\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__36699\,
            I => \c0.data_in_frame_9_1\
        );

    \I__8001\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36687\
        );

    \I__8000\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36682\
        );

    \I__7999\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36679\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__36687\,
            I => \N__36676\
        );

    \I__7997\ : InMux
    port map (
            O => \N__36686\,
            I => \N__36673\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__36685\,
            I => \N__36670\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__36682\,
            I => \N__36667\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36664\
        );

    \I__7993\ : Span4Mux_h
    port map (
            O => \N__36676\,
            I => \N__36659\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36659\
        );

    \I__7991\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36656\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__36667\,
            I => \N__36653\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__36664\,
            I => \N__36650\
        );

    \I__7988\ : Span4Mux_v
    port map (
            O => \N__36659\,
            I => \N__36645\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36645\
        );

    \I__7986\ : Span4Mux_h
    port map (
            O => \N__36653\,
            I => \N__36642\
        );

    \I__7985\ : Span4Mux_h
    port map (
            O => \N__36650\,
            I => \N__36637\
        );

    \I__7984\ : Span4Mux_v
    port map (
            O => \N__36645\,
            I => \N__36637\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__36642\,
            I => \c0.data_in_frame_10_7\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__36637\,
            I => \c0.data_in_frame_10_7\
        );

    \I__7981\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36626\
        );

    \I__7980\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36626\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__36626\,
            I => \N__36621\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__36625\,
            I => \N__36618\
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__36624\,
            I => \N__36615\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__36621\,
            I => \N__36612\
        );

    \I__7975\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36609\
        );

    \I__7974\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36606\
        );

    \I__7973\ : Span4Mux_v
    port map (
            O => \N__36612\,
            I => \N__36601\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36601\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__36606\,
            I => \N__36598\
        );

    \I__7970\ : Span4Mux_v
    port map (
            O => \N__36601\,
            I => \N__36594\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__36598\,
            I => \N__36591\
        );

    \I__7968\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36588\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__36594\,
            I => \c0.data_in_frame_9_5\
        );

    \I__7966\ : Odrv4
    port map (
            O => \N__36591\,
            I => \c0.data_in_frame_9_5\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__36588\,
            I => \c0.data_in_frame_9_5\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__36581\,
            I => \N__36576\
        );

    \I__7963\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36573\
        );

    \I__7962\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36568\
        );

    \I__7961\ : InMux
    port map (
            O => \N__36576\,
            I => \N__36568\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__36573\,
            I => \N__36565\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__36568\,
            I => \N__36562\
        );

    \I__7958\ : Odrv12
    port map (
            O => \N__36565\,
            I => \c0.data_in_frame_9_3\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__36562\,
            I => \c0.data_in_frame_9_3\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__36557\,
            I => \N__36553\
        );

    \I__7955\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36548\
        );

    \I__7954\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36548\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36544\
        );

    \I__7952\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36541\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__36544\,
            I => \N__36538\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__36541\,
            I => \N__36535\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__36538\,
            I => \N__36532\
        );

    \I__7948\ : Span12Mux_s9_h
    port map (
            O => \N__36535\,
            I => \N__36529\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__36532\,
            I => \c0.n8989\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__36529\,
            I => \c0.n8989\
        );

    \I__7945\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36520\
        );

    \I__7944\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36517\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__36520\,
            I => \N__36513\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__36517\,
            I => \N__36510\
        );

    \I__7941\ : InMux
    port map (
            O => \N__36516\,
            I => \N__36507\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__36513\,
            I => \N__36504\
        );

    \I__7939\ : Odrv4
    port map (
            O => \N__36510\,
            I => data_in_10_2
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__36507\,
            I => data_in_10_2
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__36504\,
            I => data_in_10_2
        );

    \I__7936\ : InMux
    port map (
            O => \N__36497\,
            I => \N__36494\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__36494\,
            I => \N__36489\
        );

    \I__7934\ : InMux
    port map (
            O => \N__36493\,
            I => \N__36486\
        );

    \I__7933\ : InMux
    port map (
            O => \N__36492\,
            I => \N__36483\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__36489\,
            I => \N__36480\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36477\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__36483\,
            I => data_in_9_2
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__36480\,
            I => data_in_9_2
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__36477\,
            I => data_in_9_2
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__7926\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__36464\,
            I => \N__36460\
        );

    \I__7924\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36455\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__36460\,
            I => \N__36452\
        );

    \I__7922\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36449\
        );

    \I__7921\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36446\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__36455\,
            I => \N__36443\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__36452\,
            I => \N__36438\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__36449\,
            I => \N__36438\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__36446\,
            I => \N__36434\
        );

    \I__7916\ : Span12Mux_s4_h
    port map (
            O => \N__36443\,
            I => \N__36431\
        );

    \I__7915\ : Span4Mux_h
    port map (
            O => \N__36438\,
            I => \N__36428\
        );

    \I__7914\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36425\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__36434\,
            I => \N__36422\
        );

    \I__7912\ : Odrv12
    port map (
            O => \N__36431\,
            I => rand_data_28
        );

    \I__7911\ : Odrv4
    port map (
            O => \N__36428\,
            I => rand_data_28
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__36425\,
            I => rand_data_28
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__36422\,
            I => rand_data_28
        );

    \I__7908\ : InMux
    port map (
            O => \N__36413\,
            I => n16439
        );

    \I__7907\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36403\
        );

    \I__7906\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36403\
        );

    \I__7905\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36400\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__36403\,
            I => \N__36396\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__36400\,
            I => \N__36393\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__36399\,
            I => \N__36390\
        );

    \I__7901\ : Span4Mux_v
    port map (
            O => \N__36396\,
            I => \N__36387\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__36393\,
            I => \N__36384\
        );

    \I__7899\ : InMux
    port map (
            O => \N__36390\,
            I => \N__36380\
        );

    \I__7898\ : Span4Mux_h
    port map (
            O => \N__36387\,
            I => \N__36377\
        );

    \I__7897\ : Span4Mux_v
    port map (
            O => \N__36384\,
            I => \N__36374\
        );

    \I__7896\ : InMux
    port map (
            O => \N__36383\,
            I => \N__36371\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__36380\,
            I => \N__36368\
        );

    \I__7894\ : Odrv4
    port map (
            O => \N__36377\,
            I => rand_data_29
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__36374\,
            I => rand_data_29
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__36371\,
            I => rand_data_29
        );

    \I__7891\ : Odrv12
    port map (
            O => \N__36368\,
            I => rand_data_29
        );

    \I__7890\ : InMux
    port map (
            O => \N__36359\,
            I => n16440
        );

    \I__7889\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36348\
        );

    \I__7888\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36348\
        );

    \I__7887\ : InMux
    port map (
            O => \N__36354\,
            I => \N__36345\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__36353\,
            I => \N__36342\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__36348\,
            I => \N__36339\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__36345\,
            I => \N__36336\
        );

    \I__7883\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36332\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__36339\,
            I => \N__36329\
        );

    \I__7881\ : Span12Mux_h
    port map (
            O => \N__36336\,
            I => \N__36326\
        );

    \I__7880\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36323\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__36332\,
            I => \N__36320\
        );

    \I__7878\ : Odrv4
    port map (
            O => \N__36329\,
            I => rand_data_30
        );

    \I__7877\ : Odrv12
    port map (
            O => \N__36326\,
            I => rand_data_30
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__36323\,
            I => rand_data_30
        );

    \I__7875\ : Odrv12
    port map (
            O => \N__36320\,
            I => rand_data_30
        );

    \I__7874\ : InMux
    port map (
            O => \N__36311\,
            I => n16441
        );

    \I__7873\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36301\
        );

    \I__7872\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36301\
        );

    \I__7871\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36298\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__36301\,
            I => \N__36294\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__36298\,
            I => \N__36291\
        );

    \I__7868\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36288\
        );

    \I__7867\ : Span4Mux_v
    port map (
            O => \N__36294\,
            I => \N__36284\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__36291\,
            I => \N__36281\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__36288\,
            I => \N__36278\
        );

    \I__7864\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36275\
        );

    \I__7863\ : Span4Mux_v
    port map (
            O => \N__36284\,
            I => \N__36268\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__36281\,
            I => \N__36268\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__36278\,
            I => \N__36268\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__36275\,
            I => rand_data_31
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__36268\,
            I => rand_data_31
        );

    \I__7858\ : InMux
    port map (
            O => \N__36263\,
            I => n16442
        );

    \I__7857\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36256\
        );

    \I__7856\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36253\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36250\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7852\ : Span4Mux_h
    port map (
            O => \N__36247\,
            I => \N__36239\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__36244\,
            I => \N__36236\
        );

    \I__7850\ : InMux
    port map (
            O => \N__36243\,
            I => \N__36231\
        );

    \I__7849\ : InMux
    port map (
            O => \N__36242\,
            I => \N__36231\
        );

    \I__7848\ : Odrv4
    port map (
            O => \N__36239\,
            I => data_in_1_5
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__36236\,
            I => data_in_1_5
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__36231\,
            I => data_in_1_5
        );

    \I__7845\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36220\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__36223\,
            I => \N__36217\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__36220\,
            I => \N__36214\
        );

    \I__7842\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36211\
        );

    \I__7841\ : Span4Mux_v
    port map (
            O => \N__36214\,
            I => \N__36207\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__36211\,
            I => \N__36204\
        );

    \I__7839\ : InMux
    port map (
            O => \N__36210\,
            I => \N__36201\
        );

    \I__7838\ : Span4Mux_h
    port map (
            O => \N__36207\,
            I => \N__36196\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__36204\,
            I => \N__36196\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__36201\,
            I => data_in_7_5
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__36196\,
            I => data_in_7_5
        );

    \I__7834\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36187\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__36190\,
            I => \N__36184\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__36187\,
            I => \N__36181\
        );

    \I__7831\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__36181\,
            I => \N__36174\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__36178\,
            I => \N__36171\
        );

    \I__7828\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36168\
        );

    \I__7827\ : Span4Mux_h
    port map (
            O => \N__36174\,
            I => \N__36165\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__36171\,
            I => \N__36162\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__36168\,
            I => data_in_6_5
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__36165\,
            I => data_in_6_5
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__36162\,
            I => data_in_6_5
        );

    \I__7822\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36152\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__36152\,
            I => \N__36148\
        );

    \I__7820\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36145\
        );

    \I__7819\ : Span4Mux_s2_h
    port map (
            O => \N__36148\,
            I => \N__36138\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__36138\
        );

    \I__7817\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36135\
        );

    \I__7816\ : InMux
    port map (
            O => \N__36143\,
            I => \N__36132\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__36138\,
            I => \N__36128\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36125\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__36122\
        );

    \I__7812\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36119\
        );

    \I__7811\ : Span4Mux_s1_v
    port map (
            O => \N__36128\,
            I => \N__36114\
        );

    \I__7810\ : Span4Mux_h
    port map (
            O => \N__36125\,
            I => \N__36114\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__36122\,
            I => rand_data_20
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__36119\,
            I => rand_data_20
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__36114\,
            I => rand_data_20
        );

    \I__7806\ : InMux
    port map (
            O => \N__36107\,
            I => n16431
        );

    \I__7805\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36101\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__36101\,
            I => \N__36095\
        );

    \I__7803\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36092\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36089\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__36098\,
            I => \N__36086\
        );

    \I__7800\ : Span4Mux_h
    port map (
            O => \N__36095\,
            I => \N__36083\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__36092\,
            I => \N__36080\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__36089\,
            I => \N__36077\
        );

    \I__7797\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36073\
        );

    \I__7796\ : Span4Mux_v
    port map (
            O => \N__36083\,
            I => \N__36070\
        );

    \I__7795\ : Span4Mux_h
    port map (
            O => \N__36080\,
            I => \N__36067\
        );

    \I__7794\ : Span4Mux_v
    port map (
            O => \N__36077\,
            I => \N__36064\
        );

    \I__7793\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36061\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36058\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__36070\,
            I => rand_data_21
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__36067\,
            I => rand_data_21
        );

    \I__7789\ : Odrv4
    port map (
            O => \N__36064\,
            I => rand_data_21
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__36061\,
            I => rand_data_21
        );

    \I__7787\ : Odrv12
    port map (
            O => \N__36058\,
            I => rand_data_21
        );

    \I__7786\ : InMux
    port map (
            O => \N__36047\,
            I => n16432
        );

    \I__7785\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36035\
        );

    \I__7784\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36035\
        );

    \I__7783\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36035\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__36031\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__7780\ : Sp12to4
    port map (
            O => \N__36031\,
            I => \N__36024\
        );

    \I__7779\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36021\
        );

    \I__7778\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36018\
        );

    \I__7777\ : Span12Mux_v
    port map (
            O => \N__36024\,
            I => \N__36013\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__36013\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__36018\,
            I => rand_data_22
        );

    \I__7774\ : Odrv12
    port map (
            O => \N__36013\,
            I => rand_data_22
        );

    \I__7773\ : InMux
    port map (
            O => \N__36008\,
            I => n16433
        );

    \I__7772\ : InMux
    port map (
            O => \N__36005\,
            I => \N__36000\
        );

    \I__7771\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35995\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35995\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__36000\,
            I => \N__35992\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35988\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__35992\,
            I => \N__35985\
        );

    \I__7766\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35982\
        );

    \I__7765\ : Span4Mux_h
    port map (
            O => \N__35988\,
            I => \N__35979\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__35985\,
            I => \N__35975\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35972\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__35979\,
            I => \N__35969\
        );

    \I__7761\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35966\
        );

    \I__7760\ : Span4Mux_s1_h
    port map (
            O => \N__35975\,
            I => \N__35961\
        );

    \I__7759\ : Span4Mux_h
    port map (
            O => \N__35972\,
            I => \N__35961\
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__35969\,
            I => rand_data_23
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__35966\,
            I => rand_data_23
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__35961\,
            I => rand_data_23
        );

    \I__7755\ : InMux
    port map (
            O => \N__35954\,
            I => n16434
        );

    \I__7754\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35946\
        );

    \I__7753\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35943\
        );

    \I__7752\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35940\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__35946\,
            I => \N__35936\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__35943\,
            I => \N__35933\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__35940\,
            I => \N__35930\
        );

    \I__7748\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35927\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__35936\,
            I => \N__35924\
        );

    \I__7746\ : Span4Mux_h
    port map (
            O => \N__35933\,
            I => \N__35921\
        );

    \I__7745\ : Span4Mux_h
    port map (
            O => \N__35930\,
            I => \N__35917\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35914\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__35924\,
            I => \N__35911\
        );

    \I__7742\ : Span4Mux_v
    port map (
            O => \N__35921\,
            I => \N__35908\
        );

    \I__7741\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35905\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__35917\,
            I => \N__35900\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__35914\,
            I => \N__35900\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__35911\,
            I => rand_data_24
        );

    \I__7737\ : Odrv4
    port map (
            O => \N__35908\,
            I => rand_data_24
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__35905\,
            I => rand_data_24
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__35900\,
            I => rand_data_24
        );

    \I__7734\ : InMux
    port map (
            O => \N__35891\,
            I => \bfn_9_32_0_\
        );

    \I__7733\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35883\
        );

    \I__7732\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35880\
        );

    \I__7731\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35877\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__35883\,
            I => \N__35874\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35871\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35868\
        );

    \I__7727\ : Span4Mux_h
    port map (
            O => \N__35874\,
            I => \N__35864\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__35871\,
            I => \N__35861\
        );

    \I__7725\ : Span4Mux_v
    port map (
            O => \N__35868\,
            I => \N__35857\
        );

    \I__7724\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35854\
        );

    \I__7723\ : Span4Mux_v
    port map (
            O => \N__35864\,
            I => \N__35851\
        );

    \I__7722\ : Span4Mux_v
    port map (
            O => \N__35861\,
            I => \N__35848\
        );

    \I__7721\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35845\
        );

    \I__7720\ : Sp12to4
    port map (
            O => \N__35857\,
            I => \N__35840\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35840\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__35851\,
            I => rand_data_25
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__35848\,
            I => rand_data_25
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__35845\,
            I => rand_data_25
        );

    \I__7715\ : Odrv12
    port map (
            O => \N__35840\,
            I => rand_data_25
        );

    \I__7714\ : InMux
    port map (
            O => \N__35831\,
            I => n16436
        );

    \I__7713\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35825\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35822\
        );

    \I__7711\ : Span4Mux_v
    port map (
            O => \N__35822\,
            I => \N__35818\
        );

    \I__7710\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35815\
        );

    \I__7709\ : Span4Mux_s1_h
    port map (
            O => \N__35818\,
            I => \N__35810\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__35815\,
            I => \N__35810\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__35810\,
            I => \N__35806\
        );

    \I__7706\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35803\
        );

    \I__7705\ : Span4Mux_s1_h
    port map (
            O => \N__35806\,
            I => \N__35797\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__35803\,
            I => \N__35797\
        );

    \I__7703\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35793\
        );

    \I__7702\ : Span4Mux_h
    port map (
            O => \N__35797\,
            I => \N__35790\
        );

    \I__7701\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35787\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__35793\,
            I => \N__35784\
        );

    \I__7699\ : Odrv4
    port map (
            O => \N__35790\,
            I => rand_data_26
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__35787\,
            I => rand_data_26
        );

    \I__7697\ : Odrv12
    port map (
            O => \N__35784\,
            I => rand_data_26
        );

    \I__7696\ : InMux
    port map (
            O => \N__35777\,
            I => n16437
        );

    \I__7695\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35766\
        );

    \I__7693\ : InMux
    port map (
            O => \N__35770\,
            I => \N__35763\
        );

    \I__7692\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35760\
        );

    \I__7691\ : Span4Mux_v
    port map (
            O => \N__35766\,
            I => \N__35756\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__35763\,
            I => \N__35753\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__35760\,
            I => \N__35750\
        );

    \I__7688\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35746\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__35756\,
            I => \N__35743\
        );

    \I__7686\ : Span4Mux_h
    port map (
            O => \N__35753\,
            I => \N__35740\
        );

    \I__7685\ : Span4Mux_h
    port map (
            O => \N__35750\,
            I => \N__35737\
        );

    \I__7684\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35734\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__35746\,
            I => \N__35731\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__35743\,
            I => rand_data_27
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__35740\,
            I => rand_data_27
        );

    \I__7680\ : Odrv4
    port map (
            O => \N__35737\,
            I => rand_data_27
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__35734\,
            I => rand_data_27
        );

    \I__7678\ : Odrv12
    port map (
            O => \N__35731\,
            I => rand_data_27
        );

    \I__7677\ : InMux
    port map (
            O => \N__35720\,
            I => n16438
        );

    \I__7676\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35710\
        );

    \I__7675\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35710\
        );

    \I__7674\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35707\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__35710\,
            I => \N__35701\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__35707\,
            I => \N__35701\
        );

    \I__7671\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35698\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__35701\,
            I => \N__35693\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35693\
        );

    \I__7668\ : Span4Mux_v
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__7667\ : Span4Mux_s1_h
    port map (
            O => \N__35690\,
            I => \N__35686\
        );

    \I__7666\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35682\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__35686\,
            I => \N__35679\
        );

    \I__7664\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35676\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__35682\,
            I => \N__35673\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__35679\,
            I => rand_data_11
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__35676\,
            I => rand_data_11
        );

    \I__7660\ : Odrv12
    port map (
            O => \N__35673\,
            I => rand_data_11
        );

    \I__7659\ : InMux
    port map (
            O => \N__35666\,
            I => n16422
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__35663\,
            I => \N__35659\
        );

    \I__7657\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35654\
        );

    \I__7656\ : InMux
    port map (
            O => \N__35659\,
            I => \N__35651\
        );

    \I__7655\ : InMux
    port map (
            O => \N__35658\,
            I => \N__35648\
        );

    \I__7654\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35644\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__35654\,
            I => \N__35641\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35636\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__35648\,
            I => \N__35636\
        );

    \I__7650\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35633\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__35644\,
            I => \N__35629\
        );

    \I__7648\ : Span4Mux_v
    port map (
            O => \N__35641\,
            I => \N__35626\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__35636\,
            I => \N__35621\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35621\
        );

    \I__7645\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35618\
        );

    \I__7644\ : Span4Mux_h
    port map (
            O => \N__35629\,
            I => \N__35615\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__35626\,
            I => rand_data_12
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__35621\,
            I => rand_data_12
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__35618\,
            I => rand_data_12
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__35615\,
            I => rand_data_12
        );

    \I__7639\ : InMux
    port map (
            O => \N__35606\,
            I => n16423
        );

    \I__7638\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35596\
        );

    \I__7637\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35596\
        );

    \I__7636\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35592\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35589\
        );

    \I__7634\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35586\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__35592\,
            I => \N__35582\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__35589\,
            I => \N__35579\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__35586\,
            I => \N__35576\
        );

    \I__7630\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35573\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__35582\,
            I => \N__35570\
        );

    \I__7628\ : Span4Mux_v
    port map (
            O => \N__35579\,
            I => \N__35567\
        );

    \I__7627\ : Span4Mux_s1_h
    port map (
            O => \N__35576\,
            I => \N__35564\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__35573\,
            I => \N__35560\
        );

    \I__7625\ : Span4Mux_v
    port map (
            O => \N__35570\,
            I => \N__35557\
        );

    \I__7624\ : Span4Mux_s1_h
    port map (
            O => \N__35567\,
            I => \N__35552\
        );

    \I__7623\ : Span4Mux_v
    port map (
            O => \N__35564\,
            I => \N__35552\
        );

    \I__7622\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35549\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__35560\,
            I => \N__35546\
        );

    \I__7620\ : Odrv4
    port map (
            O => \N__35557\,
            I => rand_data_13
        );

    \I__7619\ : Odrv4
    port map (
            O => \N__35552\,
            I => rand_data_13
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__35549\,
            I => rand_data_13
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__35546\,
            I => rand_data_13
        );

    \I__7616\ : InMux
    port map (
            O => \N__35537\,
            I => n16424
        );

    \I__7615\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35529\
        );

    \I__7614\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35524\
        );

    \I__7613\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35524\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__35529\,
            I => \N__35519\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35516\
        );

    \I__7610\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35513\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__35522\,
            I => \N__35510\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__35519\,
            I => \N__35507\
        );

    \I__7607\ : Span4Mux_h
    port map (
            O => \N__35516\,
            I => \N__35504\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__35513\,
            I => \N__35500\
        );

    \I__7605\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35497\
        );

    \I__7604\ : Span4Mux_v
    port map (
            O => \N__35507\,
            I => \N__35492\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__35504\,
            I => \N__35492\
        );

    \I__7602\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35489\
        );

    \I__7601\ : Span12Mux_v
    port map (
            O => \N__35500\,
            I => \N__35484\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35484\
        );

    \I__7599\ : Odrv4
    port map (
            O => \N__35492\,
            I => rand_data_14
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__35489\,
            I => rand_data_14
        );

    \I__7597\ : Odrv12
    port map (
            O => \N__35484\,
            I => rand_data_14
        );

    \I__7596\ : InMux
    port map (
            O => \N__35477\,
            I => n16425
        );

    \I__7595\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35468\
        );

    \I__7593\ : Span4Mux_h
    port map (
            O => \N__35468\,
            I => \N__35464\
        );

    \I__7592\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35461\
        );

    \I__7591\ : Span4Mux_v
    port map (
            O => \N__35464\,
            I => \N__35455\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__35461\,
            I => \N__35452\
        );

    \I__7589\ : InMux
    port map (
            O => \N__35460\,
            I => \N__35449\
        );

    \I__7588\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35446\
        );

    \I__7587\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35443\
        );

    \I__7586\ : Span4Mux_h
    port map (
            O => \N__35455\,
            I => \N__35438\
        );

    \I__7585\ : Span4Mux_h
    port map (
            O => \N__35452\,
            I => \N__35438\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__35449\,
            I => \N__35432\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35432\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__35443\,
            I => \N__35429\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__35438\,
            I => \N__35426\
        );

    \I__7580\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35423\
        );

    \I__7579\ : Span4Mux_v
    port map (
            O => \N__35432\,
            I => \N__35418\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__35429\,
            I => \N__35418\
        );

    \I__7577\ : Odrv4
    port map (
            O => \N__35426\,
            I => rand_data_15
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__35423\,
            I => rand_data_15
        );

    \I__7575\ : Odrv4
    port map (
            O => \N__35418\,
            I => rand_data_15
        );

    \I__7574\ : InMux
    port map (
            O => \N__35411\,
            I => n16426
        );

    \I__7573\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35403\
        );

    \I__7572\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35400\
        );

    \I__7571\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35397\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__35403\,
            I => \N__35393\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__35400\,
            I => \N__35390\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35387\
        );

    \I__7567\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35383\
        );

    \I__7566\ : Span4Mux_h
    port map (
            O => \N__35393\,
            I => \N__35380\
        );

    \I__7565\ : Span4Mux_h
    port map (
            O => \N__35390\,
            I => \N__35375\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__35387\,
            I => \N__35375\
        );

    \I__7563\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35372\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35369\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__35380\,
            I => rand_data_16
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__35375\,
            I => rand_data_16
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__35372\,
            I => rand_data_16
        );

    \I__7558\ : Odrv12
    port map (
            O => \N__35369\,
            I => rand_data_16
        );

    \I__7557\ : InMux
    port map (
            O => \N__35360\,
            I => \bfn_9_31_0_\
        );

    \I__7556\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35352\
        );

    \I__7555\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35349\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35355\,
            I => \N__35346\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__35352\,
            I => \N__35342\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__35349\,
            I => \N__35339\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__35346\,
            I => \N__35336\
        );

    \I__7550\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35332\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__35342\,
            I => \N__35329\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__35339\,
            I => \N__35324\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__35336\,
            I => \N__35324\
        );

    \I__7546\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35321\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35318\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__35329\,
            I => rand_data_17
        );

    \I__7543\ : Odrv4
    port map (
            O => \N__35324\,
            I => rand_data_17
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__35321\,
            I => rand_data_17
        );

    \I__7541\ : Odrv12
    port map (
            O => \N__35318\,
            I => rand_data_17
        );

    \I__7540\ : InMux
    port map (
            O => \N__35309\,
            I => n16428
        );

    \I__7539\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35302\
        );

    \I__7538\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35299\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__35302\,
            I => \N__35293\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__35299\,
            I => \N__35293\
        );

    \I__7535\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35290\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__35293\,
            I => \N__35284\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__35290\,
            I => \N__35284\
        );

    \I__7532\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35280\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__35284\,
            I => \N__35277\
        );

    \I__7530\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35274\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35271\
        );

    \I__7528\ : Odrv4
    port map (
            O => \N__35277\,
            I => rand_data_18
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__35274\,
            I => rand_data_18
        );

    \I__7526\ : Odrv12
    port map (
            O => \N__35271\,
            I => rand_data_18
        );

    \I__7525\ : InMux
    port map (
            O => \N__35264\,
            I => n16429
        );

    \I__7524\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35257\
        );

    \I__7523\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35254\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35251\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35246\
        );

    \I__7520\ : Span4Mux_v
    port map (
            O => \N__35251\,
            I => \N__35243\
        );

    \I__7519\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35240\
        );

    \I__7518\ : InMux
    port map (
            O => \N__35249\,
            I => \N__35236\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__35246\,
            I => \N__35233\
        );

    \I__7516\ : Sp12to4
    port map (
            O => \N__35243\,
            I => \N__35228\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35228\
        );

    \I__7514\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35225\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35222\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__35233\,
            I => rand_data_19
        );

    \I__7511\ : Odrv12
    port map (
            O => \N__35228\,
            I => rand_data_19
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__35225\,
            I => rand_data_19
        );

    \I__7509\ : Odrv12
    port map (
            O => \N__35222\,
            I => rand_data_19
        );

    \I__7508\ : InMux
    port map (
            O => \N__35213\,
            I => n16430
        );

    \I__7507\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35206\
        );

    \I__7506\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35201\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__35206\,
            I => \N__35198\
        );

    \I__7504\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35195\
        );

    \I__7503\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35191\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35187\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__35198\,
            I => \N__35184\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__35195\,
            I => \N__35181\
        );

    \I__7499\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35178\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__35191\,
            I => \N__35175\
        );

    \I__7497\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35172\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__35187\,
            I => \N__35165\
        );

    \I__7495\ : Span4Mux_s3_h
    port map (
            O => \N__35184\,
            I => \N__35165\
        );

    \I__7494\ : Span4Mux_h
    port map (
            O => \N__35181\,
            I => \N__35165\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__35178\,
            I => rand_data_3
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__35175\,
            I => rand_data_3
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__35172\,
            I => rand_data_3
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__35165\,
            I => rand_data_3
        );

    \I__7489\ : InMux
    port map (
            O => \N__35156\,
            I => n16414
        );

    \I__7488\ : InMux
    port map (
            O => \N__35153\,
            I => \N__35150\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__35150\,
            I => \N__35146\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__35149\,
            I => \N__35143\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__35146\,
            I => \N__35140\
        );

    \I__7484\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35134\
        );

    \I__7483\ : Span4Mux_h
    port map (
            O => \N__35140\,
            I => \N__35130\
        );

    \I__7482\ : InMux
    port map (
            O => \N__35139\,
            I => \N__35127\
        );

    \I__7481\ : InMux
    port map (
            O => \N__35138\,
            I => \N__35122\
        );

    \I__7480\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35122\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35119\
        );

    \I__7478\ : InMux
    port map (
            O => \N__35133\,
            I => \N__35116\
        );

    \I__7477\ : Sp12to4
    port map (
            O => \N__35130\,
            I => \N__35111\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__35127\,
            I => \N__35111\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__35122\,
            I => rand_data_4
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__35119\,
            I => rand_data_4
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__35116\,
            I => rand_data_4
        );

    \I__7472\ : Odrv12
    port map (
            O => \N__35111\,
            I => rand_data_4
        );

    \I__7471\ : InMux
    port map (
            O => \N__35102\,
            I => n16415
        );

    \I__7470\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35094\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35088\
        );

    \I__7468\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35088\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__35094\,
            I => \N__35084\
        );

    \I__7466\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35081\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__35088\,
            I => \N__35078\
        );

    \I__7464\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35075\
        );

    \I__7463\ : Span4Mux_v
    port map (
            O => \N__35084\,
            I => \N__35072\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__35081\,
            I => \N__35066\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__35078\,
            I => \N__35066\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__35075\,
            I => \N__35063\
        );

    \I__7459\ : Span4Mux_h
    port map (
            O => \N__35072\,
            I => \N__35060\
        );

    \I__7458\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35057\
        );

    \I__7457\ : Span4Mux_h
    port map (
            O => \N__35066\,
            I => \N__35052\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__35063\,
            I => \N__35052\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__35060\,
            I => rand_data_5
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__35057\,
            I => rand_data_5
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__35052\,
            I => rand_data_5
        );

    \I__7452\ : InMux
    port map (
            O => \N__35045\,
            I => n16416
        );

    \I__7451\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35036\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35033\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35030\
        );

    \I__7448\ : CascadeMux
    port map (
            O => \N__35039\,
            I => \N__35026\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35036\,
            I => \N__35023\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__35033\,
            I => \N__35020\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__35030\,
            I => \N__35017\
        );

    \I__7444\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35014\
        );

    \I__7443\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35010\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__35023\,
            I => \N__35007\
        );

    \I__7441\ : Span4Mux_v
    port map (
            O => \N__35020\,
            I => \N__35002\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__35017\,
            I => \N__35002\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34999\
        );

    \I__7438\ : InMux
    port map (
            O => \N__35013\,
            I => \N__34996\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__35010\,
            I => \N__34993\
        );

    \I__7436\ : Odrv4
    port map (
            O => \N__35007\,
            I => rand_data_6
        );

    \I__7435\ : Odrv4
    port map (
            O => \N__35002\,
            I => rand_data_6
        );

    \I__7434\ : Odrv12
    port map (
            O => \N__34999\,
            I => rand_data_6
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__34996\,
            I => rand_data_6
        );

    \I__7432\ : Odrv12
    port map (
            O => \N__34993\,
            I => rand_data_6
        );

    \I__7431\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__34979\,
            I => \N__34975\
        );

    \I__7429\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34972\
        );

    \I__7428\ : Odrv12
    port map (
            O => \N__34975\,
            I => rand_setpoint_6
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__34972\,
            I => rand_setpoint_6
        );

    \I__7426\ : InMux
    port map (
            O => \N__34967\,
            I => n16417
        );

    \I__7425\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34960\
        );

    \I__7424\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34957\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34952\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__34957\,
            I => \N__34948\
        );

    \I__7421\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34945\
        );

    \I__7420\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34942\
        );

    \I__7419\ : Span4Mux_h
    port map (
            O => \N__34952\,
            I => \N__34939\
        );

    \I__7418\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34935\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__34948\,
            I => \N__34932\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__34945\,
            I => \N__34927\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__34942\,
            I => \N__34927\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__34939\,
            I => \N__34924\
        );

    \I__7413\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34921\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__34935\,
            I => \N__34918\
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__34932\,
            I => rand_data_7
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__34927\,
            I => rand_data_7
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__34924\,
            I => rand_data_7
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__34921\,
            I => rand_data_7
        );

    \I__7407\ : Odrv12
    port map (
            O => \N__34918\,
            I => rand_data_7
        );

    \I__7406\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34903\
        );

    \I__7405\ : CascadeMux
    port map (
            O => \N__34906\,
            I => \N__34900\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__34903\,
            I => \N__34897\
        );

    \I__7403\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34894\
        );

    \I__7402\ : Odrv4
    port map (
            O => \N__34897\,
            I => rand_setpoint_7
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__34894\,
            I => rand_setpoint_7
        );

    \I__7400\ : InMux
    port map (
            O => \N__34889\,
            I => n16418
        );

    \I__7399\ : InMux
    port map (
            O => \N__34886\,
            I => \N__34881\
        );

    \I__7398\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34877\
        );

    \I__7397\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34874\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__34881\,
            I => \N__34871\
        );

    \I__7395\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34868\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__34877\,
            I => \N__34862\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__34874\,
            I => \N__34862\
        );

    \I__7392\ : Span4Mux_v
    port map (
            O => \N__34871\,
            I => \N__34857\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__34868\,
            I => \N__34857\
        );

    \I__7390\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34853\
        );

    \I__7389\ : Span4Mux_h
    port map (
            O => \N__34862\,
            I => \N__34850\
        );

    \I__7388\ : Span4Mux_h
    port map (
            O => \N__34857\,
            I => \N__34847\
        );

    \I__7387\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34844\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34841\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__34850\,
            I => rand_data_8
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__34847\,
            I => rand_data_8
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__34844\,
            I => rand_data_8
        );

    \I__7382\ : Odrv12
    port map (
            O => \N__34841\,
            I => rand_data_8
        );

    \I__7381\ : InMux
    port map (
            O => \N__34832\,
            I => \bfn_9_30_0_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34826\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34821\
        );

    \I__7378\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34818\
        );

    \I__7377\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34814\
        );

    \I__7376\ : Span4Mux_v
    port map (
            O => \N__34821\,
            I => \N__34808\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__34818\,
            I => \N__34808\
        );

    \I__7374\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34805\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__34814\,
            I => \N__34802\
        );

    \I__7372\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34798\
        );

    \I__7371\ : Span4Mux_h
    port map (
            O => \N__34808\,
            I => \N__34795\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__34805\,
            I => \N__34792\
        );

    \I__7369\ : Span4Mux_h
    port map (
            O => \N__34802\,
            I => \N__34789\
        );

    \I__7368\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34786\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__34798\,
            I => \N__34783\
        );

    \I__7366\ : Odrv4
    port map (
            O => \N__34795\,
            I => rand_data_9
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__34792\,
            I => rand_data_9
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__34789\,
            I => rand_data_9
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__34786\,
            I => rand_data_9
        );

    \I__7362\ : Odrv12
    port map (
            O => \N__34783\,
            I => rand_data_9
        );

    \I__7361\ : InMux
    port map (
            O => \N__34772\,
            I => n16420
        );

    \I__7360\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34761\
        );

    \I__7358\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34758\
        );

    \I__7357\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34754\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__34761\,
            I => \N__34749\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__34758\,
            I => \N__34749\
        );

    \I__7354\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34746\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34742\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__34749\,
            I => \N__34737\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__34746\,
            I => \N__34737\
        );

    \I__7350\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34733\
        );

    \I__7349\ : Span4Mux_h
    port map (
            O => \N__34742\,
            I => \N__34730\
        );

    \I__7348\ : Span4Mux_h
    port map (
            O => \N__34737\,
            I => \N__34727\
        );

    \I__7347\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34724\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34721\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__34730\,
            I => rand_data_10
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__34727\,
            I => rand_data_10
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__34724\,
            I => rand_data_10
        );

    \I__7342\ : Odrv12
    port map (
            O => \N__34721\,
            I => rand_data_10
        );

    \I__7341\ : InMux
    port map (
            O => \N__34712\,
            I => n16421
        );

    \I__7340\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34706\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__34706\,
            I => \N__34702\
        );

    \I__7338\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34699\
        );

    \I__7337\ : Odrv12
    port map (
            O => \N__34702\,
            I => data_in_13_2
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__34699\,
            I => data_in_13_2
        );

    \I__7335\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34688\
        );

    \I__7334\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34688\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__34688\,
            I => data_in_12_2
        );

    \I__7332\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34680\
        );

    \I__7331\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34676\
        );

    \I__7330\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34669\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34666\
        );

    \I__7328\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34663\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__34676\,
            I => \N__34656\
        );

    \I__7326\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34653\
        );

    \I__7325\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34648\
        );

    \I__7324\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34648\
        );

    \I__7323\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34645\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34637\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__34666\,
            I => \N__34632\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__34663\,
            I => \N__34632\
        );

    \I__7319\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34629\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__34661\,
            I => \N__34623\
        );

    \I__7317\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34619\
        );

    \I__7316\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34616\
        );

    \I__7315\ : Span4Mux_s2_h
    port map (
            O => \N__34656\,
            I => \N__34607\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__34653\,
            I => \N__34607\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__34648\,
            I => \N__34607\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__34645\,
            I => \N__34607\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__34644\,
            I => \N__34602\
        );

    \I__7310\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34598\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__34642\,
            I => \N__34595\
        );

    \I__7308\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34589\
        );

    \I__7307\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34589\
        );

    \I__7306\ : Span4Mux_v
    port map (
            O => \N__34637\,
            I => \N__34582\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__34632\,
            I => \N__34582\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__34629\,
            I => \N__34582\
        );

    \I__7303\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34577\
        );

    \I__7302\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34577\
        );

    \I__7301\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34562\
        );

    \I__7300\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34562\
        );

    \I__7299\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34562\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__34619\,
            I => \N__34555\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__34616\,
            I => \N__34555\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__34607\,
            I => \N__34555\
        );

    \I__7295\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34545\
        );

    \I__7294\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34542\
        );

    \I__7293\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34537\
        );

    \I__7292\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34537\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__34598\,
            I => \N__34534\
        );

    \I__7290\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34529\
        );

    \I__7289\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34529\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34522\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__34582\,
            I => \N__34522\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__34577\,
            I => \N__34522\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34515\
        );

    \I__7284\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34515\
        );

    \I__7283\ : InMux
    port map (
            O => \N__34574\,
            I => \N__34515\
        );

    \I__7282\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34510\
        );

    \I__7281\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34510\
        );

    \I__7280\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34503\
        );

    \I__7279\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34503\
        );

    \I__7278\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34503\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34498\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__34555\,
            I => \N__34498\
        );

    \I__7275\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34491\
        );

    \I__7274\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34491\
        );

    \I__7273\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34491\
        );

    \I__7272\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34482\
        );

    \I__7271\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34482\
        );

    \I__7270\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34482\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34482\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__34545\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__34542\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__34537\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__34534\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__34529\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__34522\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__34515\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__34510\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__34503\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__34498\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__34491\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__34482\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1\
        );

    \I__7256\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34449\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34437\
        );

    \I__7254\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34437\
        );

    \I__7253\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34437\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34430\
        );

    \I__7251\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34427\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__34449\,
            I => \N__34423\
        );

    \I__7249\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34420\
        );

    \I__7248\ : InMux
    port map (
            O => \N__34447\,
            I => \N__34417\
        );

    \I__7247\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34414\
        );

    \I__7246\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34409\
        );

    \I__7245\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34409\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__34437\,
            I => \N__34405\
        );

    \I__7243\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34400\
        );

    \I__7242\ : InMux
    port map (
            O => \N__34435\,
            I => \N__34400\
        );

    \I__7241\ : InMux
    port map (
            O => \N__34434\,
            I => \N__34395\
        );

    \I__7240\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34395\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34390\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__34427\,
            I => \N__34387\
        );

    \I__7237\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34384\
        );

    \I__7236\ : Span4Mux_v
    port map (
            O => \N__34423\,
            I => \N__34379\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34379\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__34417\,
            I => \N__34376\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__34414\,
            I => \N__34371\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34371\
        );

    \I__7231\ : CascadeMux
    port map (
            O => \N__34408\,
            I => \N__34368\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__34405\,
            I => \N__34362\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34362\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__34395\,
            I => \N__34359\
        );

    \I__7227\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34354\
        );

    \I__7226\ : InMux
    port map (
            O => \N__34393\,
            I => \N__34354\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__34390\,
            I => \N__34341\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__34387\,
            I => \N__34341\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__34384\,
            I => \N__34341\
        );

    \I__7222\ : Span4Mux_v
    port map (
            O => \N__34379\,
            I => \N__34341\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__34376\,
            I => \N__34341\
        );

    \I__7220\ : Span4Mux_v
    port map (
            O => \N__34371\,
            I => \N__34341\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34336\
        );

    \I__7218\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34336\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__34362\,
            I => n63_adj_2642
        );

    \I__7216\ : Odrv12
    port map (
            O => \N__34359\,
            I => n63_adj_2642
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__34354\,
            I => n63_adj_2642
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__34341\,
            I => n63_adj_2642
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__34336\,
            I => n63_adj_2642
        );

    \I__7212\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34322\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34319\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__34319\,
            I => \N__34315\
        );

    \I__7209\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34312\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__34315\,
            I => \N__34309\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__34312\,
            I => \N__34304\
        );

    \I__7206\ : Span4Mux_h
    port map (
            O => \N__34309\,
            I => \N__34301\
        );

    \I__7205\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34296\
        );

    \I__7204\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34296\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__34304\,
            I => n63
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__34301\,
            I => n63
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__34296\,
            I => n63
        );

    \I__7200\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34285\
        );

    \I__7199\ : CascadeMux
    port map (
            O => \N__34288\,
            I => \N__34282\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__34285\,
            I => \N__34279\
        );

    \I__7197\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34276\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__34279\,
            I => \N__34273\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__34276\,
            I => \FRAME_MATCHER_next_state_0\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__34273\,
            I => \FRAME_MATCHER_next_state_0\
        );

    \I__7193\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34265\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__34265\,
            I => \N__34261\
        );

    \I__7191\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34258\
        );

    \I__7190\ : Odrv4
    port map (
            O => \N__34261\,
            I => data_in_17_5
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34258\,
            I => data_in_17_5
        );

    \I__7188\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34247\
        );

    \I__7186\ : Span4Mux_h
    port map (
            O => \N__34247\,
            I => \N__34242\
        );

    \I__7185\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34237\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__34242\,
            I => \c0.rx.r_SM_Main_2_N_2386_0\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__34237\,
            I => \c0.rx.r_SM_Main_2_N_2386_0\
        );

    \I__7181\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__34229\,
            I => \N__34226\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__34226\,
            I => \N__34223\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__34223\,
            I => \c0.rx.n18066\
        );

    \I__7177\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34214\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34214\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__34214\,
            I => \N__34208\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34205\
        );

    \I__7173\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34202\
        );

    \I__7172\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34198\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__34208\,
            I => \N__34195\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34192\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34189\
        );

    \I__7168\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34186\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34183\
        );

    \I__7166\ : Span4Mux_h
    port map (
            O => \N__34195\,
            I => \N__34180\
        );

    \I__7165\ : Span4Mux_s3_h
    port map (
            O => \N__34192\,
            I => \N__34171\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__34189\,
            I => \N__34171\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__34186\,
            I => \N__34171\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__34183\,
            I => \N__34171\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__34180\,
            I => rand_data_0
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__34171\,
            I => rand_data_0
        );

    \I__7159\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34161\
        );

    \I__7158\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34155\
        );

    \I__7157\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34155\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__34161\,
            I => \N__34152\
        );

    \I__7155\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34149\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__34155\,
            I => \N__34145\
        );

    \I__7153\ : Span4Mux_s3_h
    port map (
            O => \N__34152\,
            I => \N__34140\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34140\
        );

    \I__7151\ : InMux
    port map (
            O => \N__34148\,
            I => \N__34136\
        );

    \I__7150\ : Span4Mux_h
    port map (
            O => \N__34145\,
            I => \N__34133\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__34140\,
            I => \N__34130\
        );

    \I__7148\ : InMux
    port map (
            O => \N__34139\,
            I => \N__34127\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__34136\,
            I => \N__34124\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__34133\,
            I => rand_data_1
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__34130\,
            I => rand_data_1
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__34127\,
            I => rand_data_1
        );

    \I__7143\ : Odrv12
    port map (
            O => \N__34124\,
            I => rand_data_1
        );

    \I__7142\ : InMux
    port map (
            O => \N__34115\,
            I => n16412
        );

    \I__7141\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34109\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__34109\,
            I => \N__34105\
        );

    \I__7139\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34102\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__34105\,
            I => \N__34095\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34095\
        );

    \I__7136\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34092\
        );

    \I__7135\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34089\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__34095\,
            I => \N__34085\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34082\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__34089\,
            I => \N__34079\
        );

    \I__7131\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34075\
        );

    \I__7130\ : Sp12to4
    port map (
            O => \N__34085\,
            I => \N__34070\
        );

    \I__7129\ : Span12Mux_s4_h
    port map (
            O => \N__34082\,
            I => \N__34070\
        );

    \I__7128\ : Span4Mux_h
    port map (
            O => \N__34079\,
            I => \N__34067\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34064\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34075\,
            I => \N__34061\
        );

    \I__7125\ : Odrv12
    port map (
            O => \N__34070\,
            I => rand_data_2
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__34067\,
            I => rand_data_2
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34064\,
            I => rand_data_2
        );

    \I__7122\ : Odrv12
    port map (
            O => \N__34061\,
            I => rand_data_2
        );

    \I__7121\ : InMux
    port map (
            O => \N__34052\,
            I => n16413
        );

    \I__7120\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34046\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34042\
        );

    \I__7118\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34039\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__34042\,
            I => data_in_16_2
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__34039\,
            I => data_in_16_2
        );

    \I__7115\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34030\
        );

    \I__7114\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34027\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__34030\,
            I => \N__34024\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34021\
        );

    \I__7111\ : Span4Mux_h
    port map (
            O => \N__34024\,
            I => \N__34018\
        );

    \I__7110\ : Span4Mux_v
    port map (
            O => \N__34021\,
            I => \N__34015\
        );

    \I__7109\ : Sp12to4
    port map (
            O => \N__34018\,
            I => \N__34012\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__34015\,
            I => \N__34009\
        );

    \I__7107\ : Span12Mux_v
    port map (
            O => \N__34012\,
            I => \N__34006\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__34009\,
            I => \N__34003\
        );

    \I__7105\ : Odrv12
    port map (
            O => \N__34006\,
            I => n4
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__34003\,
            I => n4
        );

    \I__7103\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33994\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__33997\,
            I => \N__33991\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__33994\,
            I => \N__33988\
        );

    \I__7100\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33985\
        );

    \I__7099\ : Odrv12
    port map (
            O => \N__33988\,
            I => rx_data_3
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__33985\,
            I => rx_data_3
        );

    \I__7097\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33977\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__33977\,
            I => \N__33973\
        );

    \I__7095\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33970\
        );

    \I__7094\ : Span4Mux_h
    port map (
            O => \N__33973\,
            I => \N__33965\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__33970\,
            I => \N__33965\
        );

    \I__7092\ : Span4Mux_v
    port map (
            O => \N__33965\,
            I => \N__33962\
        );

    \I__7091\ : Span4Mux_v
    port map (
            O => \N__33962\,
            I => \N__33959\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__33956\,
            I => n4_adj_2582
        );

    \I__7088\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33949\
        );

    \I__7087\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33946\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__33949\,
            I => data_in_20_6
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__33946\,
            I => data_in_20_6
        );

    \I__7084\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__33938\,
            I => \N__33935\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__33935\,
            I => \N__33932\
        );

    \I__7081\ : Span4Mux_h
    port map (
            O => \N__33932\,
            I => \N__33928\
        );

    \I__7080\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33925\
        );

    \I__7079\ : Span4Mux_v
    port map (
            O => \N__33928\,
            I => \N__33919\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33919\
        );

    \I__7077\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33916\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__33919\,
            I => data_in_8_2
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__33916\,
            I => data_in_8_2
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__33911\,
            I => \N__33907\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__33910\,
            I => \N__33904\
        );

    \I__7072\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33895\
        );

    \I__7071\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33895\
        );

    \I__7070\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33895\
        );

    \I__7069\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33892\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33887\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33887\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__33887\,
            I => \N__33884\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__33884\,
            I => n8567
        );

    \I__7064\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33878\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__33878\,
            I => \N__33874\
        );

    \I__7062\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33871\
        );

    \I__7061\ : Odrv12
    port map (
            O => \N__33874\,
            I => data_in_11_2
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__33871\,
            I => data_in_11_2
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__33866\,
            I => \n9390_cascade_\
        );

    \I__7058\ : CascadeMux
    port map (
            O => \N__33863\,
            I => \n17681_cascade_\
        );

    \I__7057\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33856\
        );

    \I__7056\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33853\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__33856\,
            I => \N__33849\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__33853\,
            I => \N__33846\
        );

    \I__7053\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33843\
        );

    \I__7052\ : Span4Mux_h
    port map (
            O => \N__33849\,
            I => \N__33840\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__33846\,
            I => n16466
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__33843\,
            I => n16466
        );

    \I__7049\ : Odrv4
    port map (
            O => \N__33840\,
            I => n16466
        );

    \I__7048\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33828\
        );

    \I__7047\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33825\
        );

    \I__7046\ : InMux
    port map (
            O => \N__33831\,
            I => \N__33822\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__33828\,
            I => \N__33819\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33814\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__33822\,
            I => \N__33814\
        );

    \I__7042\ : Span4Mux_h
    port map (
            O => \N__33819\,
            I => \N__33811\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__33814\,
            I => \N__33808\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__33811\,
            I => n17356
        );

    \I__7039\ : Odrv4
    port map (
            O => \N__33808\,
            I => n17356
        );

    \I__7038\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__7036\ : Odrv12
    port map (
            O => \N__33797\,
            I => n18102
        );

    \I__7035\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33790\
        );

    \I__7034\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33786\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__33790\,
            I => \N__33783\
        );

    \I__7032\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33780\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33773\
        );

    \I__7030\ : Span4Mux_h
    port map (
            O => \N__33783\,
            I => \N__33773\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33773\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__33773\,
            I => \r_Clock_Count_2\
        );

    \I__7027\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33767\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__33767\,
            I => n13601
        );

    \I__7025\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33760\
        );

    \I__7024\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33757\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__33760\,
            I => \N__33754\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__33757\,
            I => \N__33751\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__33754\,
            I => \N__33747\
        );

    \I__7020\ : Span4Mux_h
    port map (
            O => \N__33751\,
            I => \N__33744\
        );

    \I__7019\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33741\
        );

    \I__7018\ : Span4Mux_h
    port map (
            O => \N__33747\,
            I => \N__33738\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__33744\,
            I => data_in_7_2
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__33741\,
            I => data_in_7_2
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__33738\,
            I => data_in_7_2
        );

    \I__7014\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33728\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__33725\,
            I => \N__33721\
        );

    \I__7011\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33718\
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__33721\,
            I => n13597
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__33718\,
            I => n13597
        );

    \I__7008\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33710\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__33710\,
            I => \N__33706\
        );

    \I__7006\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33703\
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__33706\,
            I => rx_data_6
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__33703\,
            I => rx_data_6
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__33698\,
            I => \N__33694\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__33697\,
            I => \N__33689\
        );

    \I__7001\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33686\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__33693\,
            I => \N__33683\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33679\
        );

    \I__6998\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33674\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__33686\,
            I => \N__33671\
        );

    \I__6996\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33668\
        );

    \I__6995\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33663\
        );

    \I__6994\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33660\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__33678\,
            I => \N__33657\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__33677\,
            I => \N__33654\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__33674\,
            I => \N__33651\
        );

    \I__6990\ : Span4Mux_h
    port map (
            O => \N__33671\,
            I => \N__33646\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33646\
        );

    \I__6988\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33640\
        );

    \I__6987\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33640\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__33663\,
            I => \N__33637\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__33660\,
            I => \N__33634\
        );

    \I__6984\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33630\
        );

    \I__6983\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33627\
        );

    \I__6982\ : Span4Mux_s2_h
    port map (
            O => \N__33651\,
            I => \N__33622\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__33646\,
            I => \N__33622\
        );

    \I__6980\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33619\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__33640\,
            I => \N__33614\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__33637\,
            I => \N__33614\
        );

    \I__6977\ : Span4Mux_s2_h
    port map (
            O => \N__33634\,
            I => \N__33611\
        );

    \I__6976\ : SRMux
    port map (
            O => \N__33633\,
            I => \N__33608\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33605\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33600\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__33622\,
            I => \N__33600\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__33619\,
            I => \N__33595\
        );

    \I__6971\ : Sp12to4
    port map (
            O => \N__33614\,
            I => \N__33595\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__33611\,
            I => \N__33592\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33589\
        );

    \I__6968\ : Span12Mux_s3_h
    port map (
            O => \N__33605\,
            I => \N__33586\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__33600\,
            I => \N__33583\
        );

    \I__6966\ : Span12Mux_h
    port map (
            O => \N__33595\,
            I => \N__33580\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__33592\,
            I => \N__33577\
        );

    \I__6964\ : Sp12to4
    port map (
            O => \N__33589\,
            I => \N__33572\
        );

    \I__6963\ : Span12Mux_v
    port map (
            O => \N__33586\,
            I => \N__33572\
        );

    \I__6962\ : Span4Mux_v
    port map (
            O => \N__33583\,
            I => \N__33569\
        );

    \I__6961\ : Odrv12
    port map (
            O => \N__33580\,
            I => \c0.n142\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__33577\,
            I => \c0.n142\
        );

    \I__6959\ : Odrv12
    port map (
            O => \N__33572\,
            I => \c0.n142\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__33569\,
            I => \c0.n142\
        );

    \I__6957\ : SRMux
    port map (
            O => \N__33560\,
            I => \N__33557\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__33554\,
            I => \N__33551\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__33551\,
            I => \c0.n1\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__33548\,
            I => \N__33544\
        );

    \I__6952\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33541\
        );

    \I__6951\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33538\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__33541\,
            I => \N__33535\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__33538\,
            I => \FRAME_MATCHER_next_state_1\
        );

    \I__6948\ : Odrv12
    port map (
            O => \N__33535\,
            I => \FRAME_MATCHER_next_state_1\
        );

    \I__6947\ : CascadeMux
    port map (
            O => \N__33530\,
            I => \N__33526\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__33529\,
            I => \N__33523\
        );

    \I__6945\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33519\
        );

    \I__6944\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33509\
        );

    \I__6943\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33509\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__33519\,
            I => \N__33505\
        );

    \I__6941\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33498\
        );

    \I__6940\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33498\
        );

    \I__6939\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33498\
        );

    \I__6938\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33495\
        );

    \I__6937\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33492\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__33509\,
            I => \N__33488\
        );

    \I__6935\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33485\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__33505\,
            I => \N__33480\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33480\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33477\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__33492\,
            I => \N__33474\
        );

    \I__6930\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33471\
        );

    \I__6929\ : Span4Mux_s3_h
    port map (
            O => \N__33488\,
            I => \N__33468\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33465\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__33480\,
            I => \N__33462\
        );

    \I__6926\ : Sp12to4
    port map (
            O => \N__33477\,
            I => \N__33456\
        );

    \I__6925\ : Span4Mux_v
    port map (
            O => \N__33474\,
            I => \N__33453\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__33471\,
            I => \N__33448\
        );

    \I__6923\ : Sp12to4
    port map (
            O => \N__33468\,
            I => \N__33448\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__33465\,
            I => \N__33445\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__33462\,
            I => \N__33442\
        );

    \I__6920\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33435\
        );

    \I__6919\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33435\
        );

    \I__6918\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33435\
        );

    \I__6917\ : Span12Mux_v
    port map (
            O => \N__33456\,
            I => \N__33428\
        );

    \I__6916\ : Sp12to4
    port map (
            O => \N__33453\,
            I => \N__33428\
        );

    \I__6915\ : Span12Mux_s8_v
    port map (
            O => \N__33448\,
            I => \N__33428\
        );

    \I__6914\ : Span4Mux_h
    port map (
            O => \N__33445\,
            I => \N__33425\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__33442\,
            I => \N__33422\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__33435\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__6911\ : Odrv12
    port map (
            O => \N__33428\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__33425\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__33422\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__6908\ : SRMux
    port map (
            O => \N__33413\,
            I => \N__33410\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__6906\ : Span4Mux_h
    port map (
            O => \N__33407\,
            I => \N__33404\
        );

    \I__6905\ : Span4Mux_h
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__6903\ : Odrv4
    port map (
            O => \N__33398\,
            I => \c0.n1_adj_2437\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__33395\,
            I => \r_SM_Main_2_N_2323_1_cascade_\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__33392\,
            I => \n17757_cascade_\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33384\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__33388\,
            I => \N__33381\
        );

    \I__6898\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33375\
        );

    \I__6897\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33368\
        );

    \I__6896\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33368\
        );

    \I__6895\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33368\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__33379\,
            I => \N__33364\
        );

    \I__6893\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33360\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__33375\,
            I => \N__33357\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33354\
        );

    \I__6890\ : CascadeMux
    port map (
            O => \N__33367\,
            I => \N__33351\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33346\
        );

    \I__6888\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33346\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__33360\,
            I => \N__33342\
        );

    \I__6886\ : Span4Mux_h
    port map (
            O => \N__33357\,
            I => \N__33339\
        );

    \I__6885\ : Span4Mux_v
    port map (
            O => \N__33354\,
            I => \N__33336\
        );

    \I__6884\ : InMux
    port map (
            O => \N__33351\,
            I => \N__33333\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33330\
        );

    \I__6882\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33327\
        );

    \I__6881\ : Sp12to4
    port map (
            O => \N__33342\,
            I => \N__33323\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__33339\,
            I => \N__33317\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__33336\,
            I => \N__33312\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33312\
        );

    \I__6877\ : Span4Mux_s3_h
    port map (
            O => \N__33330\,
            I => \N__33307\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__33327\,
            I => \N__33307\
        );

    \I__6875\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33304\
        );

    \I__6874\ : Span12Mux_v
    port map (
            O => \N__33323\,
            I => \N__33301\
        );

    \I__6873\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33296\
        );

    \I__6872\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33296\
        );

    \I__6871\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33293\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__33317\,
            I => \N__33288\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__33312\,
            I => \N__33288\
        );

    \I__6868\ : Span4Mux_v
    port map (
            O => \N__33307\,
            I => \N__33285\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__33304\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6866\ : Odrv12
    port map (
            O => \N__33301\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__33296\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__33293\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__33288\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6862\ : Odrv4
    port map (
            O => \N__33285\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6861\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__33269\,
            I => \N__33262\
        );

    \I__6859\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33255\
        );

    \I__6858\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33255\
        );

    \I__6857\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33255\
        );

    \I__6856\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33252\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__33262\,
            I => \N__33246\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33243\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33238\
        );

    \I__6852\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33231\
        );

    \I__6851\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33231\
        );

    \I__6850\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33231\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__33246\,
            I => \N__33226\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__33243\,
            I => \N__33223\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33218\
        );

    \I__6846\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33218\
        );

    \I__6845\ : Span4Mux_h
    port map (
            O => \N__33238\,
            I => \N__33214\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33211\
        );

    \I__6843\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33208\
        );

    \I__6842\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33205\
        );

    \I__6841\ : Span4Mux_v
    port map (
            O => \N__33226\,
            I => \N__33200\
        );

    \I__6840\ : Span4Mux_h
    port map (
            O => \N__33223\,
            I => \N__33200\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__33218\,
            I => \N__33197\
        );

    \I__6838\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33194\
        );

    \I__6837\ : Sp12to4
    port map (
            O => \N__33214\,
            I => \N__33187\
        );

    \I__6836\ : Sp12to4
    port map (
            O => \N__33211\,
            I => \N__33187\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__33208\,
            I => \N__33187\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__33205\,
            I => \N__33182\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__33200\,
            I => \N__33182\
        );

    \I__6832\ : Sp12to4
    port map (
            O => \N__33197\,
            I => \N__33175\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33175\
        );

    \I__6830\ : Span12Mux_s7_v
    port map (
            O => \N__33187\,
            I => \N__33175\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__33182\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6828\ : Odrv12
    port map (
            O => \N__33175\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__6827\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33163\
        );

    \I__6825\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33160\
        );

    \I__6824\ : Span4Mux_v
    port map (
            O => \N__33163\,
            I => \N__33153\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33153\
        );

    \I__6822\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33150\
        );

    \I__6821\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33145\
        );

    \I__6820\ : Span4Mux_h
    port map (
            O => \N__33153\,
            I => \N__33140\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__33150\,
            I => \N__33140\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33137\
        );

    \I__6817\ : CascadeMux
    port map (
            O => \N__33148\,
            I => \N__33134\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33131\
        );

    \I__6815\ : Span4Mux_v
    port map (
            O => \N__33140\,
            I => \N__33126\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__33137\,
            I => \N__33126\
        );

    \I__6813\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33123\
        );

    \I__6812\ : Span4Mux_h
    port map (
            O => \N__33131\,
            I => \N__33120\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__33126\,
            I => \N__33117\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__33123\,
            I => \N__33114\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__33120\,
            I => \N__33111\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__33117\,
            I => \N__33108\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__33114\,
            I => \N__33105\
        );

    \I__6806\ : Odrv4
    port map (
            O => \N__33111\,
            I => \c0.n157\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__33108\,
            I => \c0.n157\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__33105\,
            I => \c0.n157\
        );

    \I__6803\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33095\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__33089\,
            I => n18010
        );

    \I__6799\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33083\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__33080\,
            I => n9390
        );

    \I__6796\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__33074\,
            I => n7364
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__33071\,
            I => \N__33068\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__33062\,
            I => \N__33057\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33054\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33051\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__33057\,
            I => \N__33048\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33045\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__33051\,
            I => data_in_6_2
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__33048\,
            I => data_in_6_2
        );

    \I__6784\ : Odrv12
    port map (
            O => \N__33045\,
            I => data_in_6_2
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__33038\,
            I => \N__33034\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__33037\,
            I => \N__33031\
        );

    \I__6781\ : InMux
    port map (
            O => \N__33034\,
            I => \N__33028\
        );

    \I__6780\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33024\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33021\
        );

    \I__6778\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33018\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__33015\
        );

    \I__6776\ : Span4Mux_v
    port map (
            O => \N__33021\,
            I => \N__33011\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__33008\
        );

    \I__6774\ : Span4Mux_h
    port map (
            O => \N__33015\,
            I => \N__33005\
        );

    \I__6773\ : InMux
    port map (
            O => \N__33014\,
            I => \N__33002\
        );

    \I__6772\ : Sp12to4
    port map (
            O => \N__33011\,
            I => \N__32999\
        );

    \I__6771\ : Span4Mux_h
    port map (
            O => \N__33008\,
            I => \N__32994\
        );

    \I__6770\ : Span4Mux_h
    port map (
            O => \N__33005\,
            I => \N__32994\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33002\,
            I => data_in_5_2
        );

    \I__6768\ : Odrv12
    port map (
            O => \N__32999\,
            I => data_in_5_2
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__32994\,
            I => data_in_5_2
        );

    \I__6766\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32980\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__32986\,
            I => \N__32977\
        );

    \I__6764\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32974\
        );

    \I__6763\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32971\
        );

    \I__6762\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32968\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32965\
        );

    \I__6760\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32962\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32957\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__32971\,
            I => \N__32957\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32952\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__32965\,
            I => \N__32952\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32949\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__32957\,
            I => \N__32946\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__32952\,
            I => \N__32941\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__32949\,
            I => \N__32941\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__32946\,
            I => \c0.data_in_frame_10_5\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__32941\,
            I => \c0.data_in_frame_10_5\
        );

    \I__6749\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32932\
        );

    \I__6748\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32929\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32924\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32924\
        );

    \I__6745\ : Odrv12
    port map (
            O => \N__32924\,
            I => n2562
        );

    \I__6744\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32912\
        );

    \I__6743\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32912\
        );

    \I__6742\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32912\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__32912\,
            I => data_in_10_5
        );

    \I__6740\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32905\
        );

    \I__6739\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32902\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32899\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__32902\,
            I => \N__32896\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__32899\,
            I => \N__32893\
        );

    \I__6735\ : Span4Mux_v
    port map (
            O => \N__32896\,
            I => \N__32889\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__32893\,
            I => \N__32886\
        );

    \I__6733\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32883\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__32889\,
            I => \N__32880\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__32886\,
            I => data_in_9_5
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__32883\,
            I => data_in_9_5
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__32880\,
            I => data_in_9_5
        );

    \I__6728\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32870\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__32870\,
            I => \N__32866\
        );

    \I__6726\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32863\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__32866\,
            I => data_in_12_5
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__32863\,
            I => data_in_12_5
        );

    \I__6723\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32852\
        );

    \I__6722\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32852\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__32852\,
            I => data_in_11_5
        );

    \I__6720\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__32846\,
            I => n18098
        );

    \I__6718\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32838\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__32842\,
            I => \N__32835\
        );

    \I__6716\ : CEMux
    port map (
            O => \N__32841\,
            I => \N__32829\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__32838\,
            I => \N__32806\
        );

    \I__6714\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32801\
        );

    \I__6713\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32801\
        );

    \I__6712\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32793\
        );

    \I__6711\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32784\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32781\
        );

    \I__6709\ : CEMux
    port map (
            O => \N__32828\,
            I => \N__32778\
        );

    \I__6708\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32775\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__32826\,
            I => \N__32772\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__32825\,
            I => \N__32768\
        );

    \I__6705\ : CascadeMux
    port map (
            O => \N__32824\,
            I => \N__32765\
        );

    \I__6704\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32738\
        );

    \I__6703\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32738\
        );

    \I__6702\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32729\
        );

    \I__6701\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32729\
        );

    \I__6700\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32729\
        );

    \I__6699\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32729\
        );

    \I__6698\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32724\
        );

    \I__6697\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32724\
        );

    \I__6696\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32712\
        );

    \I__6695\ : CEMux
    port map (
            O => \N__32814\,
            I => \N__32709\
        );

    \I__6694\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32706\
        );

    \I__6693\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32699\
        );

    \I__6692\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32699\
        );

    \I__6691\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32699\
        );

    \I__6690\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32696\
        );

    \I__6689\ : Span4Mux_h
    port map (
            O => \N__32806\,
            I => \N__32691\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32691\
        );

    \I__6687\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32682\
        );

    \I__6686\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32682\
        );

    \I__6685\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32682\
        );

    \I__6684\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32682\
        );

    \I__6683\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32679\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__32793\,
            I => \N__32675\
        );

    \I__6681\ : CEMux
    port map (
            O => \N__32792\,
            I => \N__32672\
        );

    \I__6680\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32661\
        );

    \I__6679\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32661\
        );

    \I__6678\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32661\
        );

    \I__6677\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32661\
        );

    \I__6676\ : InMux
    port map (
            O => \N__32787\,
            I => \N__32661\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32656\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__32781\,
            I => \N__32656\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32653\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__32775\,
            I => \N__32644\
        );

    \I__6671\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32640\
        );

    \I__6670\ : CEMux
    port map (
            O => \N__32771\,
            I => \N__32595\
        );

    \I__6669\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32588\
        );

    \I__6668\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32588\
        );

    \I__6667\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32588\
        );

    \I__6666\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32581\
        );

    \I__6665\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32581\
        );

    \I__6664\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32581\
        );

    \I__6663\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32566\
        );

    \I__6662\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32566\
        );

    \I__6661\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32566\
        );

    \I__6660\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32566\
        );

    \I__6659\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32566\
        );

    \I__6658\ : InMux
    port map (
            O => \N__32755\,
            I => \N__32566\
        );

    \I__6657\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32566\
        );

    \I__6656\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32549\
        );

    \I__6655\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32549\
        );

    \I__6654\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32549\
        );

    \I__6653\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32549\
        );

    \I__6652\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32549\
        );

    \I__6651\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32549\
        );

    \I__6650\ : InMux
    port map (
            O => \N__32747\,
            I => \N__32549\
        );

    \I__6649\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32549\
        );

    \I__6648\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32542\
        );

    \I__6647\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32542\
        );

    \I__6646\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32542\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32539\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32536\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32533\
        );

    \I__6642\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32526\
        );

    \I__6641\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32526\
        );

    \I__6640\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32526\
        );

    \I__6639\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32513\
        );

    \I__6638\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32513\
        );

    \I__6637\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32513\
        );

    \I__6636\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32513\
        );

    \I__6635\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32513\
        );

    \I__6634\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32513\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32508\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__32709\,
            I => \N__32508\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__32706\,
            I => \N__32497\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32497\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__32696\,
            I => \N__32497\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__32691\,
            I => \N__32497\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__32682\,
            I => \N__32497\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__32679\,
            I => \N__32494\
        );

    \I__6625\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32491\
        );

    \I__6624\ : Span4Mux_h
    port map (
            O => \N__32675\,
            I => \N__32488\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32485\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32478\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__32656\,
            I => \N__32478\
        );

    \I__6620\ : Span4Mux_v
    port map (
            O => \N__32653\,
            I => \N__32478\
        );

    \I__6619\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32475\
        );

    \I__6618\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32464\
        );

    \I__6617\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32464\
        );

    \I__6616\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32464\
        );

    \I__6615\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32464\
        );

    \I__6614\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32464\
        );

    \I__6613\ : Sp12to4
    port map (
            O => \N__32644\,
            I => \N__32461\
        );

    \I__6612\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32458\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__32640\,
            I => \N__32455\
        );

    \I__6610\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32438\
        );

    \I__6609\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32438\
        );

    \I__6608\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32438\
        );

    \I__6607\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32438\
        );

    \I__6606\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32438\
        );

    \I__6605\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32438\
        );

    \I__6604\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32438\
        );

    \I__6603\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32438\
        );

    \I__6602\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32421\
        );

    \I__6601\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32421\
        );

    \I__6600\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32421\
        );

    \I__6599\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32421\
        );

    \I__6598\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32421\
        );

    \I__6597\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32421\
        );

    \I__6596\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32421\
        );

    \I__6595\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32421\
        );

    \I__6594\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32404\
        );

    \I__6593\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32404\
        );

    \I__6592\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32404\
        );

    \I__6591\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32404\
        );

    \I__6590\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32404\
        );

    \I__6589\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32404\
        );

    \I__6588\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32404\
        );

    \I__6587\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32404\
        );

    \I__6586\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32387\
        );

    \I__6585\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32387\
        );

    \I__6584\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32387\
        );

    \I__6583\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32387\
        );

    \I__6582\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32387\
        );

    \I__6581\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32387\
        );

    \I__6580\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32387\
        );

    \I__6579\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32387\
        );

    \I__6578\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32372\
        );

    \I__6577\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32372\
        );

    \I__6576\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32372\
        );

    \I__6575\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32372\
        );

    \I__6574\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32372\
        );

    \I__6573\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32372\
        );

    \I__6572\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32372\
        );

    \I__6571\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32365\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32365\
        );

    \I__6569\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32365\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__32595\,
            I => \N__32360\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32360\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__32581\,
            I => \N__32345\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32345\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32345\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32345\
        );

    \I__6562\ : Span4Mux_h
    port map (
            O => \N__32539\,
            I => \N__32345\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__32536\,
            I => \N__32345\
        );

    \I__6560\ : Span4Mux_v
    port map (
            O => \N__32533\,
            I => \N__32345\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__32526\,
            I => \N__32334\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__32513\,
            I => \N__32334\
        );

    \I__6557\ : Span4Mux_h
    port map (
            O => \N__32508\,
            I => \N__32334\
        );

    \I__6556\ : Span4Mux_v
    port map (
            O => \N__32497\,
            I => \N__32334\
        );

    \I__6555\ : Span4Mux_s2_h
    port map (
            O => \N__32494\,
            I => \N__32334\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32329\
        );

    \I__6553\ : Span4Mux_s3_h
    port map (
            O => \N__32488\,
            I => \N__32329\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__32485\,
            I => \N__32324\
        );

    \I__6551\ : Span4Mux_v
    port map (
            O => \N__32478\,
            I => \N__32324\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__32475\,
            I => \N__32317\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__32464\,
            I => \N__32317\
        );

    \I__6548\ : Span12Mux_v
    port map (
            O => \N__32461\,
            I => \N__32317\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__32458\,
            I => \N__32312\
        );

    \I__6546\ : Span12Mux_v
    port map (
            O => \N__32455\,
            I => \N__32312\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__32438\,
            I => n9606
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__32421\,
            I => n9606
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32404\,
            I => n9606
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__32387\,
            I => n9606
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__32372\,
            I => n9606
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__32365\,
            I => n9606
        );

    \I__6539\ : Odrv4
    port map (
            O => \N__32360\,
            I => n9606
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__32345\,
            I => n9606
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__32334\,
            I => n9606
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__32329\,
            I => n9606
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__32324\,
            I => n9606
        );

    \I__6534\ : Odrv12
    port map (
            O => \N__32317\,
            I => n9606
        );

    \I__6533\ : Odrv12
    port map (
            O => \N__32312\,
            I => n9606
        );

    \I__6532\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__32282\,
            I => \N__32279\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__32279\,
            I => \N__32275\
        );

    \I__6529\ : InMux
    port map (
            O => \N__32278\,
            I => \N__32272\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__32275\,
            I => \N__32269\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__32272\,
            I => data_out_frame2_7_7
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__32269\,
            I => data_out_frame2_7_7
        );

    \I__6525\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32260\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__32263\,
            I => \N__32257\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__32260\,
            I => \N__32253\
        );

    \I__6522\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32250\
        );

    \I__6521\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32247\
        );

    \I__6520\ : Span4Mux_v
    port map (
            O => \N__32253\,
            I => \N__32241\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32241\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__32247\,
            I => \N__32238\
        );

    \I__6517\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32235\
        );

    \I__6516\ : Sp12to4
    port map (
            O => \N__32241\,
            I => \N__32232\
        );

    \I__6515\ : Span4Mux_s3_h
    port map (
            O => \N__32238\,
            I => \N__32229\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__32235\,
            I => \N__32226\
        );

    \I__6513\ : Span12Mux_s11_v
    port map (
            O => \N__32232\,
            I => \N__32223\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__32229\,
            I => \c0.data_in_frame_9_7\
        );

    \I__6511\ : Odrv12
    port map (
            O => \N__32226\,
            I => \c0.data_in_frame_9_7\
        );

    \I__6510\ : Odrv12
    port map (
            O => \N__32223\,
            I => \c0.data_in_frame_9_7\
        );

    \I__6509\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32208\
        );

    \I__6508\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32208\
        );

    \I__6507\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32205\
        );

    \I__6506\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32202\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32199\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32196\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32193\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__32199\,
            I => \N__32190\
        );

    \I__6501\ : Span4Mux_v
    port map (
            O => \N__32196\,
            I => \N__32187\
        );

    \I__6500\ : Span4Mux_h
    port map (
            O => \N__32193\,
            I => \N__32184\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__32190\,
            I => \N__32181\
        );

    \I__6498\ : Span4Mux_h
    port map (
            O => \N__32187\,
            I => \N__32178\
        );

    \I__6497\ : Span4Mux_h
    port map (
            O => \N__32184\,
            I => \N__32175\
        );

    \I__6496\ : Sp12to4
    port map (
            O => \N__32181\,
            I => \N__32172\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__32178\,
            I => \c0.n17433\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__32175\,
            I => \c0.n17433\
        );

    \I__6493\ : Odrv12
    port map (
            O => \N__32172\,
            I => \c0.n17433\
        );

    \I__6492\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__32162\,
            I => \N__32158\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__32161\,
            I => \N__32155\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__32158\,
            I => \N__32152\
        );

    \I__6488\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32149\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__32152\,
            I => \N__32144\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__32149\,
            I => \N__32144\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__32144\,
            I => \N__32141\
        );

    \I__6484\ : Span4Mux_s1_h
    port map (
            O => \N__32141\,
            I => \N__32137\
        );

    \I__6483\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32134\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__32137\,
            I => \N__32131\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__32134\,
            I => data_in_7_7
        );

    \I__6480\ : Odrv4
    port map (
            O => \N__32131\,
            I => data_in_7_7
        );

    \I__6479\ : InMux
    port map (
            O => \N__32126\,
            I => \N__32123\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__6477\ : Span4Mux_v
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__32117\,
            I => n2573
        );

    \I__6475\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__32111\,
            I => \N__32107\
        );

    \I__6473\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32103\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__32107\,
            I => \N__32100\
        );

    \I__6471\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32097\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32094\
        );

    \I__6469\ : Span4Mux_v
    port map (
            O => \N__32100\,
            I => \N__32089\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32089\
        );

    \I__6467\ : Span4Mux_v
    port map (
            O => \N__32094\,
            I => \N__32084\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__32089\,
            I => \N__32084\
        );

    \I__6465\ : Sp12to4
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__6464\ : Odrv12
    port map (
            O => \N__32081\,
            I => \c0.data_in_frame_9_2\
        );

    \I__6463\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__32075\,
            I => \N__32072\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__32072\,
            I => \N__32069\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__32069\,
            I => n2565
        );

    \I__6459\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32061\
        );

    \I__6458\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32058\
        );

    \I__6457\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32054\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32049\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32058\,
            I => \N__32049\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__32057\,
            I => \N__32046\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__32042\
        );

    \I__6452\ : Span4Mux_h
    port map (
            O => \N__32049\,
            I => \N__32039\
        );

    \I__6451\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32036\
        );

    \I__6450\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32033\
        );

    \I__6449\ : Span4Mux_h
    port map (
            O => \N__32042\,
            I => \N__32026\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__32039\,
            I => \N__32026\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__32026\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__32033\,
            I => \N__32023\
        );

    \I__6445\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32020\
        );

    \I__6444\ : Span12Mux_s8_h
    port map (
            O => \N__32023\,
            I => \N__32017\
        );

    \I__6443\ : Sp12to4
    port map (
            O => \N__32020\,
            I => \N__32014\
        );

    \I__6442\ : Odrv12
    port map (
            O => \N__32017\,
            I => \c0.data_in_frame_10_2\
        );

    \I__6441\ : Odrv12
    port map (
            O => \N__32014\,
            I => \c0.data_in_frame_10_2\
        );

    \I__6440\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32006\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__32003\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__32003\,
            I => \N__32000\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__32000\,
            I => n2566
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__31997\,
            I => \N__31989\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__31996\,
            I => \N__31985\
        );

    \I__6434\ : CascadeMux
    port map (
            O => \N__31995\,
            I => \N__31982\
        );

    \I__6433\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31959\
        );

    \I__6432\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31959\
        );

    \I__6431\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31959\
        );

    \I__6430\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31959\
        );

    \I__6429\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31952\
        );

    \I__6428\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31952\
        );

    \I__6427\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31952\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__31981\,
            I => \N__31947\
        );

    \I__6425\ : CascadeMux
    port map (
            O => \N__31980\,
            I => \N__31944\
        );

    \I__6424\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31938\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__31978\,
            I => \N__31934\
        );

    \I__6422\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31929\
        );

    \I__6421\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31929\
        );

    \I__6420\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31914\
        );

    \I__6419\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31911\
        );

    \I__6418\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31908\
        );

    \I__6417\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31903\
        );

    \I__6416\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31894\
        );

    \I__6415\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31894\
        );

    \I__6414\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31894\
        );

    \I__6413\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31894\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__31959\,
            I => \N__31887\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31887\
        );

    \I__6410\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31878\
        );

    \I__6409\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31878\
        );

    \I__6408\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31878\
        );

    \I__6407\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31878\
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__31943\,
            I => \N__31872\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__31942\,
            I => \N__31867\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__31941\,
            I => \N__31864\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__31938\,
            I => \N__31861\
        );

    \I__6402\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31856\
        );

    \I__6401\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31856\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31853\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__31928\,
            I => \N__31844\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__31927\,
            I => \N__31841\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__31926\,
            I => \N__31835\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__31925\,
            I => \N__31832\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__31924\,
            I => \N__31825\
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__31923\,
            I => \N__31813\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__31922\,
            I => \N__31810\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__31921\,
            I => \N__31800\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__31920\,
            I => \N__31792\
        );

    \I__6390\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31786\
        );

    \I__6389\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31783\
        );

    \I__6388\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31780\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31777\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__31911\,
            I => \N__31774\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31771\
        );

    \I__6384\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31768\
        );

    \I__6383\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31765\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__31903\,
            I => \N__31760\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__31894\,
            I => \N__31760\
        );

    \I__6380\ : InMux
    port map (
            O => \N__31893\,
            I => \N__31755\
        );

    \I__6379\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31755\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__31887\,
            I => \N__31750\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__31878\,
            I => \N__31750\
        );

    \I__6376\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31747\
        );

    \I__6375\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31740\
        );

    \I__6374\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31740\
        );

    \I__6373\ : InMux
    port map (
            O => \N__31872\,
            I => \N__31740\
        );

    \I__6372\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31731\
        );

    \I__6371\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31731\
        );

    \I__6370\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31731\
        );

    \I__6369\ : InMux
    port map (
            O => \N__31864\,
            I => \N__31731\
        );

    \I__6368\ : Span4Mux_s3_h
    port map (
            O => \N__31861\,
            I => \N__31724\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31724\
        );

    \I__6366\ : Span4Mux_s3_h
    port map (
            O => \N__31853\,
            I => \N__31724\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__31852\,
            I => \N__31720\
        );

    \I__6364\ : CascadeMux
    port map (
            O => \N__31851\,
            I => \N__31717\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__31850\,
            I => \N__31714\
        );

    \I__6362\ : InMux
    port map (
            O => \N__31849\,
            I => \N__31701\
        );

    \I__6361\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31701\
        );

    \I__6360\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31701\
        );

    \I__6359\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31701\
        );

    \I__6358\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31701\
        );

    \I__6357\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31686\
        );

    \I__6356\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31686\
        );

    \I__6355\ : InMux
    port map (
            O => \N__31838\,
            I => \N__31686\
        );

    \I__6354\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31686\
        );

    \I__6353\ : InMux
    port map (
            O => \N__31832\,
            I => \N__31686\
        );

    \I__6352\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31686\
        );

    \I__6351\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31686\
        );

    \I__6350\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31675\
        );

    \I__6349\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31675\
        );

    \I__6348\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31675\
        );

    \I__6347\ : InMux
    port map (
            O => \N__31824\,
            I => \N__31675\
        );

    \I__6346\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31675\
        );

    \I__6345\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31664\
        );

    \I__6344\ : InMux
    port map (
            O => \N__31821\,
            I => \N__31664\
        );

    \I__6343\ : InMux
    port map (
            O => \N__31820\,
            I => \N__31664\
        );

    \I__6342\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31664\
        );

    \I__6341\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31664\
        );

    \I__6340\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31655\
        );

    \I__6339\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31655\
        );

    \I__6338\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31655\
        );

    \I__6337\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31655\
        );

    \I__6336\ : InMux
    port map (
            O => \N__31809\,
            I => \N__31642\
        );

    \I__6335\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31642\
        );

    \I__6334\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31642\
        );

    \I__6333\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31642\
        );

    \I__6332\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31642\
        );

    \I__6331\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31642\
        );

    \I__6330\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31631\
        );

    \I__6329\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31631\
        );

    \I__6328\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31631\
        );

    \I__6327\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31631\
        );

    \I__6326\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31631\
        );

    \I__6325\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31618\
        );

    \I__6324\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31618\
        );

    \I__6323\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31618\
        );

    \I__6322\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31618\
        );

    \I__6321\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31618\
        );

    \I__6320\ : InMux
    port map (
            O => \N__31789\,
            I => \N__31618\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31615\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__31783\,
            I => \N__31604\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31604\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__31777\,
            I => \N__31604\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__31774\,
            I => \N__31604\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__31771\,
            I => \N__31604\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31597\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__31765\,
            I => \N__31597\
        );

    \I__6311\ : Span4Mux_h
    port map (
            O => \N__31760\,
            I => \N__31597\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__31755\,
            I => \N__31592\
        );

    \I__6309\ : Span4Mux_s3_h
    port map (
            O => \N__31750\,
            I => \N__31592\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31583\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31583\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31583\
        );

    \I__6305\ : Span4Mux_h
    port map (
            O => \N__31724\,
            I => \N__31583\
        );

    \I__6304\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31570\
        );

    \I__6303\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31570\
        );

    \I__6302\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31570\
        );

    \I__6301\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31570\
        );

    \I__6300\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31570\
        );

    \I__6299\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31570\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__31701\,
            I => n1396
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__31686\,
            I => n1396
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__31675\,
            I => n1396
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__31664\,
            I => n1396
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__31655\,
            I => n1396
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__31642\,
            I => n1396
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__31631\,
            I => n1396
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__31618\,
            I => n1396
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__31615\,
            I => n1396
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__31604\,
            I => n1396
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__31597\,
            I => n1396
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__31592\,
            I => n1396
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__31583\,
            I => n1396
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__31570\,
            I => n1396
        );

    \I__6284\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31534\
        );

    \I__6282\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31531\
        );

    \I__6281\ : Span4Mux_h
    port map (
            O => \N__31534\,
            I => \N__31528\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__31531\,
            I => \N__31525\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__31528\,
            I => n2571
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__31525\,
            I => n2571
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__31520\,
            I => \N__31517\
        );

    \I__6276\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31513\
        );

    \I__6275\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31509\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31506\
        );

    \I__6273\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31502\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__31509\,
            I => \N__31499\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__31506\,
            I => \N__31496\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__31505\,
            I => \N__31493\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31486\
        );

    \I__6268\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31486\
        );

    \I__6267\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31486\
        );

    \I__6266\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31483\
        );

    \I__6265\ : Span4Mux_v
    port map (
            O => \N__31486\,
            I => \N__31478\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31478\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__31478\,
            I => \N__31475\
        );

    \I__6262\ : Odrv4
    port map (
            O => \N__31475\,
            I => \c0.data_in_frame_9_4\
        );

    \I__6261\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31466\
        );

    \I__6259\ : Span4Mux_v
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__31463\,
            I => \N__31459\
        );

    \I__6257\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31456\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__31459\,
            I => data_in_17_7
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__31456\,
            I => data_in_17_7
        );

    \I__6254\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31447\
        );

    \I__6253\ : InMux
    port map (
            O => \N__31450\,
            I => \N__31444\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__31447\,
            I => \N__31439\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__31444\,
            I => \N__31439\
        );

    \I__6250\ : Span4Mux_v
    port map (
            O => \N__31439\,
            I => \N__31436\
        );

    \I__6249\ : Odrv4
    port map (
            O => \N__31436\,
            I => n2564
        );

    \I__6248\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__31430\,
            I => \N__31426\
        );

    \I__6246\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31423\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__31426\,
            I => data_in_14_1
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__31423\,
            I => data_in_14_1
        );

    \I__6243\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31415\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__31415\,
            I => \N__31411\
        );

    \I__6241\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31406\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__31411\,
            I => \N__31403\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__31410\,
            I => \N__31400\
        );

    \I__6238\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31397\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__31406\,
            I => \N__31392\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__31403\,
            I => \N__31392\
        );

    \I__6235\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31389\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__31397\,
            I => data_in_2_1
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__31392\,
            I => data_in_2_1
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__31389\,
            I => data_in_2_1
        );

    \I__6231\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__31379\,
            I => \N__31373\
        );

    \I__6229\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31370\
        );

    \I__6228\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31367\
        );

    \I__6227\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31364\
        );

    \I__6226\ : Span4Mux_v
    port map (
            O => \N__31373\,
            I => \N__31358\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31358\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31355\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31352\
        );

    \I__6222\ : InMux
    port map (
            O => \N__31363\,
            I => \N__31349\
        );

    \I__6221\ : Span4Mux_h
    port map (
            O => \N__31358\,
            I => \N__31346\
        );

    \I__6220\ : Span4Mux_h
    port map (
            O => \N__31355\,
            I => \N__31341\
        );

    \I__6219\ : Span4Mux_h
    port map (
            O => \N__31352\,
            I => \N__31341\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__31349\,
            I => data_in_1_1
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__31346\,
            I => data_in_1_1
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__31341\,
            I => data_in_1_1
        );

    \I__6215\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31328\
        );

    \I__6214\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31328\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31328\,
            I => data_in_13_1
        );

    \I__6212\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31319\
        );

    \I__6211\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31319\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__31319\,
            I => data_in_12_1
        );

    \I__6209\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31313\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__31313\,
            I => \N__31310\
        );

    \I__6207\ : Span4Mux_h
    port map (
            O => \N__31310\,
            I => \N__31306\
        );

    \I__6206\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31303\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__31306\,
            I => data_in_11_1
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__31303\,
            I => data_in_11_1
        );

    \I__6203\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__31295\,
            I => \N__31292\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__31292\,
            I => \N__31288\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__31291\,
            I => \N__31284\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__31288\,
            I => \N__31281\
        );

    \I__6198\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31276\
        );

    \I__6197\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31276\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__31281\,
            I => data_in_6_6
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__31276\,
            I => data_in_6_6
        );

    \I__6194\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31267\
        );

    \I__6193\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31264\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__31267\,
            I => \N__31260\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31257\
        );

    \I__6190\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31254\
        );

    \I__6189\ : Span4Mux_v
    port map (
            O => \N__31260\,
            I => \N__31251\
        );

    \I__6188\ : Sp12to4
    port map (
            O => \N__31257\,
            I => \N__31248\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31244\
        );

    \I__6186\ : Sp12to4
    port map (
            O => \N__31251\,
            I => \N__31239\
        );

    \I__6185\ : Span12Mux_s11_v
    port map (
            O => \N__31248\,
            I => \N__31239\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31236\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__31244\,
            I => \N__31233\
        );

    \I__6182\ : Odrv12
    port map (
            O => \N__31239\,
            I => data_in_5_6
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__31236\,
            I => data_in_5_6
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__31233\,
            I => data_in_5_6
        );

    \I__6179\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31223\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__31220\,
            I => \N__31216\
        );

    \I__6176\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31213\
        );

    \I__6175\ : Sp12to4
    port map (
            O => \N__31216\,
            I => \N__31210\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__31213\,
            I => data_out_frame2_9_4
        );

    \I__6173\ : Odrv12
    port map (
            O => \N__31210\,
            I => data_out_frame2_9_4
        );

    \I__6172\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31201\
        );

    \I__6171\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31198\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__31201\,
            I => \N__31195\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__31198\,
            I => data_out_frame2_8_4
        );

    \I__6168\ : Odrv12
    port map (
            O => \N__31195\,
            I => data_out_frame2_8_4
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \N__31187\
        );

    \I__6166\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31184\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__31184\,
            I => \c0.n8\
        );

    \I__6164\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31178\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__31175\,
            I => \N__31172\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__31172\,
            I => \N__31168\
        );

    \I__6160\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31165\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__31168\,
            I => \N__31162\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__31165\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__31162\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__6156\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31147\
        );

    \I__6155\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31147\
        );

    \I__6154\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31147\
        );

    \I__6153\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31144\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__31147\,
            I => \N__31135\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__31144\,
            I => \N__31135\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__31143\,
            I => \N__31125\
        );

    \I__6149\ : CascadeMux
    port map (
            O => \N__31142\,
            I => \N__31119\
        );

    \I__6148\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31113\
        );

    \I__6147\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31113\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__31135\,
            I => \N__31110\
        );

    \I__6145\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31101\
        );

    \I__6144\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31101\
        );

    \I__6143\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31101\
        );

    \I__6142\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31101\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__31130\,
            I => \N__31097\
        );

    \I__6140\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31091\
        );

    \I__6139\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31088\
        );

    \I__6138\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31085\
        );

    \I__6137\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31081\
        );

    \I__6136\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31078\
        );

    \I__6135\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31066\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31066\
        );

    \I__6133\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31066\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__31059\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__31110\,
            I => \N__31059\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31059\
        );

    \I__6129\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31054\
        );

    \I__6128\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31054\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__31096\,
            I => \N__31049\
        );

    \I__6126\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31044\
        );

    \I__6125\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31044\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31036\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__31088\,
            I => \N__31036\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31036\
        );

    \I__6121\ : CascadeMux
    port map (
            O => \N__31084\,
            I => \N__31027\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__31081\,
            I => \N__31024\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31021\
        );

    \I__6118\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31016\
        );

    \I__6117\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31016\
        );

    \I__6116\ : InMux
    port map (
            O => \N__31075\,
            I => \N__31009\
        );

    \I__6115\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31009\
        );

    \I__6114\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31009\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__31066\,
            I => \N__31002\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__31059\,
            I => \N__31002\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31002\
        );

    \I__6110\ : InMux
    port map (
            O => \N__31053\,
            I => \N__30995\
        );

    \I__6109\ : InMux
    port map (
            O => \N__31052\,
            I => \N__30995\
        );

    \I__6108\ : InMux
    port map (
            O => \N__31049\,
            I => \N__30995\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__30992\
        );

    \I__6106\ : InMux
    port map (
            O => \N__31043\,
            I => \N__30975\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__31036\,
            I => \N__30972\
        );

    \I__6104\ : InMux
    port map (
            O => \N__31035\,
            I => \N__30969\
        );

    \I__6103\ : InMux
    port map (
            O => \N__31034\,
            I => \N__30957\
        );

    \I__6102\ : InMux
    port map (
            O => \N__31033\,
            I => \N__30957\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31032\,
            I => \N__30954\
        );

    \I__6100\ : InMux
    port map (
            O => \N__31031\,
            I => \N__30951\
        );

    \I__6099\ : InMux
    port map (
            O => \N__31030\,
            I => \N__30948\
        );

    \I__6098\ : InMux
    port map (
            O => \N__31027\,
            I => \N__30945\
        );

    \I__6097\ : Span4Mux_v
    port map (
            O => \N__31024\,
            I => \N__30942\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__31021\,
            I => \N__30931\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31016\,
            I => \N__30931\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__31009\,
            I => \N__30931\
        );

    \I__6093\ : Span4Mux_h
    port map (
            O => \N__31002\,
            I => \N__30931\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__30995\,
            I => \N__30931\
        );

    \I__6091\ : Span4Mux_v
    port map (
            O => \N__30992\,
            I => \N__30927\
        );

    \I__6090\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30924\
        );

    \I__6089\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30921\
        );

    \I__6088\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30916\
        );

    \I__6087\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30916\
        );

    \I__6086\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30911\
        );

    \I__6085\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30911\
        );

    \I__6084\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30908\
        );

    \I__6083\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30899\
        );

    \I__6082\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30899\
        );

    \I__6081\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30899\
        );

    \I__6080\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30899\
        );

    \I__6079\ : InMux
    port map (
            O => \N__30980\,
            I => \N__30892\
        );

    \I__6078\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30892\
        );

    \I__6077\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30892\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30885\
        );

    \I__6075\ : Sp12to4
    port map (
            O => \N__30972\,
            I => \N__30885\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30885\
        );

    \I__6073\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30876\
        );

    \I__6072\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30876\
        );

    \I__6071\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30876\
        );

    \I__6070\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30876\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__30964\,
            I => \N__30871\
        );

    \I__6068\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30866\
        );

    \I__6067\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30866\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__30957\,
            I => \N__30861\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30861\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30854\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__30948\,
            I => \N__30854\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30854\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__30942\,
            I => \N__30849\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__30931\,
            I => \N__30849\
        );

    \I__6059\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30846\
        );

    \I__6058\ : Span4Mux_v
    port map (
            O => \N__30927\,
            I => \N__30841\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__30924\,
            I => \N__30841\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30824\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30824\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__30911\,
            I => \N__30824\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__30908\,
            I => \N__30824\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30824\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30824\
        );

    \I__6050\ : Span12Mux_h
    port map (
            O => \N__30885\,
            I => \N__30824\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30824\
        );

    \I__6048\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30817\
        );

    \I__6047\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30817\
        );

    \I__6046\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30817\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30808\
        );

    \I__6044\ : Span4Mux_v
    port map (
            O => \N__30861\,
            I => \N__30808\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__30854\,
            I => \N__30808\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__30849\,
            I => \N__30808\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__30846\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__30841\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6039\ : Odrv12
    port map (
            O => \N__30824\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__30817\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__30808\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__6036\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30782\
        );

    \I__6035\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30782\
        );

    \I__6034\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30782\
        );

    \I__6033\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30777\
        );

    \I__6032\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30777\
        );

    \I__6031\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30774\
        );

    \I__6030\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30755\
        );

    \I__6029\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30750\
        );

    \I__6028\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30747\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30740\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__30777\,
            I => \N__30740\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__30774\,
            I => \N__30740\
        );

    \I__6024\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30726\
        );

    \I__6023\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30726\
        );

    \I__6022\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30726\
        );

    \I__6021\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30723\
        );

    \I__6020\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30719\
        );

    \I__6019\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30714\
        );

    \I__6018\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30714\
        );

    \I__6017\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30699\
        );

    \I__6016\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30699\
        );

    \I__6015\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30699\
        );

    \I__6014\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30699\
        );

    \I__6013\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30699\
        );

    \I__6012\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30699\
        );

    \I__6011\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30699\
        );

    \I__6010\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30696\
        );

    \I__6009\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30691\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30688\
        );

    \I__6007\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30685\
        );

    \I__6006\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30682\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__30750\,
            I => \N__30675\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__30747\,
            I => \N__30675\
        );

    \I__6003\ : Span4Mux_s2_v
    port map (
            O => \N__30740\,
            I => \N__30675\
        );

    \I__6002\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30664\
        );

    \I__6001\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30664\
        );

    \I__6000\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30655\
        );

    \I__5999\ : InMux
    port map (
            O => \N__30736\,
            I => \N__30655\
        );

    \I__5998\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30655\
        );

    \I__5997\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30655\
        );

    \I__5996\ : InMux
    port map (
            O => \N__30733\,
            I => \N__30652\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30649\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__30723\,
            I => \N__30646\
        );

    \I__5993\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30640\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30631\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__30714\,
            I => \N__30631\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__30699\,
            I => \N__30631\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__30696\,
            I => \N__30631\
        );

    \I__5988\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30626\
        );

    \I__5987\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30626\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__30691\,
            I => \N__30622\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30617\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30617\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__30682\,
            I => \N__30612\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__30675\,
            I => \N__30612\
        );

    \I__5981\ : InMux
    port map (
            O => \N__30674\,
            I => \N__30609\
        );

    \I__5980\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30604\
        );

    \I__5979\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30604\
        );

    \I__5978\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30601\
        );

    \I__5977\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30598\
        );

    \I__5976\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30595\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30590\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30590\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30585\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__30649\,
            I => \N__30585\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__30646\,
            I => \N__30582\
        );

    \I__5970\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30575\
        );

    \I__5969\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30575\
        );

    \I__5968\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30575\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__30640\,
            I => \N__30568\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__30631\,
            I => \N__30568\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__30626\,
            I => \N__30568\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__30625\,
            I => \N__30565\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__30622\,
            I => \N__30555\
        );

    \I__5962\ : Span4Mux_v
    port map (
            O => \N__30617\,
            I => \N__30555\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__30612\,
            I => \N__30550\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30550\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__30604\,
            I => \N__30537\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__30601\,
            I => \N__30537\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__30598\,
            I => \N__30537\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__30595\,
            I => \N__30537\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__30590\,
            I => \N__30537\
        );

    \I__5954\ : Span4Mux_v
    port map (
            O => \N__30585\,
            I => \N__30537\
        );

    \I__5953\ : Span4Mux_h
    port map (
            O => \N__30582\,
            I => \N__30532\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30532\
        );

    \I__5951\ : Span4Mux_v
    port map (
            O => \N__30568\,
            I => \N__30529\
        );

    \I__5950\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30526\
        );

    \I__5949\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30523\
        );

    \I__5948\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30514\
        );

    \I__5947\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30514\
        );

    \I__5946\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30514\
        );

    \I__5945\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30514\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__30555\,
            I => \N__30509\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__30550\,
            I => \N__30509\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__30537\,
            I => \N__30504\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__30532\,
            I => \N__30504\
        );

    \I__5940\ : Span4Mux_h
    port map (
            O => \N__30529\,
            I => \N__30501\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__30526\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__30523\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__30514\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__30509\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__30504\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__30501\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5933\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30485\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30482\
        );

    \I__5931\ : Span4Mux_s3_h
    port map (
            O => \N__30482\,
            I => \N__30479\
        );

    \I__5930\ : Span4Mux_h
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__30476\,
            I => \c0.n18086\
        );

    \I__5928\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30469\
        );

    \I__5927\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30466\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__30469\,
            I => \N__30463\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30457\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__30463\,
            I => \N__30457\
        );

    \I__5923\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30454\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__30457\,
            I => \N__30451\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__30454\,
            I => data_in_10_7
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__30451\,
            I => data_in_10_7
        );

    \I__5919\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30440\
        );

    \I__5918\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30440\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__30440\,
            I => data_in_11_7
        );

    \I__5916\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30431\
        );

    \I__5915\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30431\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__30431\,
            I => data_in_12_7
        );

    \I__5913\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30422\
        );

    \I__5912\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30422\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__30422\,
            I => data_in_13_7
        );

    \I__5910\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__5909\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30413\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__30413\,
            I => data_in_14_7
        );

    \I__5907\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30403\
        );

    \I__5905\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30400\
        );

    \I__5904\ : Odrv12
    port map (
            O => \N__30403\,
            I => data_in_16_7
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__30400\,
            I => data_in_16_7
        );

    \I__5902\ : InMux
    port map (
            O => \N__30395\,
            I => \N__30389\
        );

    \I__5901\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30389\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__30389\,
            I => data_in_15_7
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__30386\,
            I => \c0.rx.n97_cascade_\
        );

    \I__5898\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__30380\,
            I => \c0.rx.n17345\
        );

    \I__5896\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30367\
        );

    \I__5895\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30367\
        );

    \I__5894\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30364\
        );

    \I__5893\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30359\
        );

    \I__5892\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30359\
        );

    \I__5891\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30356\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__30367\,
            I => n13880
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__30364\,
            I => n13880
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__30359\,
            I => n13880
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__30356\,
            I => n13880
        );

    \I__5886\ : InMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30344\,
            I => n222
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__30341\,
            I => \N__30338\
        );

    \I__5883\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30335\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N__30330\
        );

    \I__5881\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30327\
        );

    \I__5880\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30324\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__30330\,
            I => \r_Clock_Count_4_adj_2620\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__30327\,
            I => \r_Clock_Count_4_adj_2620\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__30324\,
            I => \r_Clock_Count_4_adj_2620\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \N__30311\
        );

    \I__5875\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30306\
        );

    \I__5874\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30295\
        );

    \I__5873\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30295\
        );

    \I__5872\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30295\
        );

    \I__5871\ : InMux
    port map (
            O => \N__30310\,
            I => \N__30295\
        );

    \I__5870\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30295\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__30306\,
            I => \N__30288\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__30295\,
            I => \N__30288\
        );

    \I__5867\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30283\
        );

    \I__5866\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30283\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__30288\,
            I => n3
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__30283\,
            I => n3
        );

    \I__5863\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__30275\,
            I => \c0.rx.n18001\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__30272\,
            I => \n17856_cascade_\
        );

    \I__5860\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__30266\,
            I => n17855
        );

    \I__5858\ : IoInMux
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__5856\ : IoSpan4Mux
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__30254\,
            I => \LED_c\
        );

    \I__5854\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30247\
        );

    \I__5853\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30244\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__30247\,
            I => \c0.rx.n112\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__30244\,
            I => \c0.rx.n112\
        );

    \I__5850\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30236\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__30236\,
            I => \N__30232\
        );

    \I__5848\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30229\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__30232\,
            I => \N__30226\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__30229\,
            I => data_out_frame2_7_4
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__30226\,
            I => data_out_frame2_7_4
        );

    \I__5844\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30218\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__5842\ : Span4Mux_s2_v
    port map (
            O => \N__30215\,
            I => \N__30211\
        );

    \I__5841\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30208\
        );

    \I__5840\ : Span4Mux_h
    port map (
            O => \N__30211\,
            I => \N__30205\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__30208\,
            I => data_out_frame2_6_4
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__30205\,
            I => data_out_frame2_6_4
        );

    \I__5837\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30197\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__30197\,
            I => \c0.n5_adj_2425\
        );

    \I__5835\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30191\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__30188\,
            I => \N__30185\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__30185\,
            I => \c0.rx.n79\
        );

    \I__5831\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__5829\ : Odrv12
    port map (
            O => \N__30176\,
            I => \c0.rx.n18597\
        );

    \I__5828\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30170\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__30161\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__5823\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30152\
        );

    \I__5822\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30152\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__30152\,
            I => \c0.rx.n13537\
        );

    \I__5820\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30143\
        );

    \I__5819\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30143\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__30143\,
            I => \c0.rx.n4_adj_2424\
        );

    \I__5817\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30133\
        );

    \I__5816\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30133\
        );

    \I__5815\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30130\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__30133\,
            I => \c0.rx.n17381\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__30130\,
            I => \c0.rx.n17381\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__30125\,
            I => \c0.rx.n18003_cascade_\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__30122\,
            I => \n13880_cascade_\
        );

    \I__5810\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30113\
        );

    \I__5809\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30113\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__30113\,
            I => \c0.rx.n10193\
        );

    \I__5807\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30104\
        );

    \I__5806\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30101\
        );

    \I__5805\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30096\
        );

    \I__5804\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30096\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__30104\,
            I => \r_Clock_Count_2_adj_2622\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__30101\,
            I => \r_Clock_Count_2_adj_2622\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__30096\,
            I => \r_Clock_Count_2_adj_2622\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \N__30086\
        );

    \I__5799\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30077\
        );

    \I__5798\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30077\
        );

    \I__5797\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30077\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__30077\,
            I => \c0.rx.n124\
        );

    \I__5795\ : CascadeMux
    port map (
            O => \N__30074\,
            I => \N__30071\
        );

    \I__5794\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30065\
        );

    \I__5793\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30062\
        );

    \I__5792\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30059\
        );

    \I__5791\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30056\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30065\,
            I => \r_Clock_Count_3_adj_2621\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__30062\,
            I => \r_Clock_Count_3_adj_2621\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__30059\,
            I => \r_Clock_Count_3_adj_2621\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__30056\,
            I => \r_Clock_Count_3_adj_2621\
        );

    \I__5786\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__5784\ : Span4Mux_s2_h
    port map (
            O => \N__30041\,
            I => \N__30037\
        );

    \I__5783\ : InMux
    port map (
            O => \N__30040\,
            I => \N__30034\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__30037\,
            I => \N__30031\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__30034\,
            I => data_out_frame2_13_0
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__30031\,
            I => data_out_frame2_13_0
        );

    \I__5779\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30020\
        );

    \I__5778\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30020\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__30020\,
            I => data_in_18_5
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \n8562_cascade_\
        );

    \I__5775\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30010\
        );

    \I__5774\ : InMux
    port map (
            O => \N__30013\,
            I => \N__30007\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__30010\,
            I => rx_data_2
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__30007\,
            I => rx_data_2
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__30002\,
            I => \c0.rx.n2_cascade_\
        );

    \I__5770\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__29996\,
            I => \c0.rx.n2\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__29993\,
            I => \N__29989\
        );

    \I__5767\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29985\
        );

    \I__5766\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29982\
        );

    \I__5765\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29979\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29976\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__29982\,
            I => \r_Clock_Count_0_adj_2624\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__29979\,
            I => \r_Clock_Count_0_adj_2624\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__29976\,
            I => \r_Clock_Count_0_adj_2624\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29966\
        );

    \I__5759\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29962\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__29965\,
            I => \N__29959\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29955\
        );

    \I__5756\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29952\
        );

    \I__5755\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29949\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__29955\,
            I => \r_Clock_Count_1_adj_2623\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__29952\,
            I => \r_Clock_Count_1_adj_2623\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__29949\,
            I => \r_Clock_Count_1_adj_2623\
        );

    \I__5751\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__29939\,
            I => \N__29935\
        );

    \I__5749\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29932\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__29935\,
            I => data_in_19_0
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__29932\,
            I => data_in_19_0
        );

    \I__5746\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29923\
        );

    \I__5745\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29920\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29916\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__29920\,
            I => \N__29913\
        );

    \I__5742\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29910\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__29916\,
            I => \N__29907\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__29913\,
            I => \N__29904\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__29910\,
            I => data_in_10_0
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__29907\,
            I => data_in_10_0
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__29904\,
            I => data_in_10_0
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__29897\,
            I => \N__29893\
        );

    \I__5735\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29890\
        );

    \I__5734\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29887\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__29890\,
            I => rx_data_4
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__29887\,
            I => rx_data_4
        );

    \I__5731\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29878\
        );

    \I__5730\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29875\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__29878\,
            I => data_in_15_2
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__29875\,
            I => data_in_15_2
        );

    \I__5727\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29866\
        );

    \I__5726\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29863\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__29866\,
            I => data_in_14_2
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__29863\,
            I => data_in_14_2
        );

    \I__5723\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29855\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29852\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__29852\,
            I => \N__29848\
        );

    \I__5720\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29845\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__29848\,
            I => \N__29841\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__29845\,
            I => \N__29838\
        );

    \I__5717\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29835\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__29841\,
            I => data_in_4_2
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__29838\,
            I => data_in_4_2
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__29835\,
            I => data_in_4_2
        );

    \I__5713\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29823\
        );

    \I__5712\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29820\
        );

    \I__5711\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29817\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29814\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__29820\,
            I => data_in_9_7
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__29817\,
            I => data_in_9_7
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__29814\,
            I => data_in_9_7
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__5705\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__29801\,
            I => \N__29797\
        );

    \I__5703\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29794\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__29794\,
            I => \N__29788\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__29791\,
            I => \N__29785\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__29788\,
            I => \N__29781\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__29785\,
            I => \N__29778\
        );

    \I__5697\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29775\
        );

    \I__5696\ : Span4Mux_h
    port map (
            O => \N__29781\,
            I => \N__29772\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__29778\,
            I => \N__29769\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__29775\,
            I => data_in_8_7
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__29772\,
            I => data_in_8_7
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__29769\,
            I => data_in_8_7
        );

    \I__5691\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29759\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__29759\,
            I => \c0.n10_adj_2536\
        );

    \I__5689\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29753\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__29750\,
            I => n18101
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__5685\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__29735\,
            I => \N__29730\
        );

    \I__5681\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29727\
        );

    \I__5680\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29724\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__29730\,
            I => data_in_8_3
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__29727\,
            I => data_in_8_3
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__29724\,
            I => data_in_8_3
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__29717\,
            I => \n8517_cascade_\
        );

    \I__5675\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29705\
        );

    \I__5674\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29705\
        );

    \I__5673\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29705\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__29702\,
            I => \N__29696\
        );

    \I__5670\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29689\
        );

    \I__5669\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29689\
        );

    \I__5668\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29689\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__29696\,
            I => \N__29684\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__29689\,
            I => \N__29684\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__29684\,
            I => n17366
        );

    \I__5664\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29678\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__29678\,
            I => \N__29673\
        );

    \I__5662\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29668\
        );

    \I__5661\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29668\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__29673\,
            I => \N__29665\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__29668\,
            I => data_in_9_3
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__29665\,
            I => data_in_9_3
        );

    \I__5657\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29655\
        );

    \I__5656\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29652\
        );

    \I__5655\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29649\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__29655\,
            I => \r_Clock_Count_0\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__29652\,
            I => \r_Clock_Count_0\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__29649\,
            I => \r_Clock_Count_0\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__29642\,
            I => \N__29637\
        );

    \I__5650\ : InMux
    port map (
            O => \N__29641\,
            I => \N__29634\
        );

    \I__5649\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29631\
        );

    \I__5648\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29628\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__29634\,
            I => \r_Clock_Count_5\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__29631\,
            I => \r_Clock_Count_5\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__29628\,
            I => \r_Clock_Count_5\
        );

    \I__5644\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29616\
        );

    \I__5643\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29613\
        );

    \I__5642\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29610\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__29616\,
            I => \r_Clock_Count_3\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__29613\,
            I => \r_Clock_Count_3\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__29610\,
            I => \r_Clock_Count_3\
        );

    \I__5638\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29598\
        );

    \I__5637\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29595\
        );

    \I__5636\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29592\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__29598\,
            I => \r_Clock_Count_4\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__29595\,
            I => \r_Clock_Count_4\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__29592\,
            I => \r_Clock_Count_4\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__29585\,
            I => \c0.tx.n10_cascade_\
        );

    \I__5631\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29574\
        );

    \I__5629\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29569\
        );

    \I__5628\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29569\
        );

    \I__5627\ : Odrv12
    port map (
            O => \N__29574\,
            I => \r_Clock_Count_1\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__29569\,
            I => \r_Clock_Count_1\
        );

    \I__5625\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29558\
        );

    \I__5624\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29558\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29554\
        );

    \I__5622\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29550\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__29554\,
            I => \N__29547\
        );

    \I__5620\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29544\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__29550\,
            I => \N__29541\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__29547\,
            I => \N__29538\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__29544\,
            I => data_in_5_5
        );

    \I__5616\ : Odrv12
    port map (
            O => \N__29541\,
            I => data_in_5_5
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__29538\,
            I => data_in_5_5
        );

    \I__5614\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29527\
        );

    \I__5613\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29524\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__29527\,
            I => \N__29518\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29518\
        );

    \I__5610\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29515\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__29518\,
            I => \N__29512\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__29515\,
            I => data_in_10_1
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__29512\,
            I => data_in_10_1
        );

    \I__5606\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29503\
        );

    \I__5605\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29500\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29497\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29494\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__29497\,
            I => \N__29491\
        );

    \I__5601\ : Span12Mux_v
    port map (
            O => \N__29494\,
            I => \N__29488\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__5599\ : Odrv12
    port map (
            O => \N__29488\,
            I => \c0.n17544\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__29485\,
            I => \c0.n17544\
        );

    \I__5597\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29476\
        );

    \I__5596\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29473\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__29476\,
            I => \N__29470\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__29473\,
            I => \N__29467\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__29470\,
            I => \N__29464\
        );

    \I__5592\ : Span12Mux_h
    port map (
            O => \N__29467\,
            I => \N__29461\
        );

    \I__5591\ : Span4Mux_v
    port map (
            O => \N__29464\,
            I => \N__29458\
        );

    \I__5590\ : Odrv12
    port map (
            O => \N__29461\,
            I => \c0.n8056\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__29458\,
            I => \c0.n8056\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__29453\,
            I => \n2566_cascade_\
        );

    \I__5587\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29447\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29443\
        );

    \I__5585\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29440\
        );

    \I__5584\ : Span4Mux_h
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__29437\,
            I => n2561
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__29434\,
            I => n2561
        );

    \I__5580\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29426\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__29426\,
            I => \c0.n19\
        );

    \I__5578\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29420\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29416\
        );

    \I__5576\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29413\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__29416\,
            I => \N__29409\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29406\
        );

    \I__5573\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29403\
        );

    \I__5572\ : Span4Mux_h
    port map (
            O => \N__29409\,
            I => \N__29400\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__29406\,
            I => data_in_9_0
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__29403\,
            I => data_in_9_0
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__29400\,
            I => data_in_9_0
        );

    \I__5568\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29385\
        );

    \I__5567\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29382\
        );

    \I__5566\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29375\
        );

    \I__5565\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29375\
        );

    \I__5564\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29375\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__29388\,
            I => \N__29372\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29365\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__29382\,
            I => \N__29365\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29365\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29362\
        );

    \I__5558\ : Span12Mux_s9_v
    port map (
            O => \N__29365\,
            I => \N__29357\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29357\
        );

    \I__5556\ : Span12Mux_h
    port map (
            O => \N__29357\,
            I => \N__29354\
        );

    \I__5555\ : Odrv12
    port map (
            O => \N__29354\,
            I => \c0.data_in_frame_9_0\
        );

    \I__5554\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__29345\,
            I => \N__29341\
        );

    \I__5551\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29338\
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__29341\,
            I => n2575
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__29338\,
            I => n2575
        );

    \I__5548\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29327\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__29327\,
            I => \N__29324\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__29324\,
            I => \N__29320\
        );

    \I__5544\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29317\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__29320\,
            I => \c0.n17504\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__29317\,
            I => \c0.n17504\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__29312\,
            I => \c0.n6_adj_2541_cascade_\
        );

    \I__5540\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__5538\ : Span4Mux_v
    port map (
            O => \N__29303\,
            I => \N__29300\
        );

    \I__5537\ : Sp12to4
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__5536\ : Odrv12
    port map (
            O => \N__29297\,
            I => \c0.n17591\
        );

    \I__5535\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__5533\ : Span4Mux_s2_v
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__5532\ : Span4Mux_v
    port map (
            O => \N__29285\,
            I => \N__29282\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__29282\,
            I => \c0.data_out_frame2_20_4\
        );

    \I__5530\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29276\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__29276\,
            I => \N__29273\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__29273\,
            I => \N__29270\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__29270\,
            I => \N__29266\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29263\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__29266\,
            I => \c0.n17488\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__29263\,
            I => \c0.n17488\
        );

    \I__5523\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29254\
        );

    \I__5522\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29251\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29248\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29240\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__29248\,
            I => \N__29240\
        );

    \I__5518\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29235\
        );

    \I__5517\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29235\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__29245\,
            I => \N__29232\
        );

    \I__5515\ : Sp12to4
    port map (
            O => \N__29240\,
            I => \N__29229\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29226\
        );

    \I__5513\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29223\
        );

    \I__5512\ : Span12Mux_s11_v
    port map (
            O => \N__29229\,
            I => \N__29220\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__29226\,
            I => \N__29215\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__29223\,
            I => \N__29215\
        );

    \I__5509\ : Odrv12
    port map (
            O => \N__29220\,
            I => data_in_frame_9_6
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__29215\,
            I => data_in_frame_9_6
        );

    \I__5507\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29207\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29204\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__29204\,
            I => n17479
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__29201\,
            I => \N__29198\
        );

    \I__5503\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29194\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29197\,
            I => \N__29191\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__29194\,
            I => \N__29188\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__29191\,
            I => \N__29185\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__29188\,
            I => \N__29180\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__29185\,
            I => \N__29180\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__29180\,
            I => n9051
        );

    \I__5496\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29170\
        );

    \I__5494\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29167\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__29170\,
            I => \N__29162\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__29167\,
            I => \N__29162\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__5490\ : Odrv4
    port map (
            O => \N__29159\,
            I => n6_adj_2583
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__5488\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__5486\ : Span4Mux_s2_h
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__29141\,
            I => \c0.data_out_frame2_19_2\
        );

    \I__5483\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29135\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__29135\,
            I => \N__29130\
        );

    \I__5481\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29127\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__29133\,
            I => \N__29123\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__29130\,
            I => \N__29119\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__29127\,
            I => \N__29116\
        );

    \I__5477\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29113\
        );

    \I__5476\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29110\
        );

    \I__5475\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29107\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__29119\,
            I => \N__29102\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__29116\,
            I => \N__29102\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__29113\,
            I => \c0.data_in_frame_0_1\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__29110\,
            I => \c0.data_in_frame_0_1\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__29107\,
            I => \c0.data_in_frame_0_1\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__29102\,
            I => \c0.data_in_frame_0_1\
        );

    \I__5468\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29085\
        );

    \I__5466\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29081\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29078\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__29085\,
            I => \N__29075\
        );

    \I__5463\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29072\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__29081\,
            I => \N__29069\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__29078\,
            I => \c0.data_in_frame_3_6\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__29075\,
            I => \c0.data_in_frame_3_6\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__29072\,
            I => \c0.data_in_frame_3_6\
        );

    \I__5458\ : Odrv12
    port map (
            O => \N__29069\,
            I => \c0.data_in_frame_3_6\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__29060\,
            I => \N__29057\
        );

    \I__5456\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29053\
        );

    \I__5455\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__29050\,
            I => \N__29044\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__29047\,
            I => \N__29041\
        );

    \I__5451\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__29035\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__29041\,
            I => \N__29035\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__29040\,
            I => \N__29032\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__29035\,
            I => \N__29027\
        );

    \I__5447\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29022\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29022\
        );

    \I__5445\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29019\
        );

    \I__5444\ : Odrv4
    port map (
            O => \N__29027\,
            I => \c0.data_in_frame_2_1\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__29022\,
            I => \c0.data_in_frame_2_1\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__29019\,
            I => \c0.data_in_frame_2_1\
        );

    \I__5441\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29007\
        );

    \I__5440\ : InMux
    port map (
            O => \N__29011\,
            I => \N__29002\
        );

    \I__5439\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29002\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__29007\,
            I => \N__28998\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28995\
        );

    \I__5436\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28992\
        );

    \I__5435\ : Span12Mux_v
    port map (
            O => \N__28998\,
            I => \N__28989\
        );

    \I__5434\ : Span4Mux_h
    port map (
            O => \N__28995\,
            I => \N__28986\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__28992\,
            I => \c0.data_in_frame_0_2\
        );

    \I__5432\ : Odrv12
    port map (
            O => \N__28989\,
            I => \c0.data_in_frame_0_2\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__28986\,
            I => \c0.data_in_frame_0_2\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__28979\,
            I => \N__28975\
        );

    \I__5429\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28971\
        );

    \I__5428\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28968\
        );

    \I__5427\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__28965\,
            I => \N__28956\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__28962\,
            I => \N__28953\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__28959\,
            I => \N__28950\
        );

    \I__5421\ : Span12Mux_s8_v
    port map (
            O => \N__28956\,
            I => \N__28947\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__28953\,
            I => \N__28942\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__28950\,
            I => \N__28942\
        );

    \I__5418\ : Odrv12
    port map (
            O => \N__28947\,
            I => \c0.n9043\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__28942\,
            I => \c0.n9043\
        );

    \I__5416\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__5414\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__28930\,
            I => \N__28924\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28917\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__28921\,
            I => \N__28914\
        );

    \I__5409\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28911\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__28917\,
            I => \N__28908\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__28914\,
            I => \N__28905\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28902\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__28908\,
            I => \c0.n8886\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__28905\,
            I => \c0.n8886\
        );

    \I__5403\ : Odrv12
    port map (
            O => \N__28902\,
            I => \c0.n8886\
        );

    \I__5402\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28891\
        );

    \I__5401\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28888\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28885\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__28888\,
            I => \c0.n15927\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__28885\,
            I => \c0.n15927\
        );

    \I__5397\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__28877\,
            I => \N__28874\
        );

    \I__5395\ : Span4Mux_v
    port map (
            O => \N__28874\,
            I => \N__28870\
        );

    \I__5394\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28867\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28861\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__28864\,
            I => \N__28856\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__28861\,
            I => \N__28856\
        );

    \I__5389\ : Sp12to4
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__5388\ : Odrv12
    port map (
            O => \N__28853\,
            I => \c0.n17594\
        );

    \I__5387\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28846\
        );

    \I__5386\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28843\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__28846\,
            I => \N__28840\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__28843\,
            I => \N__28837\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__28840\,
            I => \N__28832\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__28837\,
            I => \N__28832\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__28832\,
            I => \c0.n17412\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__28829\,
            I => \n2565_cascade_\
        );

    \I__5379\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__28820\,
            I => \N__28816\
        );

    \I__5376\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28813\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__28816\,
            I => n2574
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__28813\,
            I => n2574
        );

    \I__5373\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28804\
        );

    \I__5372\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28801\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__28804\,
            I => \N__28798\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28795\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__28798\,
            I => n17547
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__28795\,
            I => n17547
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__28790\,
            I => \c0.n23_cascade_\
        );

    \I__5366\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28784\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__28784\,
            I => \c0.n17536\
        );

    \I__5364\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28778\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__28778\,
            I => \c0.n28\
        );

    \I__5362\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28768\
        );

    \I__5361\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28768\
        );

    \I__5360\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28764\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28761\
        );

    \I__5358\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28756\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__28764\,
            I => \N__28753\
        );

    \I__5356\ : Span12Mux_v
    port map (
            O => \N__28761\,
            I => \N__28750\
        );

    \I__5355\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28745\
        );

    \I__5354\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28745\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__28756\,
            I => \N__28740\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__28753\,
            I => \N__28740\
        );

    \I__5351\ : Odrv12
    port map (
            O => \N__28750\,
            I => data_in_frame_8_0
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__28745\,
            I => data_in_frame_8_0
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__28740\,
            I => data_in_frame_8_0
        );

    \I__5348\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28727\
        );

    \I__5347\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28727\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__28724\,
            I => \N__28720\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__28723\,
            I => \N__28717\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__28720\,
            I => \N__28711\
        );

    \I__5342\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28706\
        );

    \I__5341\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28706\
        );

    \I__5340\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28701\
        );

    \I__5339\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28701\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__28711\,
            I => data_in_frame_1_1
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__28706\,
            I => data_in_frame_1_1
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__28701\,
            I => data_in_frame_1_1
        );

    \I__5335\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28689\
        );

    \I__5334\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28686\
        );

    \I__5333\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28683\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__28689\,
            I => \N__28680\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__28686\,
            I => \N__28672\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__28683\,
            I => \N__28672\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__28680\,
            I => \N__28672\
        );

    \I__5328\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28669\
        );

    \I__5327\ : Span4Mux_v
    port map (
            O => \N__28672\,
            I => \N__28664\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28664\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__28661\,
            I => \c0.data_in_frame_10_4\
        );

    \I__5323\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28649\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__28649\,
            I => n2563
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__28646\,
            I => \N__28642\
        );

    \I__5318\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28638\
        );

    \I__5317\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28635\
        );

    \I__5316\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28632\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28628\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__28635\,
            I => \N__28625\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__28632\,
            I => \N__28622\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__28631\,
            I => \N__28618\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__28628\,
            I => \N__28615\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__28625\,
            I => \N__28610\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__28622\,
            I => \N__28610\
        );

    \I__5308\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28607\
        );

    \I__5307\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28604\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__28615\,
            I => \c0.data_in_frame_7_2\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__28610\,
            I => \c0.data_in_frame_7_2\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__28607\,
            I => \c0.data_in_frame_7_2\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__28604\,
            I => \c0.data_in_frame_7_2\
        );

    \I__5302\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__28592\,
            I => \N__28588\
        );

    \I__5300\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28585\
        );

    \I__5299\ : Span4Mux_h
    port map (
            O => \N__28588\,
            I => \N__28582\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28579\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__28582\,
            I => \N__28576\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__28579\,
            I => \N__28573\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__28576\,
            I => \c0.n8062\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__28573\,
            I => \c0.n8062\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__28568\,
            I => \n2563_cascade_\
        );

    \I__5292\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28560\
        );

    \I__5291\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28557\
        );

    \I__5290\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28554\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28551\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__28557\,
            I => \N__28546\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28546\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__28551\,
            I => \N__28541\
        );

    \I__5285\ : Span4Mux_h
    port map (
            O => \N__28546\,
            I => \N__28541\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__28541\,
            I => \N__28538\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__28538\,
            I => \c0.n9204\
        );

    \I__5282\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28531\
        );

    \I__5281\ : InMux
    port map (
            O => \N__28534\,
            I => \N__28527\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__28531\,
            I => \N__28524\
        );

    \I__5279\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28521\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__28527\,
            I => \N__28518\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__28524\,
            I => \N__28513\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__28521\,
            I => \N__28513\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__28518\,
            I => \N__28510\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__28513\,
            I => \N__28507\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__28510\,
            I => \c0.n8890\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__28507\,
            I => \c0.n8890\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__28502\,
            I => \c0.n17592_cascade_\
        );

    \I__5270\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28496\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__28496\,
            I => \c0.n26\
        );

    \I__5268\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28488\
        );

    \I__5267\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28485\
        );

    \I__5266\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28482\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28478\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__28485\,
            I => \N__28473\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__28482\,
            I => \N__28470\
        );

    \I__5262\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28467\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__28478\,
            I => \N__28464\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28459\
        );

    \I__5259\ : InMux
    port map (
            O => \N__28476\,
            I => \N__28459\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__28473\,
            I => \N__28454\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__28470\,
            I => \N__28454\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__28467\,
            I => \N__28451\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__28464\,
            I => \N__28446\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28446\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__28454\,
            I => \c0.data_in_frame_7_5\
        );

    \I__5252\ : Odrv12
    port map (
            O => \N__28451\,
            I => \c0.data_in_frame_7_5\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__28446\,
            I => \c0.data_in_frame_7_5\
        );

    \I__5250\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28435\
        );

    \I__5249\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28429\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28426\
        );

    \I__5247\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28423\
        );

    \I__5246\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28420\
        );

    \I__5245\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28417\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__28429\,
            I => \N__28412\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__28426\,
            I => \N__28412\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28409\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__28420\,
            I => \N__28404\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28404\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__28412\,
            I => data_in_frame_8_6
        );

    \I__5238\ : Odrv12
    port map (
            O => \N__28409\,
            I => data_in_frame_8_6
        );

    \I__5237\ : Odrv12
    port map (
            O => \N__28404\,
            I => data_in_frame_8_6
        );

    \I__5236\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__28394\,
            I => \N__28391\
        );

    \I__5234\ : Span4Mux_v
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__28388\,
            I => \c0.n17473\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__28385\,
            I => \N__28381\
        );

    \I__5231\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__5230\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28375\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28372\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28369\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__28372\,
            I => \N__28366\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__28369\,
            I => \N__28362\
        );

    \I__5225\ : Span4Mux_v
    port map (
            O => \N__28366\,
            I => \N__28359\
        );

    \I__5224\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28356\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__28362\,
            I => \N__28353\
        );

    \I__5222\ : Span4Mux_v
    port map (
            O => \N__28359\,
            I => \N__28350\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__28356\,
            I => \c0.data_in_4_6\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__28353\,
            I => \c0.data_in_4_6\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__28350\,
            I => \c0.data_in_4_6\
        );

    \I__5218\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28336\
        );

    \I__5217\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28332\
        );

    \I__5216\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28329\
        );

    \I__5215\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28326\
        );

    \I__5214\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28323\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28320\
        );

    \I__5212\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28317\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__28332\,
            I => \N__28312\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__28329\,
            I => \N__28305\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28305\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__28323\,
            I => \N__28305\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__28320\,
            I => \N__28300\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__28317\,
            I => \N__28300\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28297\
        );

    \I__5204\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28294\
        );

    \I__5203\ : Span12Mux_h
    port map (
            O => \N__28312\,
            I => \N__28291\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__28305\,
            I => \N__28286\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__28300\,
            I => \N__28286\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28283\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__28294\,
            I => data_in_frame_5_7
        );

    \I__5198\ : Odrv12
    port map (
            O => \N__28291\,
            I => data_in_frame_5_7
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__28286\,
            I => data_in_frame_5_7
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__28283\,
            I => data_in_frame_5_7
        );

    \I__5195\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__5193\ : Span4Mux_v
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__28265\,
            I => \c0.n9368\
        );

    \I__5191\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28258\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__28261\,
            I => \N__28255\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__28258\,
            I => \N__28251\
        );

    \I__5188\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28248\
        );

    \I__5187\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28245\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__28251\,
            I => \N__28242\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28239\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28236\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__28242\,
            I => \N__28233\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__28239\,
            I => \N__28230\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__28236\,
            I => \N__28227\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__28233\,
            I => \c0.n9365\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__28230\,
            I => \c0.n9365\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__28227\,
            I => \c0.n9365\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__28220\,
            I => \c0.n2600_cascade_\
        );

    \I__5176\ : InMux
    port map (
            O => \N__28217\,
            I => \N__28213\
        );

    \I__5175\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28210\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28207\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28204\
        );

    \I__5172\ : Span4Mux_s2_h
    port map (
            O => \N__28207\,
            I => \N__28199\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__28204\,
            I => \N__28199\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__28199\,
            I => \c0.n9334\
        );

    \I__5169\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28193\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__28193\,
            I => \c0.n10_adj_2493\
        );

    \I__5167\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__28184\,
            I => \N__28178\
        );

    \I__5164\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28175\
        );

    \I__5163\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28171\
        );

    \I__5162\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28168\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__28178\,
            I => \N__28165\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__28175\,
            I => \N__28162\
        );

    \I__5159\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28159\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__28171\,
            I => data_in_3_6
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__28168\,
            I => data_in_3_6
        );

    \I__5156\ : Odrv4
    port map (
            O => \N__28165\,
            I => data_in_3_6
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__28162\,
            I => data_in_3_6
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__28159\,
            I => data_in_3_6
        );

    \I__5153\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__28145\,
            I => \N__28138\
        );

    \I__5151\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28131\
        );

    \I__5150\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28131\
        );

    \I__5149\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28131\
        );

    \I__5148\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28128\
        );

    \I__5147\ : Span4Mux_v
    port map (
            O => \N__28138\,
            I => \N__28125\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__28131\,
            I => data_in_1_2
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__28128\,
            I => data_in_1_2
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__28125\,
            I => data_in_1_2
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__28118\,
            I => \N__28114\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__28117\,
            I => \N__28111\
        );

    \I__5141\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28108\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__28108\,
            I => \c0.n8572\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__28105\,
            I => \c0.n8572\
        );

    \I__5137\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28095\
        );

    \I__5136\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28089\
        );

    \I__5135\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28089\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28086\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28083\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__28089\,
            I => \N__28080\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__28086\,
            I => \N__28077\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28072\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__28080\,
            I => \N__28072\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__28077\,
            I => data_in_frame_6_5
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__28072\,
            I => data_in_frame_6_5
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28063\
        );

    \I__5125\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28059\
        );

    \I__5124\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28053\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28053\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__28059\,
            I => \N__28049\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28046\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28039\
        );

    \I__5119\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28036\
        );

    \I__5118\ : Span4Mux_s3_h
    port map (
            O => \N__28049\,
            I => \N__28028\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28028\
        );

    \I__5116\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28025\
        );

    \I__5115\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28016\
        );

    \I__5114\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28016\
        );

    \I__5113\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28016\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__28039\,
            I => \N__28013\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28010\
        );

    \I__5110\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28001\
        );

    \I__5109\ : InMux
    port map (
            O => \N__28034\,
            I => \N__27998\
        );

    \I__5108\ : InMux
    port map (
            O => \N__28033\,
            I => \N__27995\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__28028\,
            I => \N__27990\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28025\,
            I => \N__27990\
        );

    \I__5105\ : InMux
    port map (
            O => \N__28024\,
            I => \N__27985\
        );

    \I__5104\ : InMux
    port map (
            O => \N__28023\,
            I => \N__27985\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__27978\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__28013\,
            I => \N__27978\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__27978\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28009\,
            I => \N__27971\
        );

    \I__5099\ : InMux
    port map (
            O => \N__28008\,
            I => \N__27971\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28007\,
            I => \N__27971\
        );

    \I__5097\ : InMux
    port map (
            O => \N__28006\,
            I => \N__27964\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27964\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27964\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__28001\,
            I => \c0.n4_adj_2512\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__27998\,
            I => \c0.n4_adj_2512\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__27995\,
            I => \c0.n4_adj_2512\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__27990\,
            I => \c0.n4_adj_2512\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__27985\,
            I => \c0.n4_adj_2512\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__27978\,
            I => \c0.n4_adj_2512\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__27971\,
            I => \c0.n4_adj_2512\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__27964\,
            I => \c0.n4_adj_2512\
        );

    \I__5086\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27943\
        );

    \I__5085\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27939\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__27943\,
            I => \N__27936\
        );

    \I__5083\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27933\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27930\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__27936\,
            I => \N__27925\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27925\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__27930\,
            I => \N__27922\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__27925\,
            I => n2594
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__27922\,
            I => n2594
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__27917\,
            I => \n2573_cascade_\
        );

    \I__5075\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27911\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__27911\,
            I => n17481
        );

    \I__5073\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27905\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__27905\,
            I => \N__27901\
        );

    \I__5071\ : InMux
    port map (
            O => \N__27904\,
            I => \N__27898\
        );

    \I__5070\ : Span4Mux_h
    port map (
            O => \N__27901\,
            I => \N__27890\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__27898\,
            I => \N__27890\
        );

    \I__5068\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27885\
        );

    \I__5067\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27885\
        );

    \I__5066\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27882\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__27890\,
            I => \N__27877\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__27885\,
            I => \N__27877\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__27882\,
            I => \c0.data_in_3_4\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__27877\,
            I => \c0.data_in_3_4\
        );

    \I__5061\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27869\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__27869\,
            I => \c0.n17743\
        );

    \I__5059\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27862\
        );

    \I__5058\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27859\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__27862\,
            I => \N__27856\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__27859\,
            I => \N__27851\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__27856\,
            I => \N__27851\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__27851\,
            I => \N__27847\
        );

    \I__5053\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27844\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__27847\,
            I => data_in_4_0
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__27844\,
            I => data_in_4_0
        );

    \I__5050\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__27836\,
            I => \N__27832\
        );

    \I__5048\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27828\
        );

    \I__5047\ : Span4Mux_s3_h
    port map (
            O => \N__27832\,
            I => \N__27825\
        );

    \I__5046\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27820\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27817\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__27825\,
            I => \N__27814\
        );

    \I__5043\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27811\
        );

    \I__5042\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27808\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__27820\,
            I => \c0.data_in_3_0\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__27817\,
            I => \c0.data_in_3_0\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__27814\,
            I => \c0.data_in_3_0\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__27811\,
            I => \c0.data_in_3_0\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__27808\,
            I => \c0.data_in_3_0\
        );

    \I__5036\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27793\
        );

    \I__5035\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27786\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__27790\,
            I => \N__27783\
        );

    \I__5032\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27779\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__27786\,
            I => \N__27773\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__27783\,
            I => \N__27773\
        );

    \I__5029\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27770\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27767\
        );

    \I__5027\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27764\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__27773\,
            I => \N__27761\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__27770\,
            I => \N__27756\
        );

    \I__5024\ : Span12Mux_v
    port map (
            O => \N__27767\,
            I => \N__27756\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__27764\,
            I => data_in_1_6
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__27761\,
            I => data_in_1_6
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__27756\,
            I => data_in_1_6
        );

    \I__5020\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27746\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__27746\,
            I => \N__27743\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__27743\,
            I => \N__27737\
        );

    \I__5017\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27734\
        );

    \I__5016\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27731\
        );

    \I__5015\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27728\
        );

    \I__5014\ : Odrv4
    port map (
            O => \N__27737\,
            I => data_in_0_6
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__27734\,
            I => data_in_0_6
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__27731\,
            I => data_in_0_6
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__27728\,
            I => data_in_0_6
        );

    \I__5010\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27715\
        );

    \I__5009\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27711\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27708\
        );

    \I__5007\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27704\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__27711\,
            I => \N__27699\
        );

    \I__5005\ : Span12Mux_v
    port map (
            O => \N__27708\,
            I => \N__27699\
        );

    \I__5004\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27696\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__27704\,
            I => data_in_2_6
        );

    \I__5002\ : Odrv12
    port map (
            O => \N__27699\,
            I => data_in_2_6
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__27696\,
            I => data_in_2_6
        );

    \I__5000\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27683\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__27683\,
            I => \N__27677\
        );

    \I__4997\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27672\
        );

    \I__4996\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__4995\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27669\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__27677\,
            I => data_in_3_1
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__27672\,
            I => data_in_3_1
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__27669\,
            I => data_in_3_1
        );

    \I__4991\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27659\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__27659\,
            I => \N__27654\
        );

    \I__4989\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27649\
        );

    \I__4988\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27649\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__27654\,
            I => data_in_9_1
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__27649\,
            I => data_in_9_1
        );

    \I__4985\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27640\
        );

    \I__4984\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__27640\,
            I => \N__27634\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__27637\,
            I => \N__27631\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__27634\,
            I => \N__27626\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__27631\,
            I => \N__27623\
        );

    \I__4979\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27618\
        );

    \I__4978\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27618\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__27626\,
            I => \c0.data_in_1_3\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__27623\,
            I => \c0.data_in_1_3\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__27618\,
            I => \c0.data_in_1_3\
        );

    \I__4974\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__4972\ : Span4Mux_s2_h
    port map (
            O => \N__27605\,
            I => \N__27601\
        );

    \I__4971\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27598\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__27601\,
            I => \N__27593\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27590\
        );

    \I__4968\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27585\
        );

    \I__4967\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27585\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__27593\,
            I => \c0.data_in_0_3\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__27590\,
            I => \c0.data_in_0_3\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__27585\,
            I => \c0.data_in_0_3\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__27578\,
            I => \N__27575\
        );

    \I__4962\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27568\
        );

    \I__4960\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__27568\,
            I => \N__27561\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27558\
        );

    \I__4957\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27555\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__27561\,
            I => data_in_4_3
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__27558\,
            I => data_in_4_3
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__27555\,
            I => data_in_4_3
        );

    \I__4953\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4951\ : Span4Mux_s2_h
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__27539\,
            I => \N__27533\
        );

    \I__4949\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27528\
        );

    \I__4948\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27528\
        );

    \I__4947\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27525\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__27533\,
            I => data_in_3_3
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__27528\,
            I => data_in_3_3
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__27525\,
            I => data_in_3_3
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__27518\,
            I => \N__27513\
        );

    \I__4942\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27510\
        );

    \I__4941\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27506\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27503\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__27510\,
            I => \N__27500\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27497\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27494\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27491\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__27500\,
            I => \N__27486\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__27497\,
            I => \N__27486\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__27494\,
            I => \N__27481\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__27491\,
            I => \N__27481\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__27486\,
            I => \N__27478\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__27481\,
            I => \c0.data_in_frame_7_4\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__27478\,
            I => \c0.data_in_frame_7_4\
        );

    \I__4928\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27470\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__27467\,
            I => \N__27463\
        );

    \I__4925\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27460\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__27463\,
            I => n2587
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__27460\,
            I => n2587
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__27455\,
            I => \N__27450\
        );

    \I__4921\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27447\
        );

    \I__4920\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27442\
        );

    \I__4919\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27442\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__27447\,
            I => \c0.data_in_7_4\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__27442\,
            I => \c0.data_in_7_4\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__27437\,
            I => \N__27434\
        );

    \I__4915\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27431\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__27428\,
            I => \N__27423\
        );

    \I__4912\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27420\
        );

    \I__4911\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27417\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__27423\,
            I => \N__27414\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__27420\,
            I => \c0.data_in_6_4\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__27417\,
            I => \c0.data_in_6_4\
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__27414\,
            I => \c0.data_in_6_4\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__27407\,
            I => \N__27404\
        );

    \I__4905\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27400\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__27403\,
            I => \N__27397\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27394\
        );

    \I__4902\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27391\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__27394\,
            I => \N__27384\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27384\
        );

    \I__4899\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27379\
        );

    \I__4898\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27379\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__27384\,
            I => \N__27376\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__27379\,
            I => data_in_5_4
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__27376\,
            I => data_in_5_4
        );

    \I__4894\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__27365\,
            I => \N__27361\
        );

    \I__4891\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27358\
        );

    \I__4890\ : Span4Mux_s3_h
    port map (
            O => \N__27361\,
            I => \N__27354\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__27358\,
            I => \N__27351\
        );

    \I__4888\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27348\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__27354\,
            I => \c0.data_in_4_4\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__27351\,
            I => \c0.data_in_4_4\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__27348\,
            I => \c0.data_in_4_4\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__27338\,
            I => \N__27335\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__27335\,
            I => \N__27332\
        );

    \I__4881\ : Span4Mux_v
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__27329\,
            I => n17952
        );

    \I__4879\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27322\
        );

    \I__4878\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27319\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27316\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__27319\,
            I => \N__27311\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__27316\,
            I => \N__27308\
        );

    \I__4874\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27305\
        );

    \I__4873\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27302\
        );

    \I__4872\ : Sp12to4
    port map (
            O => \N__27311\,
            I => \N__27299\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__27308\,
            I => \N__27296\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27293\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__27302\,
            I => data_in_2_4
        );

    \I__4868\ : Odrv12
    port map (
            O => \N__27299\,
            I => data_in_2_4
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__27296\,
            I => data_in_2_4
        );

    \I__4866\ : Odrv12
    port map (
            O => \N__27293\,
            I => data_in_2_4
        );

    \I__4865\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27277\
        );

    \I__4863\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27272\
        );

    \I__4862\ : Span4Mux_v
    port map (
            O => \N__27277\,
            I => \N__27268\
        );

    \I__4861\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27265\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27262\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27259\
        );

    \I__4858\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27256\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__27268\,
            I => data_in_2_7
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__27265\,
            I => data_in_2_7
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__27262\,
            I => data_in_2_7
        );

    \I__4854\ : Odrv12
    port map (
            O => \N__27259\,
            I => data_in_2_7
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__27256\,
            I => data_in_2_7
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__4851\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__27233\,
            I => \N__27228\
        );

    \I__4847\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27225\
        );

    \I__4846\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27222\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__27228\,
            I => data_in_4_7
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__27225\,
            I => data_in_4_7
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__27222\,
            I => data_in_4_7
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4841\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__27209\,
            I => \N__27206\
        );

    \I__4839\ : Span4Mux_s3_h
    port map (
            O => \N__27206\,
            I => \N__27203\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__27200\,
            I => \N__27195\
        );

    \I__4836\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27192\
        );

    \I__4835\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27189\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__27195\,
            I => data_in_4_5
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27192\,
            I => data_in_4_5
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__27189\,
            I => data_in_4_5
        );

    \I__4831\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27179\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27176\
        );

    \I__4829\ : Span4Mux_v
    port map (
            O => \N__27176\,
            I => \N__27169\
        );

    \I__4828\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__4827\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27161\
        );

    \I__4826\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27161\
        );

    \I__4825\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27158\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__27169\,
            I => data_in_3_5
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__27166\,
            I => data_in_3_5
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__27161\,
            I => data_in_3_5
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__27158\,
            I => data_in_3_5
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__27149\,
            I => \c0.n28_adj_2475_cascade_\
        );

    \I__4819\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__27143\,
            I => \c0.n8_adj_2474\
        );

    \I__4817\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__27134\,
            I => \N__27130\
        );

    \I__4814\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27127\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__27130\,
            I => \c0.n8559\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__27127\,
            I => \c0.n8559\
        );

    \I__4811\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27119\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__4809\ : Span4Mux_v
    port map (
            O => \N__27116\,
            I => \N__27112\
        );

    \I__4808\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27108\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__27112\,
            I => \N__27105\
        );

    \I__4806\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27100\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27097\
        );

    \I__4804\ : Sp12to4
    port map (
            O => \N__27105\,
            I => \N__27094\
        );

    \I__4803\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27091\
        );

    \I__4802\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27088\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__27100\,
            I => \c0.data_in_2_0\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__27097\,
            I => \c0.data_in_2_0\
        );

    \I__4799\ : Odrv12
    port map (
            O => \N__27094\,
            I => \c0.data_in_2_0\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__27091\,
            I => \c0.data_in_2_0\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27088\,
            I => \c0.data_in_2_0\
        );

    \I__4796\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27070\
        );

    \I__4794\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27067\
        );

    \I__4793\ : Span4Mux_s3_h
    port map (
            O => \N__27070\,
            I => \N__27064\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__27067\,
            I => \N__27059\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__27064\,
            I => \N__27056\
        );

    \I__4790\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27053\
        );

    \I__4789\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27050\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__27059\,
            I => data_in_0_1
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__27056\,
            I => data_in_0_1
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27053\,
            I => data_in_0_1
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__27050\,
            I => data_in_0_1
        );

    \I__4784\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27034\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27037\,
            I => \N__27029\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__27034\,
            I => \N__27026\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__27033\,
            I => \N__27023\
        );

    \I__4779\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27019\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__27029\,
            I => \N__27016\
        );

    \I__4777\ : Span4Mux_h
    port map (
            O => \N__27026\,
            I => \N__27013\
        );

    \I__4776\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27010\
        );

    \I__4775\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27007\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__27019\,
            I => data_in_1_7
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__27016\,
            I => data_in_1_7
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__27013\,
            I => data_in_1_7
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__27010\,
            I => data_in_1_7
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__27007\,
            I => data_in_1_7
        );

    \I__4769\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__26990\,
            I => \N__26986\
        );

    \I__4766\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26982\
        );

    \I__4765\ : Span4Mux_s2_h
    port map (
            O => \N__26986\,
            I => \N__26979\
        );

    \I__4764\ : InMux
    port map (
            O => \N__26985\,
            I => \N__26974\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__26982\,
            I => \N__26971\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__26979\,
            I => \N__26968\
        );

    \I__4761\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26965\
        );

    \I__4760\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26962\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__26974\,
            I => data_in_2_5
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__26971\,
            I => data_in_2_5
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__26968\,
            I => data_in_2_5
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__26965\,
            I => data_in_2_5
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__26962\,
            I => data_in_2_5
        );

    \I__4754\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26948\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__26945\,
            I => \c0.n17_adj_2486\
        );

    \I__4751\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26938\
        );

    \I__4750\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26935\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26930\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26926\
        );

    \I__4747\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26922\
        );

    \I__4746\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26919\
        );

    \I__4745\ : Span4Mux_v
    port map (
            O => \N__26930\,
            I => \N__26916\
        );

    \I__4744\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26913\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__26926\,
            I => \N__26910\
        );

    \I__4742\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26907\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__26922\,
            I => \N__26902\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__26919\,
            I => \N__26895\
        );

    \I__4739\ : Span4Mux_s1_h
    port map (
            O => \N__26916\,
            I => \N__26895\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__26913\,
            I => \N__26895\
        );

    \I__4737\ : Sp12to4
    port map (
            O => \N__26910\,
            I => \N__26890\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26890\
        );

    \I__4735\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26887\
        );

    \I__4734\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26884\
        );

    \I__4733\ : Span4Mux_v
    port map (
            O => \N__26902\,
            I => \N__26879\
        );

    \I__4732\ : Span4Mux_v
    port map (
            O => \N__26895\,
            I => \N__26879\
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__26890\,
            I => \c0.n134\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__26887\,
            I => \c0.n134\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__26884\,
            I => \c0.n134\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__26879\,
            I => \c0.n134\
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__26870\,
            I => \c0.n18531_cascade_\
        );

    \I__4726\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26864\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26860\
        );

    \I__4724\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26857\
        );

    \I__4723\ : Span4Mux_s2_v
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__26857\,
            I => data_out_frame2_5_4
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__26854\,
            I => data_out_frame2_5_4
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__26849\,
            I => \c0.n17955_cascade_\
        );

    \I__4719\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26835\
        );

    \I__4718\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26835\
        );

    \I__4717\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26828\
        );

    \I__4716\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26828\
        );

    \I__4715\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26823\
        );

    \I__4714\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26818\
        );

    \I__4713\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26818\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N__26815\
        );

    \I__4711\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26812\
        );

    \I__4710\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26809\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26806\
        );

    \I__4708\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26801\
        );

    \I__4707\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26801\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26795\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__26818\,
            I => \N__26786\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__26815\,
            I => \N__26786\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__26812\,
            I => \N__26786\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__26809\,
            I => \N__26786\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__26806\,
            I => \N__26775\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26775\
        );

    \I__4699\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26768\
        );

    \I__4698\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26768\
        );

    \I__4697\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26768\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__26795\,
            I => \N__26765\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__26786\,
            I => \N__26762\
        );

    \I__4694\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26759\
        );

    \I__4693\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26755\
        );

    \I__4692\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26750\
        );

    \I__4691\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26750\
        );

    \I__4690\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26745\
        );

    \I__4689\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26745\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__26775\,
            I => \N__26742\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__26768\,
            I => \N__26733\
        );

    \I__4686\ : Sp12to4
    port map (
            O => \N__26765\,
            I => \N__26733\
        );

    \I__4685\ : Sp12to4
    port map (
            O => \N__26762\,
            I => \N__26733\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__26759\,
            I => \N__26733\
        );

    \I__4683\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26730\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__26755\,
            I => \N__26719\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__26750\,
            I => \N__26719\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__26745\,
            I => \N__26719\
        );

    \I__4679\ : Sp12to4
    port map (
            O => \N__26742\,
            I => \N__26719\
        );

    \I__4678\ : Span12Mux_h
    port map (
            O => \N__26733\,
            I => \N__26719\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__26730\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__4676\ : Odrv12
    port map (
            O => \N__26719\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__4675\ : InMux
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__26711\,
            I => \N__26707\
        );

    \I__4673\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26704\
        );

    \I__4672\ : Span4Mux_s2_v
    port map (
            O => \N__26707\,
            I => \N__26701\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__26704\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__26701\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \c0.n18456_cascade_\
        );

    \I__4668\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__26690\,
            I => \c0.n18447\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__26687\,
            I => \c0.n18459_cascade_\
        );

    \I__4665\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__26681\,
            I => \c0.n22_adj_2525\
        );

    \I__4663\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26669\
        );

    \I__4662\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26654\
        );

    \I__4661\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26654\
        );

    \I__4660\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26654\
        );

    \I__4659\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26647\
        );

    \I__4658\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26647\
        );

    \I__4657\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26647\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26644\
        );

    \I__4655\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26641\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__26667\,
            I => \N__26638\
        );

    \I__4653\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26635\
        );

    \I__4652\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26628\
        );

    \I__4651\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26628\
        );

    \I__4650\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26628\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__26662\,
            I => \N__26621\
        );

    \I__4648\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26613\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__26654\,
            I => \N__26608\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__26647\,
            I => \N__26608\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__26644\,
            I => \N__26603\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26603\
        );

    \I__4643\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26599\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26594\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__26628\,
            I => \N__26594\
        );

    \I__4640\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26589\
        );

    \I__4639\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26589\
        );

    \I__4638\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26584\
        );

    \I__4637\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26584\
        );

    \I__4636\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26581\
        );

    \I__4635\ : InMux
    port map (
            O => \N__26620\,
            I => \N__26576\
        );

    \I__4634\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26576\
        );

    \I__4633\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26569\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26569\
        );

    \I__4631\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26569\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26564\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__26608\,
            I => \N__26564\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__26603\,
            I => \N__26561\
        );

    \I__4627\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26558\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__26599\,
            I => \N__26555\
        );

    \I__4625\ : Span12Mux_s10_v
    port map (
            O => \N__26594\,
            I => \N__26552\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__26589\,
            I => \N__26537\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26537\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26537\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__26576\,
            I => \N__26537\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26537\
        );

    \I__4619\ : Sp12to4
    port map (
            O => \N__26564\,
            I => \N__26537\
        );

    \I__4618\ : Sp12to4
    port map (
            O => \N__26561\,
            I => \N__26537\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__26558\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__26555\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__4615\ : Odrv12
    port map (
            O => \N__26552\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__4614\ : Odrv12
    port map (
            O => \N__26537\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__26528\,
            I => \c0.n15_cascade_\
        );

    \I__4612\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26522\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26515\
        );

    \I__4610\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26512\
        );

    \I__4609\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26509\
        );

    \I__4608\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26505\
        );

    \I__4607\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26502\
        );

    \I__4606\ : Span4Mux_s2_v
    port map (
            O => \N__26515\,
            I => \N__26495\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__26512\,
            I => \N__26495\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__26509\,
            I => \N__26492\
        );

    \I__4603\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26489\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26486\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26483\
        );

    \I__4600\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26480\
        );

    \I__4599\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26477\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__26495\,
            I => \N__26473\
        );

    \I__4597\ : Span4Mux_h
    port map (
            O => \N__26492\,
            I => \N__26466\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__26489\,
            I => \N__26466\
        );

    \I__4595\ : Span4Mux_s2_v
    port map (
            O => \N__26486\,
            I => \N__26466\
        );

    \I__4594\ : Span4Mux_s3_v
    port map (
            O => \N__26483\,
            I => \N__26459\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26459\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26459\
        );

    \I__4591\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26456\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__26473\,
            I => \N__26450\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__26466\,
            I => \N__26450\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__26459\,
            I => \N__26445\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__26456\,
            I => \N__26445\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26442\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__26450\,
            I => \N__26439\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__26445\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__26442\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__26439\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__4580\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__26420\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__4576\ : CEMux
    port map (
            O => \N__26417\,
            I => \N__26413\
        );

    \I__4575\ : CEMux
    port map (
            O => \N__26416\,
            I => \N__26410\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26406\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26401\
        );

    \I__4572\ : CEMux
    port map (
            O => \N__26409\,
            I => \N__26397\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__26406\,
            I => \N__26394\
        );

    \I__4570\ : CEMux
    port map (
            O => \N__26405\,
            I => \N__26391\
        );

    \I__4569\ : CEMux
    port map (
            O => \N__26404\,
            I => \N__26388\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__26401\,
            I => \N__26385\
        );

    \I__4567\ : CEMux
    port map (
            O => \N__26400\,
            I => \N__26382\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__26397\,
            I => \N__26379\
        );

    \I__4565\ : Sp12to4
    port map (
            O => \N__26394\,
            I => \N__26374\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__26391\,
            I => \N__26371\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26368\
        );

    \I__4562\ : Span4Mux_h
    port map (
            O => \N__26385\,
            I => \N__26365\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__26382\,
            I => \N__26362\
        );

    \I__4560\ : Span4Mux_s2_h
    port map (
            O => \N__26379\,
            I => \N__26359\
        );

    \I__4559\ : CEMux
    port map (
            O => \N__26378\,
            I => \N__26356\
        );

    \I__4558\ : CEMux
    port map (
            O => \N__26377\,
            I => \N__26353\
        );

    \I__4557\ : Span12Mux_s1_h
    port map (
            O => \N__26374\,
            I => \N__26350\
        );

    \I__4556\ : Span4Mux_v
    port map (
            O => \N__26371\,
            I => \N__26347\
        );

    \I__4555\ : Span4Mux_s1_v
    port map (
            O => \N__26368\,
            I => \N__26344\
        );

    \I__4554\ : Span4Mux_s1_h
    port map (
            O => \N__26365\,
            I => \N__26341\
        );

    \I__4553\ : Sp12to4
    port map (
            O => \N__26362\,
            I => \N__26338\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__26359\,
            I => \N__26335\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__26356\,
            I => \c0.tx2.n7727\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__26353\,
            I => \c0.tx2.n7727\
        );

    \I__4549\ : Odrv12
    port map (
            O => \N__26350\,
            I => \c0.tx2.n7727\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__26347\,
            I => \c0.tx2.n7727\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__26344\,
            I => \c0.tx2.n7727\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__26341\,
            I => \c0.tx2.n7727\
        );

    \I__4545\ : Odrv12
    port map (
            O => \N__26338\,
            I => \c0.tx2.n7727\
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__26335\,
            I => \c0.tx2.n7727\
        );

    \I__4543\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26315\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__4541\ : Span4Mux_s2_v
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__26309\,
            I => n224
        );

    \I__4539\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__26303\,
            I => n226
        );

    \I__4537\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__26297\,
            I => n221
        );

    \I__4535\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__26291\,
            I => n223
        );

    \I__4533\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__26285\,
            I => \c0.rx.n17999\
        );

    \I__4531\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__26276\,
            I => \c0.n18444\
        );

    \I__4528\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__26267\,
            I => \c0.n9\
        );

    \I__4525\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26257\
        );

    \I__4523\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26254\
        );

    \I__4522\ : Span4Mux_h
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26246\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__26251\,
            I => \N__26246\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__26246\,
            I => data_out_frame2_18_4
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__4517\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26237\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__4515\ : Span4Mux_v
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__26231\,
            I => \N__26228\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__26228\,
            I => \c0.data_out_frame2_19_4\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26218\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26215\
        );

    \I__4509\ : Span4Mux_s3_v
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__26215\,
            I => data_out_frame2_16_4
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__26212\,
            I => data_out_frame2_16_4
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__26207\,
            I => \c0.n18528_cascade_\
        );

    \I__4505\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26197\
        );

    \I__4503\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26194\
        );

    \I__4502\ : Span12Mux_s6_v
    port map (
            O => \N__26197\,
            I => \N__26191\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__26194\,
            I => data_out_frame2_17_4
        );

    \I__4500\ : Odrv12
    port map (
            O => \N__26191\,
            I => data_out_frame2_17_4
        );

    \I__4499\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26182\
        );

    \I__4498\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26177\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__26182\,
            I => \N__26174\
        );

    \I__4496\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26171\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26164\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26161\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__26174\,
            I => \N__26156\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26156\
        );

    \I__4491\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26153\
        );

    \I__4490\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26144\
        );

    \I__4489\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26144\
        );

    \I__4488\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26144\
        );

    \I__4487\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26144\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__26161\,
            I => \r_Bit_Index_1_adj_2636\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__26156\,
            I => \r_Bit_Index_1_adj_2636\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__26153\,
            I => \r_Bit_Index_1_adj_2636\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__26144\,
            I => \r_Bit_Index_1_adj_2636\
        );

    \I__4482\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26132\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__4480\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26121\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26121\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__26129\,
            I => \N__26115\
        );

    \I__4477\ : Span4Mux_h
    port map (
            O => \N__26126\,
            I => \N__26110\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26110\
        );

    \I__4475\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26103\
        );

    \I__4474\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26103\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26103\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26100\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__26110\,
            I => \r_Bit_Index_0_adj_2637\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__26103\,
            I => \r_Bit_Index_0_adj_2637\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__26100\,
            I => \r_Bit_Index_0_adj_2637\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__4467\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__26087\,
            I => n4980
        );

    \I__4465\ : InMux
    port map (
            O => \N__26084\,
            I => \bfn_6_30_0_\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26078\,
            I => n225
        );

    \I__4462\ : InMux
    port map (
            O => \N__26075\,
            I => \c0.rx.n16365\
        );

    \I__4461\ : InMux
    port map (
            O => \N__26072\,
            I => \c0.rx.n16366\
        );

    \I__4460\ : InMux
    port map (
            O => \N__26069\,
            I => \c0.rx.n16367\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26066\,
            I => \c0.rx.n16368\
        );

    \I__4458\ : InMux
    port map (
            O => \N__26063\,
            I => \c0.rx.n16369\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26060\,
            I => \c0.rx.n16370\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26057\,
            I => \c0.rx.n16371\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__26054\,
            I => \c0.n18375_cascade_\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__26048\,
            I => \N__26045\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__26042\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__4450\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__26036\,
            I => \N__26032\
        );

    \I__4448\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26029\
        );

    \I__4447\ : Span4Mux_h
    port map (
            O => \N__26032\,
            I => \N__26026\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__26029\,
            I => data_out_frame2_18_3
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__26026\,
            I => data_out_frame2_18_3
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__26015\,
            I => \N__26012\
        );

    \I__4441\ : Span4Mux_h
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__26006\,
            I => \c0.data_out_frame2_19_3\
        );

    \I__4438\ : InMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26000\,
            I => \N__25996\
        );

    \I__4436\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25993\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__25996\,
            I => \N__25990\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__25993\,
            I => data_out_frame2_16_3
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__25990\,
            I => data_out_frame2_16_3
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__25985\,
            I => \c0.n18510_cascade_\
        );

    \I__4431\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25975\
        );

    \I__4429\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25972\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__25975\,
            I => \N__25969\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__25972\,
            I => data_out_frame2_17_3
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__25969\,
            I => data_out_frame2_17_3
        );

    \I__4425\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__25955\,
            I => \c0.data_out_frame2_20_3\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__25952\,
            I => \c0.n18513_cascade_\
        );

    \I__4420\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__25946\,
            I => \c0.n22_adj_2527\
        );

    \I__4418\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25939\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__25942\,
            I => \N__25936\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__25939\,
            I => \N__25932\
        );

    \I__4415\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25927\
        );

    \I__4414\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25927\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__25932\,
            I => \N__25923\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__25927\,
            I => \N__25920\
        );

    \I__4411\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25917\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__25923\,
            I => n9652
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__25920\,
            I => n9652
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__25917\,
            I => n9652
        );

    \I__4407\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25902\
        );

    \I__4405\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25897\
        );

    \I__4404\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25897\
        );

    \I__4403\ : Span4Mux_h
    port map (
            O => \N__25902\,
            I => \N__25892\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__25897\,
            I => \N__25892\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__25892\,
            I => n9922
        );

    \I__4400\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25885\
        );

    \I__4399\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25881\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__25885\,
            I => \N__25878\
        );

    \I__4397\ : InMux
    port map (
            O => \N__25884\,
            I => \N__25875\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25872\
        );

    \I__4395\ : Sp12to4
    port map (
            O => \N__25878\,
            I => \N__25866\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__25875\,
            I => \N__25866\
        );

    \I__4393\ : Span4Mux_s3_v
    port map (
            O => \N__25872\,
            I => \N__25863\
        );

    \I__4392\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25860\
        );

    \I__4391\ : Span12Mux_s3_v
    port map (
            O => \N__25866\,
            I => \N__25857\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__25863\,
            I => \N__25854\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__25860\,
            I => \r_Bit_Index_2_adj_2635\
        );

    \I__4388\ : Odrv12
    port map (
            O => \N__25857\,
            I => \r_Bit_Index_2_adj_2635\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__25854\,
            I => \r_Bit_Index_2_adj_2635\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__4385\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__25838\,
            I => \c0.n17559\
        );

    \I__4382\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25828\
        );

    \I__4380\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25825\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__25825\,
            I => \N__25819\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__25822\,
            I => \N__25816\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__25819\,
            I => n9135
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__25816\,
            I => n9135
        );

    \I__4374\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25807\
        );

    \I__4373\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25804\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__25804\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__25801\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__4369\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__25793\,
            I => \c0.n18082\
        );

    \I__4367\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25786\
        );

    \I__4366\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25783\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__25786\,
            I => \c0.n14631\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__25783\,
            I => \c0.n14631\
        );

    \I__4363\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25774\
        );

    \I__4362\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__25774\,
            I => data_out_frame2_12_3
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__25771\,
            I => data_out_frame2_12_3
        );

    \I__4359\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25760\
        );

    \I__4358\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25760\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__25760\,
            I => data_in_20_2
        );

    \I__4356\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__25754\,
            I => \c0.n17815\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__4353\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__25745\,
            I => \c0.n17818\
        );

    \I__4351\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__4349\ : Span4Mux_h
    port map (
            O => \N__25736\,
            I => \N__25733\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__25733\,
            I => \c0.n6_adj_2432\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__25730\,
            I => \c0.n18372_cascade_\
        );

    \I__4346\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__25724\,
            I => \N__25720\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25717\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__25720\,
            I => \N__25714\
        );

    \I__4342\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25711\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__25714\,
            I => \N__25705\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__25711\,
            I => \N__25705\
        );

    \I__4339\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25702\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__25702\,
            I => data_in_7_3
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__25699\,
            I => data_in_7_3
        );

    \I__4335\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__25691\,
            I => n18054
        );

    \I__4333\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25684\
        );

    \I__4332\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25681\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__25684\,
            I => \N__25678\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__25681\,
            I => \N__25673\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__25678\,
            I => \N__25673\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__25673\,
            I => data_out_frame2_10_4
        );

    \I__4327\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25666\
        );

    \I__4326\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__25666\,
            I => \N__25658\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25658\
        );

    \I__4323\ : Odrv12
    port map (
            O => \N__25658\,
            I => data_out_frame2_11_4
        );

    \I__4322\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__25652\,
            I => \N__25648\
        );

    \I__4320\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__4319\ : Span12Mux_v
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__25645\,
            I => data_out_frame2_14_5
        );

    \I__4317\ : Odrv12
    port map (
            O => \N__25642\,
            I => data_out_frame2_14_5
        );

    \I__4316\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25632\
        );

    \I__4315\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25628\
        );

    \I__4314\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25625\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25622\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__25631\,
            I => \N__25619\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__25628\,
            I => \N__25614\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__25625\,
            I => \N__25614\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__25622\,
            I => \N__25611\
        );

    \I__4308\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25608\
        );

    \I__4307\ : Span4Mux_v
    port map (
            O => \N__25614\,
            I => \N__25605\
        );

    \I__4306\ : Span4Mux_v
    port map (
            O => \N__25611\,
            I => \N__25600\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25600\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__25605\,
            I => \N__25597\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__25600\,
            I => \N__25594\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__25597\,
            I => \c0.data_in_frame_10_0\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__25594\,
            I => \c0.data_in_frame_10_0\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__25589\,
            I => \N__25584\
        );

    \I__4299\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25579\
        );

    \I__4298\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25576\
        );

    \I__4297\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25573\
        );

    \I__4296\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25570\
        );

    \I__4295\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25567\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__25579\,
            I => \N__25564\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__25576\,
            I => \N__25561\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__25573\,
            I => \N__25556\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__25570\,
            I => \N__25556\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__25567\,
            I => \N__25550\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__25564\,
            I => \N__25550\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__25561\,
            I => \N__25545\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__25556\,
            I => \N__25545\
        );

    \I__4286\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25542\
        );

    \I__4285\ : Span4Mux_v
    port map (
            O => \N__25550\,
            I => \N__25539\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__25545\,
            I => \N__25536\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__25542\,
            I => data_in_frame_8_3
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__25539\,
            I => data_in_frame_8_3
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__25536\,
            I => data_in_frame_8_3
        );

    \I__4280\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__25526\,
            I => \N__25522\
        );

    \I__4278\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25519\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__25522\,
            I => \N__25516\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25513\
        );

    \I__4275\ : Span4Mux_h
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__25513\,
            I => \N__25507\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__25510\,
            I => n9380
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__25507\,
            I => n9380
        );

    \I__4271\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25498\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25495\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25492\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25489\
        );

    \I__4267\ : Span4Mux_s3_h
    port map (
            O => \N__25492\,
            I => \N__25486\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__25486\,
            I => \N__25480\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__25483\,
            I => n9054
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__25480\,
            I => n9054
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__25475\,
            I => \n6_adj_2604_cascade_\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25468\
        );

    \I__4260\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25465\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25462\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__25465\,
            I => \N__25458\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__25462\,
            I => \N__25455\
        );

    \I__4256\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25452\
        );

    \I__4255\ : Odrv12
    port map (
            O => \N__25458\,
            I => data_in_frame_7_0
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__25455\,
            I => data_in_frame_7_0
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__25452\,
            I => data_in_frame_7_0
        );

    \I__4252\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25440\
        );

    \I__4251\ : InMux
    port map (
            O => \N__25444\,
            I => \N__25437\
        );

    \I__4250\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25434\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__25440\,
            I => \N__25429\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__25437\,
            I => \N__25424\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__25434\,
            I => \N__25424\
        );

    \I__4246\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25421\
        );

    \I__4245\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25418\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__25429\,
            I => \N__25413\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__25424\,
            I => \N__25413\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__25421\,
            I => \N__25410\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__25418\,
            I => \c0.data_in_frame_1_7\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__25413\,
            I => \c0.data_in_frame_1_7\
        );

    \I__4239\ : Odrv12
    port map (
            O => \N__25410\,
            I => \c0.data_in_frame_1_7\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__4237\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25396\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__25399\,
            I => \N__25393\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__25396\,
            I => \N__25390\
        );

    \I__4234\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25386\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__25390\,
            I => \N__25382\
        );

    \I__4232\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25379\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__25386\,
            I => \N__25376\
        );

    \I__4230\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25373\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__25382\,
            I => \N__25366\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__25379\,
            I => \N__25366\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__25376\,
            I => \N__25366\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__25373\,
            I => \c0.data_in_frame_3_5\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__25366\,
            I => \c0.data_in_frame_3_5\
        );

    \I__4224\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25358\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__4222\ : Span4Mux_v
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__25349\,
            I => \c0.n17614\
        );

    \I__4219\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25342\
        );

    \I__4218\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25339\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25336\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25333\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25326\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__25333\,
            I => \N__25326\
        );

    \I__4213\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25321\
        );

    \I__4212\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25321\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__25326\,
            I => \c0.n8666\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__25321\,
            I => \c0.n8666\
        );

    \I__4209\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__4207\ : Span4Mux_s1_h
    port map (
            O => \N__25310\,
            I => \N__25306\
        );

    \I__4206\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25303\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__25306\,
            I => \N__25300\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__25303\,
            I => data_out_frame2_14_1
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__25300\,
            I => data_out_frame2_14_1
        );

    \I__4202\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25292\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25292\,
            I => n18104
        );

    \I__4200\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25286\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__25286\,
            I => n18097
        );

    \I__4198\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__25280\,
            I => n18103
        );

    \I__4196\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__25274\,
            I => \N__25267\
        );

    \I__4194\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25264\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__25272\,
            I => \N__25260\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \N__25257\
        );

    \I__4191\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25254\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__25267\,
            I => \N__25251\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__25264\,
            I => \N__25248\
        );

    \I__4188\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25241\
        );

    \I__4187\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25241\
        );

    \I__4186\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25241\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__25254\,
            I => data_in_frame_5_4
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__25251\,
            I => data_in_frame_5_4
        );

    \I__4183\ : Odrv12
    port map (
            O => \N__25248\,
            I => data_in_frame_5_4
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__25241\,
            I => data_in_frame_5_4
        );

    \I__4181\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__4179\ : Span4Mux_h
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__25223\,
            I => \c0.n2603\
        );

    \I__4177\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__25211\,
            I => n2568
        );

    \I__4173\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25204\
        );

    \I__4172\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25201\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25198\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__25201\,
            I => \c0.n17538\
        );

    \I__4169\ : Odrv12
    port map (
            O => \N__25198\,
            I => \c0.n17538\
        );

    \I__4168\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25186\
        );

    \I__4166\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25183\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__25186\,
            I => \c0.n9355\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__25183\,
            I => \c0.n9355\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__25178\,
            I => \n2568_cascade_\
        );

    \I__4162\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25171\
        );

    \I__4161\ : InMux
    port map (
            O => \N__25174\,
            I => \N__25168\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__25171\,
            I => \N__25165\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25168\,
            I => \N__25162\
        );

    \I__4158\ : Span4Mux_h
    port map (
            O => \N__25165\,
            I => \N__25159\
        );

    \I__4157\ : Span4Mux_v
    port map (
            O => \N__25162\,
            I => \N__25156\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__25159\,
            I => \N__25153\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__25153\,
            I => \c0.n17541\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__25150\,
            I => \c0.n17541\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \c0.n21_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__25139\,
            I => \c0.n25\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__25136\,
            I => \c0.n27_cascade_\
        );

    \I__4148\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25129\
        );

    \I__4147\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25123\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__25126\,
            I => \N__25120\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__25120\,
            I => \c0.n5_adj_2438\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__25117\,
            I => \c0.n5_adj_2438\
        );

    \I__4141\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25103\
        );

    \I__4139\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25100\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__25107\,
            I => \N__25097\
        );

    \I__4137\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25094\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__25103\,
            I => \N__25089\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25089\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25086\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25094\,
            I => \N__25083\
        );

    \I__4132\ : Span4Mux_v
    port map (
            O => \N__25089\,
            I => \N__25080\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25086\,
            I => \c0.data_in_frame_6_7\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__25083\,
            I => \c0.data_in_frame_6_7\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__25080\,
            I => \c0.data_in_frame_6_7\
        );

    \I__4128\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__4126\ : Odrv12
    port map (
            O => \N__25067\,
            I => \c0.n4_adj_2548\
        );

    \I__4125\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25059\
        );

    \I__4124\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25056\
        );

    \I__4123\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25053\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__25049\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25046\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__25043\
        );

    \I__4119\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25040\
        );

    \I__4118\ : Span4Mux_v
    port map (
            O => \N__25049\,
            I => \N__25037\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__25046\,
            I => \N__25032\
        );

    \I__4116\ : Span4Mux_s3_h
    port map (
            O => \N__25043\,
            I => \N__25032\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__25040\,
            I => data_in_frame_8_4
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__25037\,
            I => data_in_frame_8_4
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__25032\,
            I => data_in_frame_8_4
        );

    \I__4112\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__25022\,
            I => \N__25018\
        );

    \I__4110\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25015\
        );

    \I__4109\ : Span4Mux_v
    port map (
            O => \N__25018\,
            I => \N__25012\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__25006\,
            I => \N__25000\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__25003\,
            I => n19_adj_2651
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__25000\,
            I => n19_adj_2651
        );

    \I__4102\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24991\
        );

    \I__4101\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24988\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24985\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__24988\,
            I => \N__24982\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__24985\,
            I => \N__24979\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__24982\,
            I => \N__24976\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__24979\,
            I => \c0.n8658\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__24976\,
            I => \c0.n8658\
        );

    \I__4094\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24967\
        );

    \I__4093\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24964\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__24967\,
            I => \N__24960\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24957\
        );

    \I__4090\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24952\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__24960\,
            I => \N__24947\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__24957\,
            I => \N__24947\
        );

    \I__4087\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24942\
        );

    \I__4086\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24942\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__24952\,
            I => data_in_frame_5_1
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__24947\,
            I => data_in_frame_5_1
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__24942\,
            I => data_in_frame_5_1
        );

    \I__4082\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24932\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24928\
        );

    \I__4080\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24925\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__24922\,
            I => \N__24916\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__24919\,
            I => \c0.n17516\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__24916\,
            I => \c0.n17516\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__24911\,
            I => \c0.n2601_cascade_\
        );

    \I__4073\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24905\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__24905\,
            I => \N__24902\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__24902\,
            I => \N__24897\
        );

    \I__4070\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24894\
        );

    \I__4069\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24891\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__24897\,
            I => n2597
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__24894\,
            I => n2597
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__24891\,
            I => n2597
        );

    \I__4065\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24880\
        );

    \I__4064\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24876\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__24880\,
            I => \N__24873\
        );

    \I__4062\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24870\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__24876\,
            I => \N__24867\
        );

    \I__4060\ : Span4Mux_s3_h
    port map (
            O => \N__24873\,
            I => \N__24864\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__24870\,
            I => \N__24861\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__24867\,
            I => \N__24856\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__24864\,
            I => \N__24856\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__24861\,
            I => \N__24853\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__24856\,
            I => \c0.n9039\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__24853\,
            I => \c0.n9039\
        );

    \I__4053\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__24839\,
            I => \N__24835\
        );

    \I__4049\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24832\
        );

    \I__4048\ : Span4Mux_s2_h
    port map (
            O => \N__24835\,
            I => \N__24829\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__24829\,
            I => \c0.n17522\
        );

    \I__4045\ : Odrv12
    port map (
            O => \N__24826\,
            I => \c0.n17522\
        );

    \I__4044\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__24818\,
            I => \c0.n2606\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \c0.n17428_cascade_\
        );

    \I__4041\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__24809\,
            I => \c0.n11_adj_2494\
        );

    \I__4039\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__4037\ : Span4Mux_v
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__4036\ : Span4Mux_s2_h
    port map (
            O => \N__24797\,
            I => \N__24794\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__24794\,
            I => \c0.n14\
        );

    \I__4034\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24785\
        );

    \I__4033\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24785\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__24785\,
            I => \c0.n17575\
        );

    \I__4031\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24778\
        );

    \I__4030\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24775\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__24778\,
            I => \N__24772\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__24775\,
            I => \N__24769\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__24772\,
            I => \c0.n9103\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__24769\,
            I => \c0.n9103\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__24764\,
            I => \N__24760\
        );

    \I__4024\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24755\
        );

    \I__4023\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24750\
        );

    \I__4022\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24747\
        );

    \I__4021\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24744\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24741\
        );

    \I__4019\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24736\
        );

    \I__4018\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24736\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__24750\,
            I => \N__24733\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24730\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__24744\,
            I => \N__24725\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__24741\,
            I => \N__24725\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24722\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__24733\,
            I => \N__24715\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__24730\,
            I => \N__24715\
        );

    \I__4010\ : Sp12to4
    port map (
            O => \N__24725\,
            I => \N__24710\
        );

    \I__4009\ : Span12Mux_s11_v
    port map (
            O => \N__24722\,
            I => \N__24710\
        );

    \I__4008\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24705\
        );

    \I__4007\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24705\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__24715\,
            I => data_in_frame_5_2
        );

    \I__4005\ : Odrv12
    port map (
            O => \N__24710\,
            I => data_in_frame_5_2
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__24705\,
            I => data_in_frame_5_2
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__4002\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24688\
        );

    \I__4001\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24683\
        );

    \I__4000\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24683\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__24692\,
            I => \N__24679\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__24691\,
            I => \N__24674\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24670\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__24683\,
            I => \N__24667\
        );

    \I__3995\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24660\
        );

    \I__3994\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24660\
        );

    \I__3993\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24660\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__24677\,
            I => \N__24657\
        );

    \I__3991\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24654\
        );

    \I__3990\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24651\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__24670\,
            I => \N__24648\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__24667\,
            I => \N__24643\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__24660\,
            I => \N__24643\
        );

    \I__3986\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24640\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24637\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24634\
        );

    \I__3983\ : Sp12to4
    port map (
            O => \N__24648\,
            I => \N__24631\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__24643\,
            I => \N__24628\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24621\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__24637\,
            I => \N__24621\
        );

    \I__3979\ : Span4Mux_s2_h
    port map (
            O => \N__24634\,
            I => \N__24621\
        );

    \I__3978\ : Odrv12
    port map (
            O => \N__24631\,
            I => data_in_frame_5_6
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__24628\,
            I => data_in_frame_5_6
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__24621\,
            I => data_in_frame_5_6
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__3974\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__24608\,
            I => \c0.n17430\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__3971\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24595\
        );

    \I__3969\ : InMux
    port map (
            O => \N__24598\,
            I => \N__24591\
        );

    \I__3968\ : Span12Mux_s4_h
    port map (
            O => \N__24595\,
            I => \N__24588\
        );

    \I__3967\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24585\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__24591\,
            I => data_in_7_0
        );

    \I__3965\ : Odrv12
    port map (
            O => \N__24588\,
            I => data_in_7_0
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__24585\,
            I => data_in_7_0
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__24578\,
            I => \c0.n4_adj_2512_cascade_\
        );

    \I__3962\ : InMux
    port map (
            O => \N__24575\,
            I => \N__24572\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__3960\ : Span4Mux_s3_h
    port map (
            O => \N__24569\,
            I => \N__24566\
        );

    \I__3959\ : Span4Mux_v
    port map (
            O => \N__24566\,
            I => \N__24563\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__24563\,
            I => n2591
        );

    \I__3957\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__24557\,
            I => \N__24552\
        );

    \I__3955\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24549\
        );

    \I__3954\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24546\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__24552\,
            I => \N__24543\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__24549\,
            I => \N__24540\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__24546\,
            I => \N__24537\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__24543\,
            I => \N__24532\
        );

    \I__3949\ : Span4Mux_s3_h
    port map (
            O => \N__24540\,
            I => \N__24532\
        );

    \I__3948\ : Span4Mux_h
    port map (
            O => \N__24537\,
            I => \N__24529\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__24532\,
            I => \c0.n8751\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__24529\,
            I => \c0.n8751\
        );

    \I__3945\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24520\
        );

    \I__3944\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24517\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__24520\,
            I => \N__24514\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24509\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__24514\,
            I => \N__24509\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__24509\,
            I => \c0.n17532\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__24506\,
            I => \n2591_cascade_\
        );

    \I__3938\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24496\
        );

    \I__3936\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24487\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__24490\,
            I => \c0.n9324\
        );

    \I__3932\ : Odrv12
    port map (
            O => \N__24487\,
            I => \c0.n9324\
        );

    \I__3931\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__24479\,
            I => \c0.n17533\
        );

    \I__3929\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__24473\,
            I => \c0.n2605\
        );

    \I__3927\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__24461\,
            I => n2570
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__24458\,
            I => \n2570_cascade_\
        );

    \I__3922\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__24449\,
            I => \c0.n8556\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__24446\,
            I => \c0.n17_adj_2514_cascade_\
        );

    \I__3918\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24440\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24435\
        );

    \I__3916\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24430\
        );

    \I__3915\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24430\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__24435\,
            I => \N__24427\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24424\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__24427\,
            I => \c0.data_in_frame_6_2\
        );

    \I__3911\ : Odrv12
    port map (
            O => \N__24424\,
            I => \c0.data_in_frame_6_2\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__24419\,
            I => \FRAME_MATCHER_next_state_31_N_2026_1_cascade_\
        );

    \I__3909\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24412\
        );

    \I__3908\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24409\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24406\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__24409\,
            I => \N__24403\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__24406\,
            I => \N__24400\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__24403\,
            I => n2567
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__24400\,
            I => n2567
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__24395\,
            I => \c0.n8556_cascade_\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__24392\,
            I => \c0.n7_cascade_\
        );

    \I__3900\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__24386\,
            I => \c0.n6_adj_2478\
        );

    \I__3898\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__3896\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24371\
        );

    \I__3895\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24367\
        );

    \I__3894\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24364\
        );

    \I__3893\ : Span4Mux_v
    port map (
            O => \N__24374\,
            I => \N__24361\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24358\
        );

    \I__3891\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24355\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24367\,
            I => data_in_2_2
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__24364\,
            I => data_in_2_2
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__24361\,
            I => data_in_2_2
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__24358\,
            I => data_in_2_2
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__24355\,
            I => data_in_2_2
        );

    \I__3885\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24340\
        );

    \I__3884\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24337\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__24340\,
            I => \c0.n8460\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__24337\,
            I => \c0.n8460\
        );

    \I__3881\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__3879\ : Odrv12
    port map (
            O => \N__24326\,
            I => \c0.n17745\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \c0.n16_adj_2485_cascade_\
        );

    \I__3877\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24310\
        );

    \I__3876\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24310\
        );

    \I__3875\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24307\
        );

    \I__3874\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24304\
        );

    \I__3873\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24299\
        );

    \I__3872\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24299\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__24310\,
            I => \N__24294\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__24307\,
            I => \N__24294\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__24304\,
            I => \N__24291\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__24299\,
            I => \N__24284\
        );

    \I__3867\ : Span4Mux_v
    port map (
            O => \N__24294\,
            I => \N__24284\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__24291\,
            I => \N__24284\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__24284\,
            I => data_in_frame_10_6
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \n63_adj_2642_cascade_\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__24278\,
            I => \N__24247\
        );

    \I__3862\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24230\
        );

    \I__3861\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24230\
        );

    \I__3860\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24230\
        );

    \I__3859\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24227\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24222\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24222\
        );

    \I__3856\ : InMux
    port map (
            O => \N__24271\,
            I => \N__24219\
        );

    \I__3855\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24205\
        );

    \I__3854\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24205\
        );

    \I__3853\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24205\
        );

    \I__3852\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24202\
        );

    \I__3851\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24193\
        );

    \I__3850\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24193\
        );

    \I__3849\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24193\
        );

    \I__3848\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24193\
        );

    \I__3847\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24184\
        );

    \I__3846\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24184\
        );

    \I__3845\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24184\
        );

    \I__3844\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24184\
        );

    \I__3843\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24181\
        );

    \I__3842\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24176\
        );

    \I__3841\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24176\
        );

    \I__3840\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24171\
        );

    \I__3839\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24171\
        );

    \I__3838\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24162\
        );

    \I__3837\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24162\
        );

    \I__3836\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24162\
        );

    \I__3835\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24162\
        );

    \I__3834\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24159\
        );

    \I__3833\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24152\
        );

    \I__3832\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24152\
        );

    \I__3831\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24152\
        );

    \I__3830\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24143\
        );

    \I__3829\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24143\
        );

    \I__3828\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24143\
        );

    \I__3827\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24143\
        );

    \I__3826\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24136\
        );

    \I__3825\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24136\
        );

    \I__3824\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24136\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24131\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__24227\,
            I => \N__24131\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__24222\,
            I => \N__24126\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__24219\,
            I => \N__24126\
        );

    \I__3819\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24122\
        );

    \I__3818\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24119\
        );

    \I__3817\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24115\
        );

    \I__3816\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24106\
        );

    \I__3815\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24106\
        );

    \I__3814\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24106\
        );

    \I__3813\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24106\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__24205\,
            I => \N__24103\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24096\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N__24096\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__24184\,
            I => \N__24096\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__24181\,
            I => \N__24091\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24091\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24171\,
            I => \N__24086\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24086\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24073\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24073\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__24143\,
            I => \N__24073\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__24136\,
            I => \N__24073\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__24131\,
            I => \N__24073\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__24126\,
            I => \N__24073\
        );

    \I__3798\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24066\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__24122\,
            I => \N__24061\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__24119\,
            I => \N__24061\
        );

    \I__3795\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24058\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24049\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__24106\,
            I => \N__24049\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__24103\,
            I => \N__24049\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__24096\,
            I => \N__24049\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__24091\,
            I => \N__24044\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24044\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__24073\,
            I => \N__24041\
        );

    \I__3787\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24032\
        );

    \I__3786\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24032\
        );

    \I__3785\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24032\
        );

    \I__3784\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24032\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__24066\,
            I => \N__24025\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__24061\,
            I => \N__24025\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24025\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__24049\,
            I => n16468
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__24044\,
            I => n16468
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__24041\,
            I => n16468
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__24032\,
            I => n16468
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__24025\,
            I => n16468
        );

    \I__3775\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__24008\,
            I => \N__24004\
        );

    \I__3772\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23999\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__24004\,
            I => \N__23996\
        );

    \I__3770\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23991\
        );

    \I__3769\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23991\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__23999\,
            I => \c0.data_in_1_0\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__23996\,
            I => \c0.data_in_1_0\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__23991\,
            I => \c0.data_in_1_0\
        );

    \I__3765\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23981\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__23978\,
            I => \N__23974\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__23977\,
            I => \N__23970\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__23974\,
            I => \N__23966\
        );

    \I__3760\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23959\
        );

    \I__3759\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23959\
        );

    \I__3758\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23959\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__23966\,
            I => \c0.data_in_0_0\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__23959\,
            I => \c0.data_in_0_0\
        );

    \I__3755\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3753\ : Span4Mux_v
    port map (
            O => \N__23948\,
            I => \N__23941\
        );

    \I__3752\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23938\
        );

    \I__3751\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23931\
        );

    \I__3750\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23931\
        );

    \I__3749\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23931\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__23941\,
            I => data_in_3_7
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__23938\,
            I => data_in_3_7
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__23931\,
            I => data_in_3_7
        );

    \I__3745\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__23921\,
            I => \c0.n6_adj_2473\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__3742\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3740\ : Span4Mux_v
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__23906\,
            I => \N__23902\
        );

    \I__3738\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23899\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__23902\,
            I => \N__23894\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23894\
        );

    \I__3735\ : Span4Mux_v
    port map (
            O => \N__23894\,
            I => \N__23890\
        );

    \I__3734\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23887\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__23890\,
            I => data_in_8_0
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__23887\,
            I => data_in_8_0
        );

    \I__3731\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23878\
        );

    \I__3730\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23874\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__23878\,
            I => \N__23870\
        );

    \I__3728\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23867\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23863\
        );

    \I__3726\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23860\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__23870\,
            I => \N__23856\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__23867\,
            I => \N__23853\
        );

    \I__3723\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23850\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__23863\,
            I => \N__23845\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23845\
        );

    \I__3720\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23842\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__23856\,
            I => \c0.n81\
        );

    \I__3718\ : Odrv12
    port map (
            O => \N__23853\,
            I => \c0.n81\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__23850\,
            I => \c0.n81\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__23845\,
            I => \c0.n81\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__23842\,
            I => \c0.n81\
        );

    \I__3714\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23827\
        );

    \I__3713\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23824\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23820\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23817\
        );

    \I__3710\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23814\
        );

    \I__3709\ : Span12Mux_h
    port map (
            O => \N__23820\,
            I => \N__23811\
        );

    \I__3708\ : Odrv12
    port map (
            O => \N__23817\,
            I => data_in_6_0
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__23814\,
            I => data_in_6_0
        );

    \I__3706\ : Odrv12
    port map (
            O => \N__23811\,
            I => data_in_6_0
        );

    \I__3705\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__3703\ : Span4Mux_v
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__3702\ : Span4Mux_h
    port map (
            O => \N__23795\,
            I => \N__23790\
        );

    \I__3701\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23787\
        );

    \I__3700\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23784\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__23790\,
            I => \c0.data_in_frame_6_0\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__23787\,
            I => \c0.data_in_frame_6_0\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__23784\,
            I => \c0.data_in_frame_6_0\
        );

    \I__3696\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23774\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__23774\,
            I => \N__23770\
        );

    \I__3694\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23767\
        );

    \I__3693\ : Span4Mux_h
    port map (
            O => \N__23770\,
            I => \N__23764\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__23767\,
            I => \N__23761\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__23764\,
            I => n2599
        );

    \I__3690\ : Odrv12
    port map (
            O => \N__23761\,
            I => n2599
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \n2599_cascade_\
        );

    \I__3688\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23747\
        );

    \I__3686\ : Span4Mux_h
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__23744\,
            I => \c0.n20_adj_2452\
        );

    \I__3684\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23733\
        );

    \I__3682\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23730\
        );

    \I__3681\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23727\
        );

    \I__3680\ : Odrv12
    port map (
            O => \N__23733\,
            I => data_in_0_2
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__23730\,
            I => data_in_0_2
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__23727\,
            I => data_in_0_2
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__23720\,
            I => \c0.n12_adj_2472_cascade_\
        );

    \I__3676\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__23708\,
            I => \c0.n17765\
        );

    \I__3672\ : InMux
    port map (
            O => \N__23705\,
            I => n16349
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__3670\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23695\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__23698\,
            I => \N__23692\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__23695\,
            I => \N__23689\
        );

    \I__3667\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23686\
        );

    \I__3666\ : Span4Mux_s2_h
    port map (
            O => \N__23689\,
            I => \N__23683\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__23686\,
            I => \N__23680\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__23683\,
            I => \N__23675\
        );

    \I__3663\ : Span4Mux_v
    port map (
            O => \N__23680\,
            I => \N__23672\
        );

    \I__3662\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23669\
        );

    \I__3661\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23666\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__23675\,
            I => \N__23663\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__23672\,
            I => data_in_5_3
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__23669\,
            I => data_in_5_3
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__23666\,
            I => data_in_5_3
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__23663\,
            I => data_in_5_3
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__23654\,
            I => \c0.n17715_cascade_\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__3653\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__3651\ : Span4Mux_h
    port map (
            O => \N__23642\,
            I => \N__23638\
        );

    \I__3650\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23635\
        );

    \I__3649\ : Span4Mux_v
    port map (
            O => \N__23638\,
            I => \N__23632\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__23635\,
            I => data_out_frame2_15_5
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__23632\,
            I => data_out_frame2_15_5
        );

    \I__3646\ : InMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3644\ : Span4Mux_h
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__23615\,
            I => \c0.n18540\
        );

    \I__3641\ : InMux
    port map (
            O => \N__23612\,
            I => n16340
        );

    \I__3640\ : InMux
    port map (
            O => \N__23609\,
            I => n16341
        );

    \I__3639\ : InMux
    port map (
            O => \N__23606\,
            I => \bfn_5_32_0_\
        );

    \I__3638\ : InMux
    port map (
            O => \N__23603\,
            I => n16343
        );

    \I__3637\ : InMux
    port map (
            O => \N__23600\,
            I => n16344
        );

    \I__3636\ : InMux
    port map (
            O => \N__23597\,
            I => n16345
        );

    \I__3635\ : InMux
    port map (
            O => \N__23594\,
            I => n16346
        );

    \I__3634\ : InMux
    port map (
            O => \N__23591\,
            I => n16347
        );

    \I__3633\ : InMux
    port map (
            O => \N__23588\,
            I => n16348
        );

    \I__3632\ : InMux
    port map (
            O => \N__23585\,
            I => n16330
        );

    \I__3631\ : InMux
    port map (
            O => \N__23582\,
            I => n16331
        );

    \I__3630\ : InMux
    port map (
            O => \N__23579\,
            I => n16332
        );

    \I__3629\ : InMux
    port map (
            O => \N__23576\,
            I => n16333
        );

    \I__3628\ : InMux
    port map (
            O => \N__23573\,
            I => \bfn_5_31_0_\
        );

    \I__3627\ : InMux
    port map (
            O => \N__23570\,
            I => n16335
        );

    \I__3626\ : InMux
    port map (
            O => \N__23567\,
            I => n16336
        );

    \I__3625\ : InMux
    port map (
            O => \N__23564\,
            I => n16337
        );

    \I__3624\ : InMux
    port map (
            O => \N__23561\,
            I => n16338
        );

    \I__3623\ : InMux
    port map (
            O => \N__23558\,
            I => n16339
        );

    \I__3622\ : InMux
    port map (
            O => \N__23555\,
            I => n16321
        );

    \I__3621\ : InMux
    port map (
            O => \N__23552\,
            I => n16322
        );

    \I__3620\ : InMux
    port map (
            O => \N__23549\,
            I => n16323
        );

    \I__3619\ : InMux
    port map (
            O => \N__23546\,
            I => n16324
        );

    \I__3618\ : InMux
    port map (
            O => \N__23543\,
            I => n16325
        );

    \I__3617\ : InMux
    port map (
            O => \N__23540\,
            I => \bfn_5_30_0_\
        );

    \I__3616\ : InMux
    port map (
            O => \N__23537\,
            I => n16327
        );

    \I__3615\ : InMux
    port map (
            O => \N__23534\,
            I => n16328
        );

    \I__3614\ : InMux
    port map (
            O => \N__23531\,
            I => n16329
        );

    \I__3613\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23524\
        );

    \I__3612\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__23524\,
            I => \N__23516\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__23521\,
            I => \N__23516\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__23513\,
            I => \c0.n17482\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__23510\,
            I => \N__23506\
        );

    \I__3606\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__3605\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23500\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23497\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__23500\,
            I => data_out_frame2_9_3
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__23497\,
            I => data_out_frame2_9_3
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__23492\,
            I => \N__23488\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__23491\,
            I => \N__23485\
        );

    \I__3599\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23480\
        );

    \I__3598\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23480\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__23480\,
            I => data_out_frame2_8_3
        );

    \I__3596\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3594\ : Odrv12
    port map (
            O => \N__23471\,
            I => \c0.n18522\
        );

    \I__3593\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23461\
        );

    \I__3591\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23458\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__23461\,
            I => \N__23455\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__23458\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__23455\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3586\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__3584\ : Sp12to4
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__3583\ : Odrv12
    port map (
            O => \N__23438\,
            I => \c0.n18076\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__3581\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23428\
        );

    \I__3580\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23425\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__23428\,
            I => data_out_frame2_9_7
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__23425\,
            I => data_out_frame2_9_7
        );

    \I__3577\ : CascadeMux
    port map (
            O => \N__23420\,
            I => \N__23416\
        );

    \I__3576\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23413\
        );

    \I__3575\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23410\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__23413\,
            I => data_out_frame2_8_7
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__23410\,
            I => data_out_frame2_8_7
        );

    \I__3572\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__23399\,
            I => \c0.n18588\
        );

    \I__3569\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__23390\,
            I => \c0.n17785\
        );

    \I__3566\ : InMux
    port map (
            O => \N__23387\,
            I => \bfn_5_29_0_\
        );

    \I__3565\ : InMux
    port map (
            O => \N__23384\,
            I => n16319
        );

    \I__3564\ : InMux
    port map (
            O => \N__23381\,
            I => n16320
        );

    \I__3563\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23374\
        );

    \I__3562\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23371\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__23374\,
            I => \N__23368\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__23371\,
            I => data_out_frame2_9_6
        );

    \I__3559\ : Odrv12
    port map (
            O => \N__23368\,
            I => data_out_frame2_9_6
        );

    \I__3558\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23359\
        );

    \I__3557\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23356\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__23359\,
            I => data_out_frame2_15_3
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__23356\,
            I => data_out_frame2_15_3
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23347\
        );

    \I__3553\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23344\
        );

    \I__3552\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23341\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__23344\,
            I => data_out_frame2_14_3
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__23341\,
            I => data_out_frame2_14_3
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__23336\,
            I => \c0.n18516_cascade_\
        );

    \I__3548\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23326\
        );

    \I__3546\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23323\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__23326\,
            I => \N__23320\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__23323\,
            I => data_out_frame2_13_3
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__23320\,
            I => data_out_frame2_13_3
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3541\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23308\
        );

    \I__3540\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23305\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__23308\,
            I => data_out_frame2_11_1
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__23305\,
            I => data_out_frame2_11_1
        );

    \I__3537\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23296\
        );

    \I__3536\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__23296\,
            I => data_out_frame2_10_1
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__23293\,
            I => data_out_frame2_10_1
        );

    \I__3533\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__3531\ : Span4Mux_h
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__23279\,
            I => \c0.n18480\
        );

    \I__3529\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23273\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__23273\,
            I => \c0.n136\
        );

    \I__3527\ : InMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23264\
        );

    \I__3525\ : Span4Mux_v
    port map (
            O => \N__23264\,
            I => \N__23260\
        );

    \I__3524\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23257\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__23260\,
            I => \c0.n1_adj_2443\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__23257\,
            I => \c0.n1_adj_2443\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__23252\,
            I => \c0.n14631_cascade_\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__3519\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23239\
        );

    \I__3517\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__3516\ : Span4Mux_h
    port map (
            O => \N__23239\,
            I => \N__23233\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__23236\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__23233\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__3513\ : InMux
    port map (
            O => \N__23228\,
            I => \c0.tx.n16358\
        );

    \I__3512\ : InMux
    port map (
            O => \N__23225\,
            I => \c0.tx.n16359\
        );

    \I__3511\ : InMux
    port map (
            O => \N__23222\,
            I => \c0.tx.n16360\
        );

    \I__3510\ : InMux
    port map (
            O => \N__23219\,
            I => \c0.tx.n16361\
        );

    \I__3509\ : InMux
    port map (
            O => \N__23216\,
            I => \c0.tx.n16362\
        );

    \I__3508\ : InMux
    port map (
            O => \N__23213\,
            I => \c0.tx.n16363\
        );

    \I__3507\ : InMux
    port map (
            O => \N__23210\,
            I => \bfn_5_26_0_\
        );

    \I__3506\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23203\
        );

    \I__3505\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23200\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__23203\,
            I => \N__23195\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__23200\,
            I => \N__23192\
        );

    \I__3502\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23187\
        );

    \I__3501\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23187\
        );

    \I__3500\ : Span4Mux_v
    port map (
            O => \N__23195\,
            I => \N__23184\
        );

    \I__3499\ : Span4Mux_v
    port map (
            O => \N__23192\,
            I => \N__23181\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__23187\,
            I => \c0.n31\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__23184\,
            I => \c0.n31\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__23181\,
            I => \c0.n31\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__23174\,
            I => \c0.n17582_cascade_\
        );

    \I__3494\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__3492\ : Span4Mux_h
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__3491\ : Span4Mux_v
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__23159\,
            I => \c0.data_out_frame2_20_7\
        );

    \I__3489\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__3487\ : Span4Mux_h
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__23147\,
            I => n2560
        );

    \I__3485\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__23138\,
            I => \c0.n17588\
        );

    \I__3482\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__23132\,
            I => \c0.n17582\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \n2560_cascade_\
        );

    \I__3479\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23122\
        );

    \I__3478\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23119\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__23119\,
            I => \N__23113\
        );

    \I__3475\ : Odrv12
    port map (
            O => \N__23116\,
            I => n17585
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__23113\,
            I => n17585
        );

    \I__3473\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__23105\,
            I => \c0.n17648\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__23102\,
            I => \c0.n18_cascade_\
        );

    \I__3470\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23095\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23092\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__23095\,
            I => \c0.n17418\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__23092\,
            I => \c0.n17418\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23084\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23080\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23077\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__23080\,
            I => n2572
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23077\,
            I => n2572
        );

    \I__3461\ : InMux
    port map (
            O => \N__23072\,
            I => \bfn_5_25_0_\
        );

    \I__3460\ : InMux
    port map (
            O => \N__23069\,
            I => \c0.tx.n16357\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23062\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23059\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__23056\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__23059\,
            I => \c0.n8695\
        );

    \I__3455\ : Odrv12
    port map (
            O => \N__23056\,
            I => \c0.n8695\
        );

    \I__3454\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23047\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23044\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23040\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23037\
        );

    \I__3450\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23034\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__23040\,
            I => \N__23029\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__23037\,
            I => \N__23029\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__23034\,
            I => \c0.data_in_frame_6_6\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__23029\,
            I => \c0.data_in_frame_6_6\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23019\
        );

    \I__3444\ : InMux
    port map (
            O => \N__23023\,
            I => \N__23016\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23013\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__23019\,
            I => \N__23010\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__23007\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__23013\,
            I => \N__23004\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__23010\,
            I => \N__23001\
        );

    \I__3438\ : Span4Mux_v
    port map (
            O => \N__23007\,
            I => \N__22998\
        );

    \I__3437\ : Odrv12
    port map (
            O => \N__23004\,
            I => \c0.n9208\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__23001\,
            I => \c0.n9208\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__22998\,
            I => \c0.n9208\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__22991\,
            I => \c0.n22_cascade_\
        );

    \I__3433\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__22985\,
            I => n16_adj_2656
        );

    \I__3431\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__22979\,
            I => \c0.n17519\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \c0.n24_cascade_\
        );

    \I__3428\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__22967\,
            I => \N__22964\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__22964\,
            I => \c0.n11_adj_2453\
        );

    \I__3424\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22957\
        );

    \I__3423\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22954\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22949\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__22954\,
            I => \N__22946\
        );

    \I__3420\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22943\
        );

    \I__3419\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22940\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__22949\,
            I => \N__22935\
        );

    \I__3417\ : Span4Mux_s2_h
    port map (
            O => \N__22946\,
            I => \N__22935\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__22943\,
            I => data_in_frame_8_2
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__22940\,
            I => data_in_frame_8_2
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__22935\,
            I => data_in_frame_8_2
        );

    \I__3413\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22922\
        );

    \I__3412\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22917\
        );

    \I__3411\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22917\
        );

    \I__3410\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22914\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N__22909\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22909\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__22914\,
            I => data_in_frame_8_1
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__22909\,
            I => data_in_frame_8_1
        );

    \I__3405\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22897\
        );

    \I__3404\ : InMux
    port map (
            O => \N__22903\,
            I => \N__22897\
        );

    \I__3403\ : InMux
    port map (
            O => \N__22902\,
            I => \N__22894\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22890\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22887\
        );

    \I__3400\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22884\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__22890\,
            I => \N__22881\
        );

    \I__3398\ : Span4Mux_h
    port map (
            O => \N__22887\,
            I => \N__22876\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22876\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__22881\,
            I => \c0.data_in_frame_6_3\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__22876\,
            I => \c0.data_in_frame_6_3\
        );

    \I__3394\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22865\
        );

    \I__3393\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22865\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__22865\,
            I => \c0.n17605\
        );

    \I__3391\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__22859\,
            I => \c0.n20\
        );

    \I__3389\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__22847\,
            I => \N__22843\
        );

    \I__3385\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22840\
        );

    \I__3384\ : Span4Mux_s1_h
    port map (
            O => \N__22843\,
            I => \N__22836\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__22840\,
            I => \N__22833\
        );

    \I__3382\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22828\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__22836\,
            I => \N__22823\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__22833\,
            I => \N__22823\
        );

    \I__3379\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22820\
        );

    \I__3378\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22817\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22814\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__22823\,
            I => \c0.data_in_frame_7_6\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__22820\,
            I => \c0.data_in_frame_7_6\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__22817\,
            I => \c0.data_in_frame_7_6\
        );

    \I__3373\ : Odrv12
    port map (
            O => \N__22814\,
            I => \c0.data_in_frame_7_6\
        );

    \I__3372\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22798\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22795\
        );

    \I__3369\ : Span4Mux_v
    port map (
            O => \N__22798\,
            I => \N__22792\
        );

    \I__3368\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__22792\,
            I => \c0.n9144\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__22789\,
            I => \c0.n9144\
        );

    \I__3365\ : InMux
    port map (
            O => \N__22784\,
            I => \N__22780\
        );

    \I__3364\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22777\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22774\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__22777\,
            I => \c0.n8064\
        );

    \I__3361\ : Odrv12
    port map (
            O => \N__22774\,
            I => \c0.n8064\
        );

    \I__3360\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22762\
        );

    \I__3359\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22762\
        );

    \I__3358\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22759\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22756\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__22759\,
            I => \N__22752\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__22756\,
            I => \N__22749\
        );

    \I__3354\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22746\
        );

    \I__3353\ : Span4Mux_v
    port map (
            O => \N__22752\,
            I => \N__22739\
        );

    \I__3352\ : Span4Mux_h
    port map (
            O => \N__22749\,
            I => \N__22739\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22739\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__22739\,
            I => \c0.n8687\
        );

    \I__3349\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__22730\,
            I => \N__22726\
        );

    \I__3346\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22723\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__22726\,
            I => n2585
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__22723\,
            I => n2585
        );

    \I__3343\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__22715\,
            I => \c0.n17\
        );

    \I__3341\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__22709\,
            I => n2590
        );

    \I__3339\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22702\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__22705\,
            I => \N__22699\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22696\
        );

    \I__3336\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22692\
        );

    \I__3335\ : Span4Mux_h
    port map (
            O => \N__22696\,
            I => \N__22689\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__22695\,
            I => \N__22686\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22683\
        );

    \I__3332\ : Span4Mux_h
    port map (
            O => \N__22689\,
            I => \N__22680\
        );

    \I__3331\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22677\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__22683\,
            I => \c0.data_in_frame_7_1\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__22680\,
            I => \c0.data_in_frame_7_1\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__22677\,
            I => \c0.data_in_frame_7_1\
        );

    \I__3327\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22665\
        );

    \I__3326\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22662\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__22668\,
            I => \N__22659\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__22665\,
            I => \N__22654\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__22662\,
            I => \N__22654\
        );

    \I__3322\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22650\
        );

    \I__3321\ : Span4Mux_s3_h
    port map (
            O => \N__22654\,
            I => \N__22647\
        );

    \I__3320\ : InMux
    port map (
            O => \N__22653\,
            I => \N__22644\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__22650\,
            I => \c0.data_in_frame_1_0\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__22647\,
            I => \c0.data_in_frame_1_0\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__22644\,
            I => \c0.data_in_frame_1_0\
        );

    \I__3316\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22632\
        );

    \I__3315\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22629\
        );

    \I__3314\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22624\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__22632\,
            I => \N__22621\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__22629\,
            I => \N__22618\
        );

    \I__3311\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22615\
        );

    \I__3310\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22612\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22609\
        );

    \I__3308\ : Span4Mux_s2_h
    port map (
            O => \N__22621\,
            I => \N__22604\
        );

    \I__3307\ : Span4Mux_h
    port map (
            O => \N__22618\,
            I => \N__22604\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__22615\,
            I => \c0.data_in_frame_4_6\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__22612\,
            I => \c0.data_in_frame_4_6\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__22609\,
            I => \c0.data_in_frame_4_6\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__22604\,
            I => \c0.data_in_frame_4_6\
        );

    \I__3302\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__22592\,
            I => \N__22587\
        );

    \I__3300\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22584\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__22590\,
            I => \N__22581\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__22587\,
            I => \N__22577\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22574\
        );

    \I__3296\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22571\
        );

    \I__3295\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22568\
        );

    \I__3294\ : Span4Mux_v
    port map (
            O => \N__22577\,
            I => \N__22563\
        );

    \I__3293\ : Span4Mux_v
    port map (
            O => \N__22574\,
            I => \N__22563\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22560\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__22568\,
            I => \c0.data_in_frame_3_0\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__22563\,
            I => \c0.data_in_frame_3_0\
        );

    \I__3289\ : Odrv12
    port map (
            O => \N__22560\,
            I => \c0.data_in_frame_3_0\
        );

    \I__3288\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22549\
        );

    \I__3287\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22545\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22539\
        );

    \I__3285\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22536\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22533\
        );

    \I__3283\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22530\
        );

    \I__3282\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22525\
        );

    \I__3281\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22525\
        );

    \I__3280\ : Span4Mux_v
    port map (
            O => \N__22539\,
            I => \N__22518\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__22536\,
            I => \N__22518\
        );

    \I__3278\ : Span4Mux_v
    port map (
            O => \N__22533\,
            I => \N__22518\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__22530\,
            I => \c0.data_in_frame_4_7\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__22525\,
            I => \c0.data_in_frame_4_7\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__22518\,
            I => \c0.data_in_frame_4_7\
        );

    \I__3274\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__22502\,
            I => \c0.n17403\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__22499\,
            I => \c0.n17403_cascade_\
        );

    \I__3269\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22489\
        );

    \I__3267\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22486\
        );

    \I__3266\ : Span4Mux_v
    port map (
            O => \N__22489\,
            I => \N__22481\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22477\
        );

    \I__3264\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22474\
        );

    \I__3263\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22471\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__22481\,
            I => \N__22468\
        );

    \I__3261\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22465\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__22477\,
            I => \N__22460\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22460\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__22471\,
            I => \c0.data_in_frame_2_6\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__22468\,
            I => \c0.data_in_frame_2_6\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__22465\,
            I => \c0.data_in_frame_2_6\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__22460\,
            I => \c0.data_in_frame_2_6\
        );

    \I__3254\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22447\
        );

    \I__3253\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22444\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22441\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22438\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__22441\,
            I => \N__22433\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__22438\,
            I => \N__22433\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__22433\,
            I => n9283
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__22430\,
            I => \n9283_cascade_\
        );

    \I__3246\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__22424\,
            I => \N__22421\
        );

    \I__3244\ : Sp12to4
    port map (
            O => \N__22421\,
            I => \N__22417\
        );

    \I__3243\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22414\
        );

    \I__3242\ : Span12Mux_s7_v
    port map (
            O => \N__22417\,
            I => \N__22411\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__22414\,
            I => data_out_frame2_16_7
        );

    \I__3240\ : Odrv12
    port map (
            O => \N__22411\,
            I => data_out_frame2_16_7
        );

    \I__3239\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22402\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__22405\,
            I => \N__22399\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__22402\,
            I => \N__22396\
        );

    \I__3236\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22393\
        );

    \I__3235\ : Span4Mux_v
    port map (
            O => \N__22396\,
            I => \N__22390\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22387\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__22390\,
            I => \N__22382\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__22387\,
            I => \N__22382\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__22382\,
            I => \c0.n9219\
        );

    \I__3230\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22372\
        );

    \I__3228\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22369\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__22372\,
            I => \N__22366\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__22369\,
            I => n2593
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__22366\,
            I => n2593
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__22361\,
            I => \n2593_cascade_\
        );

    \I__3223\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__22355\,
            I => \c0.n22_adj_2461\
        );

    \I__3221\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__22346\,
            I => \N__22342\
        );

    \I__3218\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22339\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__22342\,
            I => n2586
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__22339\,
            I => n2586
        );

    \I__3215\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22330\
        );

    \I__3214\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22327\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22324\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22321\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__22324\,
            I => \N__22316\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__22321\,
            I => \N__22316\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__22316\,
            I => \c0.n9279\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \n2590_cascade_\
        );

    \I__3207\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__22307\,
            I => \c0.n10_adj_2450\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__3204\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22293\
        );

    \I__3202\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22288\
        );

    \I__3201\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22288\
        );

    \I__3200\ : Span4Mux_v
    port map (
            O => \N__22293\,
            I => \N__22285\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__22288\,
            I => data_in_6_3
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__22285\,
            I => data_in_6_3
        );

    \I__3197\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__22274\,
            I => \N__22270\
        );

    \I__3194\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22267\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__22270\,
            I => n2596
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__22267\,
            I => n2596
        );

    \I__3191\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22258\
        );

    \I__3190\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22255\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22250\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__22255\,
            I => \N__22250\
        );

    \I__3187\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__22247\,
            I => \c0.n17529\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__22244\,
            I => \n2596_cascade_\
        );

    \I__3184\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__22232\,
            I => \c0.n10_adj_2498\
        );

    \I__3180\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22221\
        );

    \I__3178\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22218\
        );

    \I__3177\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22215\
        );

    \I__3176\ : Span4Mux_s3_h
    port map (
            O => \N__22221\,
            I => \N__22212\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22209\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__22215\,
            I => \c0.data_in_frame_7_3\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__22212\,
            I => \c0.data_in_frame_7_3\
        );

    \I__3172\ : Odrv12
    port map (
            O => \N__22209\,
            I => \c0.data_in_frame_7_3\
        );

    \I__3171\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22196\
        );

    \I__3170\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22196\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__22196\,
            I => n2588
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__22193\,
            I => \c0.n8695_cascade_\
        );

    \I__3167\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22180\
        );

    \I__3164\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22177\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__22180\,
            I => \c0.n8867\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__22177\,
            I => \c0.n8867\
        );

    \I__3161\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22165\
        );

    \I__3159\ : InMux
    port map (
            O => \N__22168\,
            I => \N__22162\
        );

    \I__3158\ : Span4Mux_v
    port map (
            O => \N__22165\,
            I => \N__22156\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__22162\,
            I => \N__22156\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22152\
        );

    \I__3155\ : Span4Mux_v
    port map (
            O => \N__22156\,
            I => \N__22149\
        );

    \I__3154\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22146\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__22152\,
            I => \c0.data_in_frame_0_6\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__22149\,
            I => \c0.data_in_frame_0_6\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__22146\,
            I => \c0.data_in_frame_0_6\
        );

    \I__3150\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22135\
        );

    \I__3149\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22130\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__22135\,
            I => \N__22127\
        );

    \I__3147\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22124\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \N__22121\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22114\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__22127\,
            I => \N__22114\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__22124\,
            I => \N__22114\
        );

    \I__3142\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22111\
        );

    \I__3141\ : Span4Mux_h
    port map (
            O => \N__22114\,
            I => \N__22108\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__22111\,
            I => \c0.data_in_frame_3_4\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__22108\,
            I => \c0.data_in_frame_3_4\
        );

    \I__3138\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22099\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__22102\,
            I => \N__22095\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22092\
        );

    \I__3135\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22087\
        );

    \I__3134\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22087\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__22092\,
            I => \N__22083\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__22087\,
            I => \N__22080\
        );

    \I__3131\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22077\
        );

    \I__3130\ : Sp12to4
    port map (
            O => \N__22083\,
            I => \N__22074\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__22080\,
            I => \N__22071\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22077\,
            I => data_in_5_0
        );

    \I__3127\ : Odrv12
    port map (
            O => \N__22074\,
            I => data_in_5_0
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__22071\,
            I => data_in_5_0
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__22064\,
            I => \N__22060\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__22063\,
            I => \N__22056\
        );

    \I__3123\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22049\
        );

    \I__3122\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22049\
        );

    \I__3121\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22049\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__22049\,
            I => data_in_7_6
        );

    \I__3119\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__22043\,
            I => \N__22038\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \N__22035\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__22041\,
            I => \N__22030\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__22038\,
            I => \N__22027\
        );

    \I__3114\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22022\
        );

    \I__3113\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22022\
        );

    \I__3112\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22017\
        );

    \I__3111\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22017\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__22027\,
            I => \c0.data_in_frame_1_2\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__22022\,
            I => \c0.data_in_frame_1_2\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__22017\,
            I => \c0.data_in_frame_1_2\
        );

    \I__3107\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22006\
        );

    \I__3106\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22003\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__21999\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21996\
        );

    \I__3103\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21993\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__21999\,
            I => \N__21990\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__21996\,
            I => \N__21985\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__21993\,
            I => \N__21985\
        );

    \I__3099\ : Span4Mux_h
    port map (
            O => \N__21990\,
            I => \N__21982\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__21985\,
            I => \c0.data_in_frame_6_1\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__21982\,
            I => \c0.data_in_frame_6_1\
        );

    \I__3096\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21973\
        );

    \I__3095\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21970\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21967\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__3092\ : Span4Mux_h
    port map (
            O => \N__21967\,
            I => \N__21961\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__21964\,
            I => \N__21958\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__21961\,
            I => \c0.n9328\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__21958\,
            I => \c0.n9328\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__3087\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21943\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__21946\,
            I => \N__21940\
        );

    \I__3084\ : Span4Mux_v
    port map (
            O => \N__21943\,
            I => \N__21937\
        );

    \I__3083\ : InMux
    port map (
            O => \N__21940\,
            I => \N__21934\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__21937\,
            I => \c0.n8645\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__21934\,
            I => \c0.n8645\
        );

    \I__3080\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21925\
        );

    \I__3079\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21922\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__21925\,
            I => \N__21919\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__3076\ : Span12Mux_s4_h
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__21916\,
            I => n9100
        );

    \I__3074\ : Odrv12
    port map (
            O => \N__21913\,
            I => n9100
        );

    \I__3073\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21902\
        );

    \I__3072\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21899\
        );

    \I__3071\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21896\
        );

    \I__3070\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21892\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__21902\,
            I => \N__21885\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21885\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21885\
        );

    \I__3066\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21882\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__21892\,
            I => \N__21877\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__21885\,
            I => \N__21877\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21874\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__21877\,
            I => \c0.data_in_frame_4_5\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__21874\,
            I => \c0.data_in_frame_4_5\
        );

    \I__3060\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21865\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__21868\,
            I => \N__21862\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21859\
        );

    \I__3057\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21854\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__21859\,
            I => \N__21851\
        );

    \I__3055\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21846\
        );

    \I__3054\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21846\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__21854\,
            I => \c0.data_in_frame_0_5\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__21851\,
            I => \c0.data_in_frame_0_5\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__21846\,
            I => \c0.data_in_frame_0_5\
        );

    \I__3050\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21834\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__21838\,
            I => \N__21830\
        );

    \I__3048\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21826\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__21834\,
            I => \N__21823\
        );

    \I__3046\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21820\
        );

    \I__3045\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21817\
        );

    \I__3044\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21814\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__21826\,
            I => \N__21811\
        );

    \I__3042\ : Span4Mux_s2_h
    port map (
            O => \N__21823\,
            I => \N__21808\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__21820\,
            I => \N__21805\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21802\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21795\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__21811\,
            I => \N__21795\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__21808\,
            I => \N__21795\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__21805\,
            I => \N__21790\
        );

    \I__3035\ : Span4Mux_h
    port map (
            O => \N__21802\,
            I => \N__21790\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__21795\,
            I => \c0.data_in_frame_4_4\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__21790\,
            I => \c0.data_in_frame_4_4\
        );

    \I__3032\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__3030\ : Span4Mux_h
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__21776\,
            I => \c0.n9176\
        );

    \I__3028\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21769\
        );

    \I__3027\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21765\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21761\
        );

    \I__3025\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21758\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__21765\,
            I => \N__21755\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__21764\,
            I => \N__21751\
        );

    \I__3022\ : Span4Mux_s3_h
    port map (
            O => \N__21761\,
            I => \N__21748\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21745\
        );

    \I__3020\ : Span4Mux_s2_h
    port map (
            O => \N__21755\,
            I => \N__21742\
        );

    \I__3019\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21737\
        );

    \I__3018\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21737\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__21748\,
            I => \c0.data_in_frame_4_2\
        );

    \I__3016\ : Odrv12
    port map (
            O => \N__21745\,
            I => \c0.data_in_frame_4_2\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__21742\,
            I => \c0.data_in_frame_4_2\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__21737\,
            I => \c0.data_in_frame_4_2\
        );

    \I__3013\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21724\
        );

    \I__3012\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21719\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__21724\,
            I => \N__21715\
        );

    \I__3010\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21712\
        );

    \I__3009\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21709\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21706\
        );

    \I__3007\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21703\
        );

    \I__3006\ : Span4Mux_s1_h
    port map (
            O => \N__21715\,
            I => \N__21700\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__21712\,
            I => \c0.data_in_frame_2_3\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__21709\,
            I => \c0.data_in_frame_2_3\
        );

    \I__3003\ : Odrv12
    port map (
            O => \N__21706\,
            I => \c0.data_in_frame_2_3\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__21703\,
            I => \c0.data_in_frame_2_3\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__21700\,
            I => \c0.data_in_frame_2_3\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \c0.n10_adj_2430_cascade_\
        );

    \I__2999\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21680\
        );

    \I__2998\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21677\
        );

    \I__2997\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21674\
        );

    \I__2996\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21671\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__21680\,
            I => \N__21668\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21665\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__21674\,
            I => \N__21662\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__21671\,
            I => \c0.data_in_frame_4_1\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__21668\,
            I => \c0.data_in_frame_4_1\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__21665\,
            I => \c0.data_in_frame_4_1\
        );

    \I__2989\ : Odrv12
    port map (
            O => \N__21662\,
            I => \c0.data_in_frame_4_1\
        );

    \I__2988\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__21647\,
            I => \N__21642\
        );

    \I__2985\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21637\
        );

    \I__2984\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21637\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__21642\,
            I => data_in_0_7
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__21637\,
            I => data_in_0_7
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__21632\,
            I => \c0.n17697_cascade_\
        );

    \I__2980\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21625\
        );

    \I__2979\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21621\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__21625\,
            I => \N__21618\
        );

    \I__2977\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21615\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__21621\,
            I => data_in_0_4
        );

    \I__2975\ : Odrv12
    port map (
            O => \N__21618\,
            I => data_in_0_4
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__21615\,
            I => data_in_0_4
        );

    \I__2973\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__2972\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21599\
        );

    \I__2971\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21596\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__21605\,
            I => \N__21593\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21589\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21584\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__21596\,
            I => \N__21584\
        );

    \I__2966\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21579\
        );

    \I__2965\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21576\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__21589\,
            I => \N__21573\
        );

    \I__2963\ : Span4Mux_h
    port map (
            O => \N__21584\,
            I => \N__21570\
        );

    \I__2962\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21565\
        );

    \I__2961\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21565\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__21579\,
            I => data_in_frame_5_0
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__21576\,
            I => data_in_frame_5_0
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__21573\,
            I => data_in_frame_5_0
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__21570\,
            I => data_in_frame_5_0
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__21565\,
            I => data_in_frame_5_0
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__21554\,
            I => \N__21549\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21546\
        );

    \I__2953\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21543\
        );

    \I__2952\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21540\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__21546\,
            I => \c0.n9306\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__21543\,
            I => \c0.n9306\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__21540\,
            I => \c0.n9306\
        );

    \I__2948\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__21530\,
            I => \c0.tx2.n4\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__21527\,
            I => \c0.tx2.n9568_cascade_\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21520\
        );

    \I__2944\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__21520\,
            I => \c0.tx2.tx2_active\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__21517\,
            I => \c0.tx2.tx2_active\
        );

    \I__2941\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21509\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__21509\,
            I => \c0.tx2.n23\
        );

    \I__2939\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21502\
        );

    \I__2938\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21497\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21494\
        );

    \I__2936\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21491\
        );

    \I__2935\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21488\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__21497\,
            I => \c0.r_SM_Main_2_N_2326_0\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__21494\,
            I => \c0.r_SM_Main_2_N_2326_0\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__21491\,
            I => \c0.r_SM_Main_2_N_2326_0\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__21488\,
            I => \c0.r_SM_Main_2_N_2326_0\
        );

    \I__2930\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__21473\,
            I => \c0.tx2.n17990\
        );

    \I__2927\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21462\
        );

    \I__2926\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21455\
        );

    \I__2925\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21455\
        );

    \I__2924\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21455\
        );

    \I__2923\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21452\
        );

    \I__2922\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21449\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21444\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21444\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21452\,
            I => \c0.tx2.r_SM_Main_2_N_2323_1\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__21449\,
            I => \c0.tx2.r_SM_Main_2_N_2323_1\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__21444\,
            I => \c0.tx2.r_SM_Main_2_N_2323_1\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__21437\,
            I => \c0.tx2.n12_cascade_\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__21434\,
            I => \N__21427\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__21433\,
            I => \N__21422\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__21432\,
            I => \N__21418\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21406\
        );

    \I__2911\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21401\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21401\
        );

    \I__2909\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21398\
        );

    \I__2908\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21391\
        );

    \I__2907\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21391\
        );

    \I__2906\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21391\
        );

    \I__2905\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21382\
        );

    \I__2904\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21382\
        );

    \I__2903\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21382\
        );

    \I__2902\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21382\
        );

    \I__2901\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21379\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21368\
        );

    \I__2899\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21368\
        );

    \I__2898\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21368\
        );

    \I__2897\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21368\
        );

    \I__2896\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21368\
        );

    \I__2895\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21365\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__21401\,
            I => \N__21360\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21360\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__21391\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__21382\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__21379\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__21368\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__21365\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__21360\,
            I => \r_SM_Main_2_adj_2628\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21337\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21330\
        );

    \I__2883\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21330\
        );

    \I__2882\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21330\
        );

    \I__2881\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21327\
        );

    \I__2880\ : Span4Mux_s3_h
    port map (
            O => \N__21337\,
            I => \N__21320\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__21330\,
            I => \N__21315\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__21327\,
            I => \N__21315\
        );

    \I__2877\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21312\
        );

    \I__2876\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21305\
        );

    \I__2875\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21305\
        );

    \I__2874\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21305\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__21320\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__2872\ : Odrv12
    port map (
            O => \N__21315\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__21312\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__21305\,
            I => \c0.tx2.r_SM_Main_0\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__21296\,
            I => \N__21289\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \N__21285\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__21294\,
            I => \N__21280\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21276\
        );

    \I__2865\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21267\
        );

    \I__2864\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21267\
        );

    \I__2863\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21267\
        );

    \I__2862\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21267\
        );

    \I__2861\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21261\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21261\
        );

    \I__2859\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21258\
        );

    \I__2858\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21255\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__21276\,
            I => \N__21250\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21250\
        );

    \I__2855\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21247\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__21261\,
            I => \c0.tx2.r_SM_Main_1\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__21258\,
            I => \c0.tx2.r_SM_Main_1\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__21255\,
            I => \c0.tx2.r_SM_Main_1\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__21250\,
            I => \c0.tx2.r_SM_Main_1\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__21247\,
            I => \c0.tx2.r_SM_Main_1\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__21236\,
            I => \c0.tx2.n6812_cascade_\
        );

    \I__2848\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21229\
        );

    \I__2847\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__21229\,
            I => data_out_frame2_18_7
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__21226\,
            I => data_out_frame2_18_7
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__2843\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__2841\ : Odrv12
    port map (
            O => \N__21212\,
            I => \c0.data_out_frame2_19_7\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \c0.n18576_cascade_\
        );

    \I__2839\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21202\
        );

    \I__2838\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21199\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21196\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__21199\,
            I => data_out_frame2_17_7
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__21196\,
            I => data_out_frame2_17_7
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__21191\,
            I => \c0.n18579_cascade_\
        );

    \I__2833\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__21185\,
            I => \c0.n22_adj_2520\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__2830\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21176\,
            I => \c0.n17788\
        );

    \I__2828\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__21170\,
            I => \c0.n18420\
        );

    \I__2826\ : SRMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__21164\,
            I => \c0.n4_adj_2480\
        );

    \I__2824\ : IoInMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__2822\ : Odrv12
    port map (
            O => \N__21155\,
            I => tx_enable
        );

    \I__2821\ : IoInMux
    port map (
            O => \N__21152\,
            I => \N__21149\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__21149\,
            I => \N__21145\
        );

    \I__2819\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21142\
        );

    \I__2818\ : Span4Mux_s0_h
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21136\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__21139\,
            I => \N__21130\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__21136\,
            I => \N__21130\
        );

    \I__2814\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21127\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__21130\,
            I => tx2_o
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__21127\,
            I => tx2_o
        );

    \I__2811\ : IoInMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__2809\ : IoSpan4Mux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2808\ : Span4Mux_s3_h
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__2807\ : Span4Mux_h
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__21107\,
            I => tx2_enable
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__21104\,
            I => \c0.n17535_cascade_\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2803\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__2801\ : Span4Mux_s3_h
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__21089\,
            I => \c0.data_out_frame2_19_6\
        );

    \I__2799\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__21080\,
            I => \c0.n9240\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__21077\,
            I => \c0.n9240_cascade_\
        );

    \I__2795\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21068\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21068\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__2792\ : Span4Mux_v
    port map (
            O => \N__21065\,
            I => \N__21061\
        );

    \I__2791\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21058\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__21061\,
            I => \c0.n9131\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__21058\,
            I => \c0.n9131\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__21053\,
            I => \c0.n17409_cascade_\
        );

    \I__2787\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__21047\,
            I => \c0.n10_adj_2470\
        );

    \I__2785\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__2783\ : Span4Mux_s3_v
    port map (
            O => \N__21038\,
            I => \N__21035\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__21035\,
            I => \c0.data_out_frame2_20_1\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__2780\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__21023\,
            I => \c0.data_out_frame2_19_1\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__2775\ : Span4Mux_h
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__21011\,
            I => \c0.n6_adj_2464\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__21008\,
            I => \c0.n18423_cascade_\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__20999\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__2769\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20992\
        );

    \I__2768\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20989\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__20992\,
            I => \N__20986\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__20989\,
            I => data_out_frame2_15_4
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__20986\,
            I => data_out_frame2_15_4
        );

    \I__2764\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20977\
        );

    \I__2763\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20974\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__20977\,
            I => \N__20971\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__20974\,
            I => data_out_frame2_12_4
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__20971\,
            I => data_out_frame2_12_4
        );

    \I__2759\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20963\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__2757\ : Span4Mux_v
    port map (
            O => \N__20960\,
            I => \N__20956\
        );

    \I__2756\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20953\
        );

    \I__2755\ : Span4Mux_h
    port map (
            O => \N__20956\,
            I => \N__20950\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__20953\,
            I => data_out_frame2_13_6
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__20950\,
            I => data_out_frame2_13_6
        );

    \I__2752\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__20939\,
            I => \N__20935\
        );

    \I__2749\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20932\
        );

    \I__2748\ : Span4Mux_s1_h
    port map (
            O => \N__20935\,
            I => \N__20929\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__20932\,
            I => data_out_frame2_8_0
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__20929\,
            I => data_out_frame2_8_0
        );

    \I__2745\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20920\
        );

    \I__2744\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__20920\,
            I => data_out_frame2_10_7
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__20917\,
            I => data_out_frame2_10_7
        );

    \I__2741\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__20909\,
            I => \c0.n17647\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__20906\,
            I => \N__20902\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__20905\,
            I => \N__20899\
        );

    \I__2737\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20894\
        );

    \I__2736\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20894\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__20894\,
            I => \c0.n8995\
        );

    \I__2734\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__2732\ : Span4Mux_h
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__20882\,
            I => \c0.n6_adj_2550\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__2729\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__2727\ : Span12Mux_s3_h
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__20867\,
            I => \c0.data_out_frame2_20_0\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__20864\,
            I => \c0.n6_adj_2502_cascade_\
        );

    \I__2724\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__2722\ : Span4Mux_s3_h
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__20852\,
            I => \c0.data_out_frame2_20_2\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__2719\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__2717\ : Span4Mux_s1_h
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__20837\,
            I => \c0.data_out_frame2_19_5\
        );

    \I__2715\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__20831\,
            I => \N__20827\
        );

    \I__2713\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20824\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__20827\,
            I => \N__20821\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__20824\,
            I => data_out_frame2_14_0
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__20821\,
            I => data_out_frame2_14_0
        );

    \I__2709\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20809\
        );

    \I__2707\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20806\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__20809\,
            I => \N__20803\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__20806\,
            I => data_out_frame2_18_2
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__20803\,
            I => data_out_frame2_18_2
        );

    \I__2703\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__20792\,
            I => \N__20788\
        );

    \I__2700\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20785\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__20788\,
            I => \N__20782\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__20785\,
            I => data_out_frame2_5_6
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__20782\,
            I => data_out_frame2_5_6
        );

    \I__2696\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20770\
        );

    \I__2694\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__2693\ : Span4Mux_s3_v
    port map (
            O => \N__20770\,
            I => \N__20764\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__20767\,
            I => data_out_frame2_6_3
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__20764\,
            I => data_out_frame2_6_3
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2689\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__20753\,
            I => \N__20749\
        );

    \I__2687\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20746\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__20746\,
            I => data_out_frame2_12_6
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__20743\,
            I => data_out_frame2_12_6
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__20738\,
            I => \c0.n17647_cascade_\
        );

    \I__2682\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__20732\,
            I => \c0.n12_adj_2549\
        );

    \I__2680\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20725\
        );

    \I__2679\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20722\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20719\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20716\
        );

    \I__2676\ : Sp12to4
    port map (
            O => \N__20719\,
            I => \N__20713\
        );

    \I__2675\ : Span4Mux_s3_h
    port map (
            O => \N__20716\,
            I => \N__20709\
        );

    \I__2674\ : Span12Mux_v
    port map (
            O => \N__20713\,
            I => \N__20706\
        );

    \I__2673\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20703\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__20709\,
            I => data_in_8_5
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__20706\,
            I => data_in_8_5
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__20703\,
            I => data_in_8_5
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__2668\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__20690\,
            I => \N__20686\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__20689\,
            I => \N__20683\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__20686\,
            I => \N__20680\
        );

    \I__2664\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20677\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__20680\,
            I => \N__20674\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__20677\,
            I => \c0.n17602\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__20674\,
            I => \c0.n17602\
        );

    \I__2660\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20665\
        );

    \I__2659\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20662\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20659\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20656\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__20659\,
            I => \N__20653\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__20656\,
            I => \c0.n30_adj_2489\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__20653\,
            I => \c0.n30_adj_2489\
        );

    \I__2653\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__20645\,
            I => \c0.n9345\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__20642\,
            I => \c0.n9345_cascade_\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__20639\,
            I => \c0.n10_cascade_\
        );

    \I__2649\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__2647\ : Span4Mux_s3_v
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__20624\,
            I => \c0.data_out_frame2_20_6\
        );

    \I__2644\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__20618\,
            I => \N__20615\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__20612\,
            I => \N__20608\
        );

    \I__2640\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20605\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__20608\,
            I => \c0.n9163\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__20605\,
            I => \c0.n9163\
        );

    \I__2637\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20596\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__20599\,
            I => \N__20593\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__20596\,
            I => \N__20590\
        );

    \I__2634\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__2633\ : Span4Mux_s3_h
    port map (
            O => \N__20590\,
            I => \N__20584\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__20587\,
            I => \c0.n17470\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__20584\,
            I => \c0.n17470\
        );

    \I__2630\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20576\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__20576\,
            I => n9148
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__20573\,
            I => \n9148_cascade_\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__2626\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20563\
        );

    \I__2625\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20560\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20557\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20553\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__20557\,
            I => \N__20550\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20547\
        );

    \I__2620\ : Span12Mux_h
    port map (
            O => \N__20553\,
            I => \N__20544\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__20550\,
            I => \c0.n22_adj_2508\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__20547\,
            I => \c0.n22_adj_2508\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__20544\,
            I => \c0.n22_adj_2508\
        );

    \I__2616\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__2614\ : Odrv12
    port map (
            O => \N__20531\,
            I => \c0.n12_adj_2542\
        );

    \I__2613\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20524\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20520\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__20524\,
            I => \N__20517\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__20523\,
            I => \N__20514\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__20520\,
            I => \N__20510\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__20517\,
            I => \N__20507\
        );

    \I__2607\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20502\
        );

    \I__2606\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20502\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__20510\,
            I => \N__20499\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__20507\,
            I => \c0.data_in_frame_2_2\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__20502\,
            I => \c0.data_in_frame_2_2\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__20499\,
            I => \c0.data_in_frame_2_2\
        );

    \I__2601\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20486\
        );

    \I__2600\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20486\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__20483\,
            I => \N__20478\
        );

    \I__2597\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20475\
        );

    \I__2596\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20472\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__20478\,
            I => \N__20467\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20467\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__20472\,
            I => \c0.n9058\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__20467\,
            I => \c0.n9058\
        );

    \I__2591\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20458\
        );

    \I__2590\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20455\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__20452\,
            I => \N__20446\
        );

    \I__2586\ : Odrv12
    port map (
            O => \N__20449\,
            I => \c0.n17467\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__20446\,
            I => \c0.n17467\
        );

    \I__2584\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__20438\,
            I => \N__20434\
        );

    \I__2582\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20431\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__20434\,
            I => \N__20428\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__20431\,
            I => \N__20419\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__20428\,
            I => \N__20419\
        );

    \I__2578\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20414\
        );

    \I__2577\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20414\
        );

    \I__2576\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20409\
        );

    \I__2575\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20409\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__20419\,
            I => \c0.data_in_frame_4_3\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__20414\,
            I => \c0.data_in_frame_4_3\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__20409\,
            I => \c0.data_in_frame_4_3\
        );

    \I__2571\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20398\
        );

    \I__2570\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20395\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20392\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__20395\,
            I => \N__20389\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__20392\,
            I => \N__20386\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__20389\,
            I => \c0.n17562\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__20386\,
            I => \c0.n17562\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__20381\,
            I => \N__20377\
        );

    \I__2563\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20372\
        );

    \I__2562\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20369\
        );

    \I__2561\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20366\
        );

    \I__2560\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20363\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__20372\,
            I => \N__20360\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__20369\,
            I => \N__20355\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20355\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20350\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__20360\,
            I => \N__20350\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__20355\,
            I => data_in_frame_8_7
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__20350\,
            I => data_in_frame_8_7
        );

    \I__2552\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__20342\,
            I => \N__20338\
        );

    \I__2550\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20335\
        );

    \I__2549\ : Span4Mux_h
    port map (
            O => \N__20338\,
            I => \N__20332\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__20335\,
            I => data_out_frame2_6_7
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__20332\,
            I => data_out_frame2_6_7
        );

    \I__2546\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__20315\,
            I => \c0.n5_adj_2501\
        );

    \I__2541\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__20309\,
            I => \c0.n17534\
        );

    \I__2539\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20302\
        );

    \I__2538\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20299\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20296\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20291\
        );

    \I__2535\ : Span4Mux_s3_h
    port map (
            O => \N__20296\,
            I => \N__20291\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__20291\,
            I => \N__20286\
        );

    \I__2533\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20281\
        );

    \I__2532\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20281\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__20286\,
            I => \c0.n8674\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__20281\,
            I => \c0.n8674\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20270\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \N__20267\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20262\
        );

    \I__2526\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20254\
        );

    \I__2525\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20254\
        );

    \I__2524\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20254\
        );

    \I__2523\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20247\
        );

    \I__2522\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20247\
        );

    \I__2521\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20247\
        );

    \I__2520\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20244\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__20254\,
            I => n9419
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__20247\,
            I => n9419
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__20244\,
            I => n9419
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__2515\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__20228\,
            I => \c0.n8061\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__2511\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__2508\ : Span4Mux_s1_h
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__20210\,
            I => \c0.n8857\
        );

    \I__2506\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__20204\,
            I => \c0.n18_adj_2468\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__20201\,
            I => \c0.n26_adj_2469_cascade_\
        );

    \I__2503\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__20192\,
            I => \c0.n30\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__20189\,
            I => \c0.n12_adj_2449_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20179\
        );

    \I__2497\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20175\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__20179\,
            I => \N__20172\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20169\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__20175\,
            I => \N__20166\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__20172\,
            I => n2598
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__20169\,
            I => n2598
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__20166\,
            I => n2598
        );

    \I__2490\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__20150\,
            I => \c0.n23_adj_2462\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__20147\,
            I => \c0.n24_adj_2454_cascade_\
        );

    \I__2485\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20140\
        );

    \I__2484\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20137\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__20140\,
            I => \N__20132\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20129\
        );

    \I__2481\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20126\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \N__20123\
        );

    \I__2479\ : Span4Mux_s3_h
    port map (
            O => \N__20132\,
            I => \N__20115\
        );

    \I__2478\ : Span4Mux_s3_h
    port map (
            O => \N__20129\,
            I => \N__20115\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__20126\,
            I => \N__20115\
        );

    \I__2476\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20112\
        );

    \I__2475\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20109\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__20115\,
            I => \N__20104\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__20112\,
            I => \N__20104\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__20109\,
            I => data_in_frame_5_3
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__20104\,
            I => data_in_frame_5_3
        );

    \I__2470\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20095\
        );

    \I__2469\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20090\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__20095\,
            I => \N__20087\
        );

    \I__2467\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20082\
        );

    \I__2466\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20082\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20090\,
            I => \c0.data_in_frame_2_7\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__20087\,
            I => \c0.data_in_frame_2_7\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__20082\,
            I => \c0.data_in_frame_2_7\
        );

    \I__2462\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20068\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__20074\,
            I => \N__20065\
        );

    \I__2460\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20062\
        );

    \I__2459\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20057\
        );

    \I__2458\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20057\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20054\
        );

    \I__2456\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20051\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__20062\,
            I => \N__20048\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20045\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__20054\,
            I => \N__20036\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20036\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__20048\,
            I => \N__20036\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__20045\,
            I => \N__20036\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__20036\,
            I => \c0.data_in_frame_7_7\
        );

    \I__2448\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__2446\ : Span4Mux_s3_h
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__20024\,
            I => n2584
        );

    \I__2444\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__2442\ : Span4Mux_h
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__20009\,
            I => \c0.n9151\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__20006\,
            I => \n2584_cascade_\
        );

    \I__2438\ : InMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__20000\,
            I => \c0.n21_adj_2465\
        );

    \I__2436\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19993\
        );

    \I__2435\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__19993\,
            I => \N__19987\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__2432\ : Span4Mux_s3_h
    port map (
            O => \N__19987\,
            I => \N__19981\
        );

    \I__2431\ : Span4Mux_s3_h
    port map (
            O => \N__19984\,
            I => \N__19978\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__19981\,
            I => \N__19975\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__19975\,
            I => \c0.n8874\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__19972\,
            I => \c0.n8874\
        );

    \I__2426\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19960\
        );

    \I__2424\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19955\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__19960\,
            I => \N__19952\
        );

    \I__2422\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19947\
        );

    \I__2421\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19947\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__19955\,
            I => \c0.data_in_frame_1_4\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__19952\,
            I => \c0.data_in_frame_1_4\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__19947\,
            I => \c0.data_in_frame_1_4\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \c0.n8874_cascade_\
        );

    \I__2416\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19933\
        );

    \I__2415\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19930\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__19933\,
            I => \c0.n9349\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__19930\,
            I => \c0.n9349\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__19925\,
            I => \c0.n9368_cascade_\
        );

    \I__2411\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19915\
        );

    \I__2409\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19912\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__19912\,
            I => \c0.n23_adj_2426\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__19909\,
            I => \c0.n23_adj_2426\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19899\
        );

    \I__2404\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19893\
        );

    \I__2403\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19893\
        );

    \I__2402\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19888\
        );

    \I__2401\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19888\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19885\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__19888\,
            I => \c0.data_in_frame_1_6\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__19885\,
            I => \c0.data_in_frame_1_6\
        );

    \I__2397\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__19874\,
            I => \c0.n17632\
        );

    \I__2394\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__2392\ : Span4Mux_s3_h
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__19862\,
            I => \c0.n17485\
        );

    \I__2390\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19855\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__19858\,
            I => \N__19852\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__19855\,
            I => \N__19848\
        );

    \I__2387\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19845\
        );

    \I__2386\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19842\
        );

    \I__2385\ : Span4Mux_s3_h
    port map (
            O => \N__19848\,
            I => \N__19839\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__19845\,
            I => \c0.data_in_frame_3_1\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__19842\,
            I => \c0.data_in_frame_3_1\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__19839\,
            I => \c0.data_in_frame_3_1\
        );

    \I__2381\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__2379\ : Odrv12
    port map (
            O => \N__19826\,
            I => \c0.n17406\
        );

    \I__2378\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19817\
        );

    \I__2377\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19817\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__19817\,
            I => \c0.n13530\
        );

    \I__2375\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__19808\,
            I => \N__19804\
        );

    \I__2372\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19801\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__19804\,
            I => \c0.n17656\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__19801\,
            I => \c0.n17656\
        );

    \I__2369\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__19790\,
            I => \c0.n20_adj_2427\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \c0.n10_adj_2428_cascade_\
        );

    \I__2365\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__19778\,
            I => \c0.n17442\
        );

    \I__2362\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__19769\,
            I => \c0.n17553\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__19766\,
            I => \c0.n17442_cascade_\
        );

    \I__2358\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__19757\,
            I => \c0.n17550\
        );

    \I__2355\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19750\
        );

    \I__2354\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19745\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19742\
        );

    \I__2352\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19737\
        );

    \I__2351\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19737\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__19745\,
            I => \c0.data_in_frame_4_0\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__19742\,
            I => \c0.data_in_frame_4_0\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__19737\,
            I => \c0.data_in_frame_4_0\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19726\
        );

    \I__2346\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19721\
        );

    \I__2345\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19721\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__19721\,
            I => data_out_frame2_5_3
        );

    \I__2343\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19714\
        );

    \I__2342\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19711\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__19714\,
            I => \N__19708\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__19711\,
            I => data_out_frame2_7_3
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__19708\,
            I => data_out_frame2_7_3
        );

    \I__2338\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__19700\,
            I => \c0.n5_adj_2509\
        );

    \I__2336\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__2334\ : Span4Mux_s2_v
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__19688\,
            I => \N__19684\
        );

    \I__2332\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19681\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__19684\,
            I => \N__19678\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__19681\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__19678\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__2328\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__2326\ : Span4Mux_s2_v
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__2325\ : Span4Mux_v
    port map (
            O => \N__19664\,
            I => \N__19660\
        );

    \I__2324\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19657\
        );

    \I__2323\ : Span4Mux_v
    port map (
            O => \N__19660\,
            I => \N__19654\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__19657\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__19654\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__19649\,
            I => \c0.n18_adj_2544_cascade_\
        );

    \I__2319\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__2317\ : Span4Mux_s2_v
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__19637\,
            I => \N__19633\
        );

    \I__2315\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19630\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__19633\,
            I => \N__19627\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__19630\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__19627\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__19622\,
            I => \c0.n19_adj_2540_cascade_\
        );

    \I__2310\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__2308\ : Span12Mux_s2_h
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__2307\ : Odrv12
    port map (
            O => \N__19610\,
            I => \c0.tx2_transmit_N_2287\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__19607\,
            I => \c0.tx2_transmit_N_2287_cascade_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__19598\,
            I => \c0.n19_adj_2540\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__19595\,
            I => \c0.n67_cascade_\
        );

    \I__2301\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__2299\ : Span4Mux_s3_v
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__19583\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__2297\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__19574\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__19571\,
            I => \c0.tx2.n18612_cascade_\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__19565\,
            I => \c0.tx2.n18615\
        );

    \I__2291\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__19559\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__2289\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19552\
        );

    \I__2288\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19549\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__19552\,
            I => data_out_frame2_17_6
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__19549\,
            I => data_out_frame2_17_6
        );

    \I__2285\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19537\
        );

    \I__2283\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__2282\ : Span12Mux_s8_v
    port map (
            O => \N__19537\,
            I => \N__19531\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__19534\,
            I => data_out_frame2_13_4
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__19531\,
            I => data_out_frame2_13_4
        );

    \I__2279\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__19517\,
            I => \c0.n12\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \c0.n11_cascade_\
        );

    \I__2274\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__19499\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__2269\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__19493\,
            I => \c0.tx2.n18450\
        );

    \I__2267\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__19487\,
            I => \c0.tx2.n18453\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__2264\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__19475\,
            I => \N__19471\
        );

    \I__2261\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__2260\ : Span4Mux_s3_v
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__19468\,
            I => data_out_frame2_19_0
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__19465\,
            I => data_out_frame2_19_0
        );

    \I__2257\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__19457\,
            I => \c0.n18603\
        );

    \I__2255\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__19448\,
            I => \c0.n22_adj_2510\
        );

    \I__2252\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19441\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__19438\,
            I => data_out_frame2_14_7
        );

    \I__2248\ : Odrv12
    port map (
            O => \N__19435\,
            I => data_out_frame2_14_7
        );

    \I__2247\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19426\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__19423\,
            I => data_out_frame2_15_7
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__19420\,
            I => data_out_frame2_15_7
        );

    \I__2242\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19409\
        );

    \I__2241\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19409\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__19409\,
            I => data_out_frame2_12_7
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__19406\,
            I => \c0.n18582_cascade_\
        );

    \I__2238\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19399\
        );

    \I__2237\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19396\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__19396\,
            I => data_out_frame2_13_7
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__19393\,
            I => data_out_frame2_13_7
        );

    \I__2233\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19384\
        );

    \I__2232\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__19384\,
            I => data_out_frame2_9_2
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__19381\,
            I => data_out_frame2_9_2
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__2228\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19369\
        );

    \I__2227\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19366\,
            I => data_out_frame2_8_2
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__19363\,
            I => data_out_frame2_8_2
        );

    \I__2223\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__19355\,
            I => \c0.n18504\
        );

    \I__2221\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__2219\ : Span4Mux_s2_h
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__19343\,
            I => \c0.n17824\
        );

    \I__2217\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__19331\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__2212\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19321\
        );

    \I__2211\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__19318\,
            I => data_out_frame2_6_0
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__19315\,
            I => data_out_frame2_6_0
        );

    \I__2207\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19306\
        );

    \I__2206\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19303\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__19303\,
            I => data_out_frame2_7_1
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__19300\,
            I => data_out_frame2_7_1
        );

    \I__2202\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19288\
        );

    \I__2200\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19285\
        );

    \I__2199\ : Span4Mux_s2_h
    port map (
            O => \N__19288\,
            I => \N__19282\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__19285\,
            I => data_out_frame2_16_6
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__19282\,
            I => data_out_frame2_16_6
        );

    \I__2196\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19271\
        );

    \I__2195\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19271\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__19271\,
            I => data_out_frame2_11_7
        );

    \I__2193\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19264\
        );

    \I__2192\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19261\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__19264\,
            I => \N__19258\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__19261\,
            I => data_out_frame2_9_1
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__19258\,
            I => data_out_frame2_9_1
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__19253\,
            I => \N__19249\
        );

    \I__2187\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19244\
        );

    \I__2186\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19244\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__19244\,
            I => data_out_frame2_8_1
        );

    \I__2184\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__2182\ : Span4Mux_s2_h
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__19232\,
            I => \c0.n17833\
        );

    \I__2180\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19225\
        );

    \I__2179\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19222\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19219\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__2176\ : Span4Mux_s3_h
    port map (
            O => \N__19219\,
            I => \N__19213\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__19216\,
            I => data_out_frame2_6_1
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__19213\,
            I => data_out_frame2_6_1
        );

    \I__2173\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19204\
        );

    \I__2172\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19201\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19198\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__19201\,
            I => data_out_frame2_17_2
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__19198\,
            I => data_out_frame2_17_2
        );

    \I__2168\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19189\
        );

    \I__2167\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19186\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__19189\,
            I => data_out_frame2_5_7
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__19186\,
            I => data_out_frame2_5_7
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__2163\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19171\
        );

    \I__2161\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__19171\,
            I => \N__19165\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__19168\,
            I => data_out_frame2_6_5
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__19165\,
            I => data_out_frame2_6_5
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__2156\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__19154\,
            I => \N__19150\
        );

    \I__2154\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19147\
        );

    \I__2153\ : Span4Mux_s2_h
    port map (
            O => \N__19150\,
            I => \N__19144\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__19147\,
            I => data_out_frame2_12_1
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__19144\,
            I => data_out_frame2_12_1
        );

    \I__2150\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19132\
        );

    \I__2148\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19129\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__19132\,
            I => \N__19126\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__19129\,
            I => data_out_frame2_7_0
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__19126\,
            I => data_out_frame2_7_0
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__19121\,
            I => \n9606_cascade_\
        );

    \I__2143\ : InMux
    port map (
            O => \N__19118\,
            I => \N__19114\
        );

    \I__2142\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19111\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19108\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19103\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__19108\,
            I => \N__19103\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__19103\,
            I => data_out_frame2_10_5
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__2136\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19093\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19090\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19087\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__19090\,
            I => data_out_frame2_13_5
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__19087\,
            I => data_out_frame2_13_5
        );

    \I__2131\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__19079\,
            I => \N__19075\
        );

    \I__2129\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19072\
        );

    \I__2128\ : Span4Mux_s2_h
    port map (
            O => \N__19075\,
            I => \N__19069\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__19072\,
            I => data_out_frame2_9_0
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__19069\,
            I => data_out_frame2_9_0
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__19064\,
            I => \c0.n9151_cascade_\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__19061\,
            I => \c0.n17588_cascade_\
        );

    \I__2123\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19054\
        );

    \I__2122\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19050\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__19054\,
            I => \N__19047\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19044\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19050\,
            I => \N__19041\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__19047\,
            I => \N__19038\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19044\,
            I => data_in_frame_8_5
        );

    \I__2116\ : Odrv12
    port map (
            O => \N__19041\,
            I => data_in_frame_8_5
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__19038\,
            I => data_in_frame_8_5
        );

    \I__2114\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19028\,
            I => \c0.n6_adj_2429\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__2110\ : Span4Mux_s2_h
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__19016\,
            I => \c0.data_out_frame2_20_5\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__19013\,
            I => \N__19009\
        );

    \I__2107\ : InMux
    port map (
            O => \N__19012\,
            I => \N__19006\
        );

    \I__2106\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19003\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__19006\,
            I => data_out_frame2_12_2
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__19003\,
            I => data_out_frame2_12_2
        );

    \I__2103\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18991\
        );

    \I__2101\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__2100\ : Span4Mux_s2_h
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__18988\,
            I => data_out_frame2_13_1
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__18985\,
            I => data_out_frame2_13_1
        );

    \I__2097\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__18968\,
            I => \c0.n17424\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__2091\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__18956\,
            I => \c0.n17569\
        );

    \I__2088\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__18950\,
            I => \c0.n10_adj_2505\
        );

    \I__2086\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__18944\,
            I => \c0.n9028\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \c0.n8061_cascade_\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \N__18933\
        );

    \I__2082\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18930\
        );

    \I__2081\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18927\
        );

    \I__2080\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18924\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__18930\,
            I => \N__18919\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__18927\,
            I => \N__18919\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18916\
        );

    \I__2076\ : Span4Mux_s3_h
    port map (
            O => \N__18919\,
            I => \N__18911\
        );

    \I__2075\ : Span4Mux_s3_h
    port map (
            O => \N__18916\,
            I => \N__18911\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__18911\,
            I => \c0.data_in_frame_6_4\
        );

    \I__2073\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18904\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__18907\,
            I => \N__18900\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__18904\,
            I => \N__18897\
        );

    \I__2070\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18894\
        );

    \I__2069\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18891\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__18897\,
            I => n2595
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__18894\,
            I => n2595
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__18891\,
            I => n2595
        );

    \I__2065\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18880\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__18883\,
            I => \N__18877\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18873\
        );

    \I__2062\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18868\
        );

    \I__2061\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18868\
        );

    \I__2060\ : Odrv12
    port map (
            O => \N__18873\,
            I => \c0.data_in_frame_0_0\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__18868\,
            I => \c0.data_in_frame_0_0\
        );

    \I__2058\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18859\
        );

    \I__2057\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18856\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__18859\,
            I => \N__18850\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__2054\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18847\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__18850\,
            I => \N__18842\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__18847\,
            I => \N__18842\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__18842\,
            I => \c0.n2839\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \n1396_cascade_\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__18836\,
            I => \n2589_cascade_\
        );

    \I__2048\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__18830\,
            I => n2589
        );

    \I__2046\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__18818\,
            I => \c0.n18558\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__2041\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2039\ : Span4Mux_s3_v
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__18800\,
            I => \c0.n17797\
        );

    \I__2036\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__18794\,
            I => \N__18790\
        );

    \I__2034\ : InMux
    port map (
            O => \N__18793\,
            I => \N__18786\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__18790\,
            I => \N__18783\
        );

    \I__2032\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18780\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__18786\,
            I => \c0.n25_adj_2491\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__18783\,
            I => \c0.n25_adj_2491\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__18780\,
            I => \c0.n25_adj_2491\
        );

    \I__2028\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__18770\,
            I => \N__18764\
        );

    \I__2026\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18761\
        );

    \I__2025\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18758\
        );

    \I__2024\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18755\
        );

    \I__2023\ : Span4Mux_s2_h
    port map (
            O => \N__18764\,
            I => \N__18750\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18750\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__18758\,
            I => data_in_frame_5_5
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__18755\,
            I => data_in_frame_5_5
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__18750\,
            I => data_in_frame_5_5
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__2017\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18736\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__18739\,
            I => \N__18732\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__18736\,
            I => \N__18728\
        );

    \I__2014\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18725\
        );

    \I__2013\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18722\
        );

    \I__2012\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18719\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__18728\,
            I => \N__18714\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__18725\,
            I => \N__18714\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__18722\,
            I => \c0.data_in_frame_2_4\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__18719\,
            I => \c0.data_in_frame_2_4\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__18714\,
            I => \c0.data_in_frame_2_4\
        );

    \I__2006\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18700\
        );

    \I__2005\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__2004\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18697\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__18700\,
            I => \N__18694\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__18697\,
            I => \c0.data_in_frame_1_5\
        );

    \I__2001\ : Odrv12
    port map (
            O => \N__18694\,
            I => \c0.data_in_frame_1_5\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \n9419_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__18683\,
            I => \c0.n12_adj_2492\
        );

    \I__1997\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18675\
        );

    \I__1996\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18672\
        );

    \I__1995\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18669\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__18675\,
            I => \c0.data_in_frame_0_7\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__18672\,
            I => \c0.data_in_frame_0_7\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__18669\,
            I => \c0.data_in_frame_0_7\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__1990\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18654\
        );

    \I__1989\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18649\
        );

    \I__1988\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18649\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__18654\,
            I => \c0.data_in_frame_2_0\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__18649\,
            I => \c0.data_in_frame_2_0\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \c0.n17553_cascade_\
        );

    \I__1984\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18635\
        );

    \I__1983\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18632\
        );

    \I__1982\ : InMux
    port map (
            O => \N__18639\,
            I => \N__18629\
        );

    \I__1981\ : InMux
    port map (
            O => \N__18638\,
            I => \N__18626\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__18635\,
            I => \c0.data_in_frame_3_7\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__18632\,
            I => \c0.data_in_frame_3_7\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__18629\,
            I => \c0.data_in_frame_3_7\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18626\,
            I => \c0.data_in_frame_3_7\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__18617\,
            I => \c0.n17406_cascade_\
        );

    \I__1975\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__18611\,
            I => \c0.tx2.o_Tx_Serial_N_2354\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__18608\,
            I => \c0.tx2.n12306_cascade_\
        );

    \I__1972\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18600\
        );

    \I__1971\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18595\
        );

    \I__1970\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18595\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__18600\,
            I => \r_Clock_Count_0_adj_2634\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__18595\,
            I => \r_Clock_Count_0_adj_2634\
        );

    \I__1967\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18585\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18582\
        );

    \I__1965\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18579\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__18585\,
            I => \r_Clock_Count_2_adj_2632\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__18582\,
            I => \r_Clock_Count_2_adj_2632\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__18579\,
            I => \r_Clock_Count_2_adj_2632\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__18572\,
            I => \N__18567\
        );

    \I__1960\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18564\
        );

    \I__1959\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18559\
        );

    \I__1958\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18559\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__18564\,
            I => \r_Clock_Count_4_adj_2630\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__18559\,
            I => \r_Clock_Count_4_adj_2630\
        );

    \I__1955\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18549\
        );

    \I__1954\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18544\
        );

    \I__1953\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18544\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__18549\,
            I => \r_Clock_Count_3_adj_2631\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__18544\,
            I => \r_Clock_Count_3_adj_2631\
        );

    \I__1950\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18534\
        );

    \I__1949\ : InMux
    port map (
            O => \N__18538\,
            I => \N__18531\
        );

    \I__1948\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18528\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__18534\,
            I => \r_Clock_Count_5_adj_2629\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18531\,
            I => \r_Clock_Count_5_adj_2629\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__18528\,
            I => \r_Clock_Count_5_adj_2629\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__18521\,
            I => \c0.tx2.n10_cascade_\
        );

    \I__1943\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18513\
        );

    \I__1942\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18510\
        );

    \I__1941\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18507\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__18513\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__18510\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__18507\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1937\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18495\
        );

    \I__1936\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18492\
        );

    \I__1935\ : InMux
    port map (
            O => \N__18498\,
            I => \N__18489\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__18495\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__18492\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__18489\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1930\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18474\
        );

    \I__1929\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18469\
        );

    \I__1928\ : InMux
    port map (
            O => \N__18477\,
            I => \N__18469\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__18474\,
            I => \N__18466\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__18469\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__18466\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1924\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__18458\,
            I => \c0.tx2.n16452\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__18455\,
            I => \c0.tx2.r_SM_Main_2_N_2323_1_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__18449\,
            I => n320
        );

    \I__1919\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18435\
        );

    \I__1918\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18432\
        );

    \I__1917\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18423\
        );

    \I__1916\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18423\
        );

    \I__1915\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18423\
        );

    \I__1914\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18423\
        );

    \I__1913\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18420\
        );

    \I__1912\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18417\
        );

    \I__1911\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18414\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__18435\,
            I => n10244
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__18432\,
            I => n10244
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__18423\,
            I => n10244
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__18420\,
            I => n10244
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__18417\,
            I => n10244
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__18414\,
            I => n10244
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1903\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18393\
        );

    \I__1902\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18390\
        );

    \I__1901\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18387\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__18393\,
            I => \r_Clock_Count_1_adj_2633\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__18390\,
            I => \r_Clock_Count_1_adj_2633\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18387\,
            I => \r_Clock_Count_1_adj_2633\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__18380\,
            I => \c0.n18411_cascade_\
        );

    \I__1896\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18373\
        );

    \I__1895\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__18373\,
            I => data_out_frame2_18_6
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__18370\,
            I => data_out_frame2_18_6
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \c0.n18552_cascade_\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__18362\,
            I => \c0.n18555_cascade_\
        );

    \I__1890\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__18356\,
            I => \c0.n22_adj_2521\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__1887\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__18347\,
            I => n317
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__1884\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__18338\,
            I => n318
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__1881\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__18326\,
            I => n319
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__1877\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__18317\,
            I => n321
        );

    \I__1875\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18307\
        );

    \I__1873\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18304\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__18307\,
            I => \N__18301\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__18304\,
            I => data_out_frame2_5_0
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__18301\,
            I => data_out_frame2_5_0
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__18296\,
            I => \c0.n5_adj_2477_cascade_\
        );

    \I__1868\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__18287\,
            I => \c0.n6_adj_2436\
        );

    \I__1865\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18280\
        );

    \I__1864\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18277\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18274\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__18277\,
            I => data_out_frame2_18_1
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__18274\,
            I => data_out_frame2_18_1
        );

    \I__1860\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__18266\,
            I => \c0.n18468\
        );

    \I__1858\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18259\
        );

    \I__1857\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18256\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__18259\,
            I => data_out_frame2_5_1
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__18256\,
            I => data_out_frame2_5_1
        );

    \I__1854\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18247\
        );

    \I__1853\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18244\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__18244\,
            I => data_out_frame2_10_2
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__18241\,
            I => data_out_frame2_10_2
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__1848\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__18227\,
            I => \N__18223\
        );

    \I__1845\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__1844\ : Span4Mux_v
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__18220\,
            I => data_out_frame2_11_2
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__18217\,
            I => data_out_frame2_11_2
        );

    \I__1841\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18208\
        );

    \I__1840\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18205\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__18208\,
            I => data_out_frame2_12_0
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__18205\,
            I => data_out_frame2_12_0
        );

    \I__1837\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__1835\ : Odrv12
    port map (
            O => \N__18194\,
            I => \c0.n17794\
        );

    \I__1834\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__18179\,
            I => \c0.n18078\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \c0.n18408_cascade_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__1826\ : Span12Mux_v
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__1825\ : Odrv12
    port map (
            O => \N__18164\,
            I => \c0.n6_adj_2506\
        );

    \I__1824\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__18158\,
            I => \c0.n5_adj_2495\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__1821\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__18149\,
            I => \N__18145\
        );

    \I__1819\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18142\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__18145\,
            I => \N__18139\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__18142\,
            I => data_out_frame2_5_5
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__18139\,
            I => data_out_frame2_5_5
        );

    \I__1815\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__1813\ : Span4Mux_s1_h
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__18125\,
            I => \c0.n6_adj_2496\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__18122\,
            I => \N__18118\
        );

    \I__1810\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__1809\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18112\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__18115\,
            I => data_out_frame2_11_3
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__18112\,
            I => data_out_frame2_11_3
        );

    \I__1806\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__18101\,
            I => \c0.n17629\
        );

    \I__1803\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__1801\ : Span4Mux_h
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__18083\,
            I => \c0.n8725\
        );

    \I__1797\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18076\
        );

    \I__1796\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18073\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__18076\,
            I => data_out_frame2_10_0
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__18073\,
            I => data_out_frame2_10_0
        );

    \I__1793\ : InMux
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18061\
        );

    \I__1791\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18058\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__18061\,
            I => \N__18055\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__18058\,
            I => data_out_frame2_17_0
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__18055\,
            I => data_out_frame2_17_0
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18043\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18040\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__18037\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__18040\,
            I => data_out_frame2_16_0
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__18037\,
            I => data_out_frame2_16_0
        );

    \I__1781\ : InMux
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__18029\,
            I => \c0.n18600\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__18026\,
            I => \N__18022\
        );

    \I__1778\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18017\
        );

    \I__1777\ : InMux
    port map (
            O => \N__18022\,
            I => \N__18017\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__18017\,
            I => data_out_frame2_8_6
        );

    \I__1775\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__1773\ : Span12Mux_s7_v
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__18005\,
            I => \c0.n18564\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__1770\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17995\
        );

    \I__1769\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17992\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__17995\,
            I => \N__17989\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__17992\,
            I => \N__17984\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__17989\,
            I => \N__17984\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__17984\,
            I => data_out_frame2_16_1
        );

    \I__1764\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17974\
        );

    \I__1762\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__1761\ : Span4Mux_s1_h
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__17971\,
            I => data_out_frame2_17_1
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__17968\,
            I => data_out_frame2_17_1
        );

    \I__1758\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17959\
        );

    \I__1757\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17956\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__17959\,
            I => data_out_frame2_18_0
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__17956\,
            I => data_out_frame2_18_0
        );

    \I__1754\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17947\
        );

    \I__1753\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17944\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__17947\,
            I => data_out_frame2_10_3
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__17944\,
            I => data_out_frame2_10_3
        );

    \I__1750\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17935\
        );

    \I__1749\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17932\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__17935\,
            I => data_out_frame2_14_4
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__17932\,
            I => data_out_frame2_14_4
        );

    \I__1746\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17924\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__1744\ : Span4Mux_h
    port map (
            O => \N__17921\,
            I => \N__17917\
        );

    \I__1743\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17914\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__17917\,
            I => \N__17911\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__17914\,
            I => data_out_frame2_7_6
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__17911\,
            I => data_out_frame2_7_6
        );

    \I__1739\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17902\
        );

    \I__1738\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17899\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__17902\,
            I => data_out_frame2_8_5
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__17899\,
            I => data_out_frame2_8_5
        );

    \I__1735\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17890\
        );

    \I__1734\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17887\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__17890\,
            I => \N__17884\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__17887\,
            I => data_out_frame2_15_1
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__17884\,
            I => data_out_frame2_15_1
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__1729\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17872\
        );

    \I__1728\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17869\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__17872\,
            I => \N__17866\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__17869\,
            I => data_out_frame2_11_6
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__17866\,
            I => data_out_frame2_11_6
        );

    \I__1724\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17857\
        );

    \I__1723\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17854\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__17857\,
            I => \N__17851\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__17854\,
            I => data_out_frame2_15_6
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__17851\,
            I => data_out_frame2_15_6
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__1718\ : InMux
    port map (
            O => \N__17843\,
            I => \N__17839\
        );

    \I__1717\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17836\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__17839\,
            I => \N__17833\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__17836\,
            I => data_out_frame2_5_2
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__17833\,
            I => data_out_frame2_5_2
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__1712\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17821\
        );

    \I__1711\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17818\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__17821\,
            I => \N__17815\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__17818\,
            I => data_out_frame2_15_2
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__17815\,
            I => data_out_frame2_15_2
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__1706\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17803\
        );

    \I__1705\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17800\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17797\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__17800\,
            I => data_out_frame2_15_0
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__17797\,
            I => data_out_frame2_15_0
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__1700\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17783\
        );

    \I__1699\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17783\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__17783\,
            I => data_out_frame2_13_2
        );

    \I__1697\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__1695\ : Span4Mux_h
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__17771\,
            I => \c0.n18492\
        );

    \I__1693\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17765\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__17765\,
            I => \N__17762\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__17762\,
            I => \c0.n17827\
        );

    \I__1690\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__1689\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17753\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__17753\,
            I => data_out_frame2_12_5
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__17750\,
            I => \c0.n9043_cascade_\
        );

    \I__1686\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17744\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17740\
        );

    \I__1684\ : InMux
    port map (
            O => \N__17743\,
            I => \N__17737\
        );

    \I__1683\ : Span12Mux_v
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__17737\,
            I => data_out_frame2_14_6
        );

    \I__1681\ : Odrv12
    port map (
            O => \N__17734\,
            I => data_out_frame2_14_6
        );

    \I__1680\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__17726\,
            I => \N__17722\
        );

    \I__1678\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17719\
        );

    \I__1677\ : Sp12to4
    port map (
            O => \N__17722\,
            I => \N__17716\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__17719\,
            I => data_out_frame2_10_6
        );

    \I__1675\ : Odrv12
    port map (
            O => \N__17716\,
            I => data_out_frame2_10_6
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__1673\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17705\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17701\
        );

    \I__1671\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17698\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__17701\,
            I => \N__17695\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__17698\,
            I => data_out_frame2_11_0
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__17695\,
            I => data_out_frame2_11_0
        );

    \I__1667\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__17681\,
            I => \N__17677\
        );

    \I__1663\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__17677\,
            I => \N__17671\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__17674\,
            I => data_out_frame2_6_6
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__17671\,
            I => data_out_frame2_6_6
        );

    \I__1659\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__1657\ : Odrv12
    port map (
            O => \N__17660\,
            I => \c0.n9_adj_2507\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__17657\,
            I => \c0.n17325_cascade_\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__17654\,
            I => \c0.n8_adj_2459_cascade_\
        );

    \I__1654\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__17648\,
            I => \c0.n2604\
        );

    \I__1652\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__17642\,
            I => \c0.n11_adj_2460\
        );

    \I__1650\ : CEMux
    port map (
            O => \N__17639\,
            I => \N__17636\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__1648\ : Span4Mux_s2_h
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__17630\,
            I => \c0.n9605\
        );

    \I__1646\ : SRMux
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__17624\,
            I => \c0.n9900\
        );

    \I__1644\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__17618\,
            I => \c0.n17806\
        );

    \I__1642\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17611\
        );

    \I__1641\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17608\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__17611\,
            I => data_out_frame2_18_5
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__17608\,
            I => data_out_frame2_18_5
        );

    \I__1638\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17600\,
            I => \c0.n2607\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__1635\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__17591\,
            I => \c0.n17513\
        );

    \I__1633\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__17585\,
            I => \c0.n2602\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__1630\ : InMux
    port map (
            O => \N__17579\,
            I => \N__17569\
        );

    \I__1629\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17569\
        );

    \I__1628\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17569\
        );

    \I__1627\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17566\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__17569\,
            I => \N__17563\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__17566\,
            I => \c0.data_in_frame_3_2\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__17563\,
            I => \c0.data_in_frame_3_2\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__1622\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__17552\,
            I => \c0.n9_adj_2500\
        );

    \I__1620\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17545\
        );

    \I__1619\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17542\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__17545\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17542\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__17537\,
            I => \N__17533\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__17536\,
            I => \N__17530\
        );

    \I__1614\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17527\
        );

    \I__1613\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17524\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__17527\,
            I => \c0.data_in_frame_3_3\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__17524\,
            I => \c0.data_in_frame_3_3\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__17519\,
            I => \c0.n17629_cascade_\
        );

    \I__1609\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__17513\,
            I => \c0.n16_adj_2546\
        );

    \I__1607\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__17507\,
            I => \c0.n9254\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__17504\,
            I => \c0.n9254_cascade_\
        );

    \I__1604\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__1603\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17489\
        );

    \I__1602\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17489\
        );

    \I__1601\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17486\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__17495\,
            I => \N__17483\
        );

    \I__1599\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17480\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__17489\,
            I => \c0.data_in_frame_2_5\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__17486\,
            I => \c0.data_in_frame_2_5\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__17483\,
            I => \c0.data_in_frame_2_5\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__17480\,
            I => \c0.data_in_frame_2_5\
        );

    \I__1594\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17467\
        );

    \I__1593\ : InMux
    port map (
            O => \N__17470\,
            I => \N__17464\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__17467\,
            I => \c0.n8976\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__17464\,
            I => \c0.n8976\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__1589\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__17453\,
            I => \N__17448\
        );

    \I__1587\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17443\
        );

    \I__1586\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17443\
        );

    \I__1585\ : Odrv12
    port map (
            O => \N__17448\,
            I => \c0.data_in_frame_1_3\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__17443\,
            I => \c0.data_in_frame_1_3\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__1582\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__1580\ : Span4Mux_v
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__17426\,
            I => \c0.n5_adj_2515\
        );

    \I__1578\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17420\,
            I => \c0.n17507\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \c0.n17476_cascade_\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17411\,
            I => \c0.n17476\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__17408\,
            I => \c0.n17478_cascade_\
        );

    \I__1572\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__17402\,
            I => n316
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__17399\,
            I => \c0.n17507_cascade_\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__1568\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17385\
        );

    \I__1567\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17385\
        );

    \I__1566\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17382\
        );

    \I__1565\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17379\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__17385\,
            I => \c0.data_in_frame_0_4\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__17382\,
            I => \c0.data_in_frame_0_4\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__17379\,
            I => \c0.data_in_frame_0_4\
        );

    \I__1561\ : InMux
    port map (
            O => \N__17372\,
            I => \c0.tx2.n16374\
        );

    \I__1560\ : InMux
    port map (
            O => \N__17369\,
            I => \c0.tx2.n16375\
        );

    \I__1559\ : InMux
    port map (
            O => \N__17366\,
            I => \c0.tx2.n16376\
        );

    \I__1558\ : InMux
    port map (
            O => \N__17363\,
            I => \c0.tx2.n16377\
        );

    \I__1557\ : InMux
    port map (
            O => \N__17360\,
            I => \c0.tx2.n16378\
        );

    \I__1556\ : InMux
    port map (
            O => \N__17357\,
            I => \bfn_1_32_0_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__17351\,
            I => \c0.tx2.n17953\
        );

    \I__1553\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__17345\,
            I => \c0.tx2.n18013\
        );

    \I__1551\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__17339\,
            I => \c0.tx2.n17939\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__17336\,
            I => \c0.n18435_cascade_\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__17333\,
            I => \N__17330\
        );

    \I__1547\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__1545\ : Span12Mux_s3_v
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__17321\,
            I => \c0.n17836\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__17318\,
            I => \c0.n18360_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17309\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__17309\,
            I => \c0.n6_adj_2504\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__17306\,
            I => \c0.n18471_cascade_\
        );

    \I__1538\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__17300\,
            I => \c0.n18363\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \c0.n22_adj_2530_cascade_\
        );

    \I__1535\ : InMux
    port map (
            O => \N__17294\,
            I => \bfn_1_31_0_\
        );

    \I__1534\ : InMux
    port map (
            O => \N__17291\,
            I => \c0.tx2.n16372\
        );

    \I__1533\ : InMux
    port map (
            O => \N__17288\,
            I => \c0.tx2.n16373\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__17285\,
            I => \c0.n5_adj_2503_cascade_\
        );

    \I__1531\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17276\
        );

    \I__1530\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17276\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__17276\,
            I => data_out_frame2_14_2
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__17273\,
            I => \c0.n18606_cascade_\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \c0.n18570_cascade_\
        );

    \I__1526\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__17264\,
            I => \c0.n17779\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__17261\,
            I => \c0.n17773_cascade_\
        );

    \I__1523\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__17252\,
            I => \c0.n18074\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__17249\,
            I => \c0.n18432_cascade_\
        );

    \I__1519\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17242\
        );

    \I__1518\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__17242\,
            I => \N__17236\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__17239\,
            I => data_out_frame2_16_2
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__17236\,
            I => data_out_frame2_16_2
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \c0.n18486_cascade_\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \c0.n18489_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__17222\,
            I => \c0.n18084\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__17219\,
            I => \c0.n18366_cascade_\
        );

    \I__1509\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__17210\,
            I => \c0.n6_adj_2466\
        );

    \I__1506\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__17204\,
            I => \c0.n22_adj_2529\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__17201\,
            I => \c0.n18369_cascade_\
        );

    \I__1503\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17194\
        );

    \I__1502\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__17191\,
            I => data_out_frame2_7_5
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__17188\,
            I => data_out_frame2_7_5
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__17183\,
            I => \c0.n18387_cascade_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__17174\,
            I => \c0.n5_adj_2463\
        );

    \I__1494\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17167\
        );

    \I__1493\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__17167\,
            I => data_out_frame2_16_5
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__17164\,
            I => data_out_frame2_16_5
        );

    \I__1490\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17155\
        );

    \I__1489\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__17152\,
            I => data_out_frame2_9_5
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__17149\,
            I => data_out_frame2_9_5
        );

    \I__1485\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__17141\,
            I => \N__17137\
        );

    \I__1483\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__1482\ : Span4Mux_s1_h
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__17134\,
            I => data_out_frame2_6_2
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__17131\,
            I => data_out_frame2_6_2
        );

    \I__1479\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__17123\,
            I => \c0.n18474\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__17120\,
            I => \c0.n18534_cascade_\
        );

    \I__1476\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17113\
        );

    \I__1475\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17110\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__17113\,
            I => data_out_frame2_17_5
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__17110\,
            I => data_out_frame2_17_5
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__17105\,
            I => \c0.n18537_cascade_\
        );

    \I__1471\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__17099\,
            I => \c0.n17803\
        );

    \I__1469\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17093\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__17093\,
            I => \N__17090\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__17090\,
            I => \c0.n18080\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__17087\,
            I => \c0.n18384_cascade_\
        );

    \I__1465\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__17081\,
            I => \c0.n22_adj_2523\
        );

    \I__1463\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17072\
        );

    \I__1462\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17072\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__17072\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__1460\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17063\
        );

    \I__1459\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17063\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__17063\,
            I => data_out_frame2_7_2
        );

    \I__1457\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17056\
        );

    \I__1456\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17053\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17050\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__17053\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__17050\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__17045\,
            I => \c0.n18546_cascade_\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \N__17038\
        );

    \I__1450\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17033\
        );

    \I__1449\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17033\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__17033\,
            I => data_out_frame2_11_5
        );

    \I__1447\ : InMux
    port map (
            O => \N__17030\,
            I => \c0.n16405\
        );

    \I__1446\ : InMux
    port map (
            O => \N__17027\,
            I => \c0.n16406\
        );

    \I__1445\ : InMux
    port map (
            O => \N__17024\,
            I => \c0.n16407\
        );

    \I__1444\ : InMux
    port map (
            O => \N__17021\,
            I => \c0.n16408\
        );

    \I__1443\ : InMux
    port map (
            O => \N__17018\,
            I => \c0.n16409\
        );

    \I__1442\ : InMux
    port map (
            O => \N__17015\,
            I => \c0.n16410\
        );

    \I__1441\ : InMux
    port map (
            O => \N__17012\,
            I => \c0.n16411\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__17009\,
            I => \c0.n20_adj_2547_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__16999\
        );

    \I__1437\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__16999\,
            I => \c0.n9317\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__16996\,
            I => \c0.n9317\
        );

    \I__1434\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__16988\,
            I => \c0.n8063\
        );

    \I__1432\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__16982\,
            I => \c0.n17650\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__16979\,
            I => \c0.n8645_cascade_\
        );

    \I__1429\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__16970\,
            I => \c0.n9186\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__16967\,
            I => \c0.n30_adj_2489_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__16961\,
            I => \c0.n18_adj_2545\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__16958\,
            I => \c0.n9186_cascade_\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__16955\,
            I => \c0.n8857_cascade_\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \c0.n8725_cascade_\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__16949\,
            I => \c0.n8063_cascade_\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__16946\,
            I => \N__16942\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__16945\,
            I => \N__16938\
        );

    \I__1417\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16928\
        );

    \I__1416\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16928\
        );

    \I__1415\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16928\
        );

    \I__1414\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16928\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__16928\,
            I => \c0.data_in_frame_0_3\
        );

    \I__1412\ : IoInMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__1410\ : IoSpan4Mux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__1409\ : IoSpan4Mux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__1408\ : IoSpan4Mux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__16910\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_9_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_29_0_\
        );

    \IN_MUX_bfv_9_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16419,
            carryinitout => \bfn_9_30_0_\
        );

    \IN_MUX_bfv_9_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16427,
            carryinitout => \bfn_9_31_0_\
        );

    \IN_MUX_bfv_9_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16435,
            carryinitout => \bfn_9_32_0_\
        );

    \IN_MUX_bfv_5_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_29_0_\
        );

    \IN_MUX_bfv_5_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16326,
            carryinitout => \bfn_5_30_0_\
        );

    \IN_MUX_bfv_5_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16334,
            carryinitout => \bfn_5_31_0_\
        );

    \IN_MUX_bfv_5_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16342,
            carryinitout => \bfn_5_32_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n16379\,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n16364\,
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_6_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_30_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16312\,
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_16_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_29_0_\
        );

    \IN_MUX_bfv_16_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16387,
            carryinitout => \bfn_16_30_0_\
        );

    \IN_MUX_bfv_16_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16395,
            carryinitout => \bfn_16_31_0_\
        );

    \IN_MUX_bfv_16_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16403,
            carryinitout => \bfn_16_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16925\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_998_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29030\,
            in1 => \N__21728\,
            in2 => \_gnd_net_\,
            in3 => \N__17501\,
            lcout => \c0.n17602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_995_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29011\,
            in1 => \_gnd_net_\,
            in2 => \N__16945\,
            in3 => \N__22168\,
            lcout => \c0.n9163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45511\,
            in1 => \N__27778\,
            in2 => \_gnd_net_\,
            in3 => \N__27719\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i33_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22103\,
            in1 => \N__27850\,
            in2 => \_gnd_net_\,
            in3 => \N__45512\,
            lcout => data_in_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_945_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16937\,
            in2 => \_gnd_net_\,
            in3 => \N__29010\,
            lcout => \c0.n17550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i4_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__27611\,
            in1 => \N__24272\,
            in2 => \N__16946\,
            in3 => \N__31976\,
            lcout => \c0.data_in_frame_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_987_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17392\,
            in2 => \_gnd_net_\,
            in3 => \N__16941\,
            lcout => \c0.n22_adj_2508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i5_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__21629\,
            in1 => \N__24273\,
            in2 => \N__17396\,
            in3 => \N__31977\,
            lcout => \c0.data_in_frame_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i18_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24271\,
            in1 => \N__31418\,
            in2 => \N__29040\,
            in3 => \N__31975\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_988_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29031\,
            in2 => \_gnd_net_\,
            in3 => \N__21718\,
            lcout => \c0.n9186\,
            ltout => \c0.n9186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1015_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20556\,
            in1 => \N__18797\,
            in2 => \N__16958\,
            in3 => \N__18773\,
            lcout => \c0.n8857\,
            ltout => \c0.n8857_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_931_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20072\,
            in1 => \N__23022\,
            in2 => \N__16955\,
            in3 => \N__22229\,
            lcout => \c0.n17541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_996_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20482\,
            in1 => \N__20071\,
            in2 => \N__25589\,
            in3 => \N__20425\,
            lcout => \c0.n8725\,
            ltout => \c0.n8725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_864_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17510\,
            in1 => \N__25025\,
            in2 => \N__16952\,
            in3 => \N__17006\,
            lcout => \c0.n17594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1024_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20424\,
            lcout => \c0.n9176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_960_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24673\,
            lcout => \c0.n8063\,
            ltout => \c0.n8063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1115_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__22450\,
            in2 => \N__16949\,
            in3 => \N__16964\,
            lcout => OPEN,
            ltout => \c0.n20_adj_2547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1116_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17002\,
            in1 => \N__20600\,
            in2 => \N__17009\,
            in3 => \N__17516\,
            lcout => \c0.n8056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i49_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23823\,
            in1 => \_gnd_net_\,
            in2 => \N__24605\,
            in3 => \N__45481\,
            lcout => data_in_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_857_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22002\,
            in1 => \N__28759\,
            in2 => \_gnd_net_\,
            in3 => \N__17498\,
            lcout => \c0.n9317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_958_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28760\,
            in1 => \N__22406\,
            in2 => \N__27518\,
            in3 => \N__16991\,
            lcout => \c0.n17544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_952_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25583\,
            in2 => \_gnd_net_\,
            in3 => \N__20073\,
            lcout => \c0.n17650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_830_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19958\,
            in1 => \N__17452\,
            in2 => \N__17536\,
            in3 => \N__19859\,
            lcout => \c0.n8645\,
            ltout => \c0.n8645_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1089_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18706\,
            in1 => \N__17577\,
            in2 => \N__16979\,
            in3 => \N__19871\,
            lcout => \c0.n30_adj_2489\,
            ltout => \c0.n30_adj_2489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1108_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16976\,
            in1 => \N__22333\,
            in2 => \N__16967\,
            in3 => \N__17470\,
            lcout => \c0.n18_adj_2545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_2_lut_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17578\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17451\,
            lcout => \c0.n9365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i7_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__33170\,
            in1 => \N__17059\,
            in2 => \N__33678\,
            in3 => \N__23873\,
            lcout => \c0.data_out_frame2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1090_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19959\,
            in1 => \N__22139\,
            in2 => \N__17582\,
            in3 => \N__18707\,
            lcout => \c0.n17516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1074_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22225\,
            in1 => \N__23793\,
            in2 => \N__20074\,
            in3 => \N__22831\,
            lcout => \c0.n9204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1034_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24955\,
            in2 => \_gnd_net_\,
            in3 => \N__21582\,
            lcout => \c0.n9328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15831_3_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__17548\,
            in1 => \N__30985\,
            in2 => \_gnd_net_\,
            in3 => \N__30564\,
            lcout => \c0.n18080\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i43_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__24721\,
            in1 => \N__24274\,
            in2 => \N__33038\,
            in3 => \N__31918\,
            lcout => data_in_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i81_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24415\,
            in2 => \_gnd_net_\,
            in3 => \N__31917\,
            lcout => \c0.data_in_frame_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1051_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24720\,
            in1 => \N__24956\,
            in2 => \_gnd_net_\,
            in3 => \N__21583\,
            lcout => \c0.n8976\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_832_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__22553\,
            in1 => \_gnd_net_\,
            in2 => \N__21946\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2272__i0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19619\,
            in2 => \N__30625\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => \c0.n16405\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i1_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30930\,
            in2 => \_gnd_net_\,
            in3 => \N__17030\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n16405\,
            carryout => \c0.n16406\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i2_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26758\,
            in2 => \_gnd_net_\,
            in3 => \N__17027\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \c0.n16406\,
            carryout => \c0.n16407\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__17024\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \c0.n16407\,
            carryout => \c0.n16408\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i4_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26455\,
            in2 => \_gnd_net_\,
            in3 => \N__17021\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \c0.n16408\,
            carryout => \c0.n16409\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19687\,
            in2 => \_gnd_net_\,
            in3 => \N__17018\,
            lcout => \c0.byte_transmit_counter2_5\,
            ltout => OPEN,
            carryin => \c0.n16409\,
            carryout => \c0.n16410\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i6_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19663\,
            in2 => \_gnd_net_\,
            in3 => \N__17015\,
            lcout => \c0.byte_transmit_counter2_6\,
            ltout => OPEN,
            carryin => \c0.n16410\,
            carryout => \c0.n16411\,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_2272__i7_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19636\,
            in2 => \_gnd_net_\,
            in3 => \N__17012\,
            lcout => \c0.byte_transmit_counter2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50266\,
            ce => \N__17639\,
            sr => \N__17627\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16006_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__17894\,
            in1 => \N__25316\,
            in2 => \N__30964\,
            in3 => \N__30560\,
            lcout => \c0.n18474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i131_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32816\,
            in1 => \N__34112\,
            in2 => \_gnd_net_\,
            in3 => \N__17245\,
            lcout => data_out_frame2_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15805_3_lut_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__30875\,
            in1 => \N__17077\,
            in2 => \_gnd_net_\,
            in3 => \N__30563\,
            lcout => \c0.n18074\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i1_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__17078\,
            in1 => \N__33159\,
            in2 => \N__33692\,
            in3 => \N__23881\,
            lcout => \c0.data_out_frame2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1080_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20380\,
            in1 => \N__18936\,
            in2 => \_gnd_net_\,
            in3 => \N__22960\,
            lcout => n9380,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i59_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32817\,
            in1 => \N__34769\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => data_out_frame2_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17068\,
            in1 => \N__17144\,
            in2 => \_gnd_net_\,
            in3 => \N__30561\,
            lcout => \c0.n5_adj_2463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15818_3_lut_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__30562\,
            in1 => \N__17060\,
            in2 => \_gnd_net_\,
            in3 => \N__30874\,
            lcout => \c0.n18078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16066_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19118\,
            in1 => \N__30979\,
            in2 => \N__17042\,
            in3 => \N__30669\,
            lcout => OPEN,
            ltout => \c0.n18546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18546_bdd_4_lut_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30980\,
            in1 => \N__17905\,
            in2 => \N__17045\,
            in3 => \N__17159\,
            lcout => \c0.n17803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i91_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34765\,
            in1 => \N__18226\,
            in2 => \_gnd_net_\,
            in3 => \N__32821\,
            lcout => data_out_frame2_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i94_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32819\,
            in1 => \N__35603\,
            in2 => \_gnd_net_\,
            in3 => \N__17041\,
            lcout => data_out_frame2_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3957_3_lut_4_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20143\,
            in1 => \N__34684\,
            in2 => \N__23702\,
            in3 => \N__28066\,
            lcout => \c0.n2604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18474_bdd_4_lut_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__30978\,
            in1 => \N__17126\,
            in2 => \N__19160\,
            in3 => \N__18998\,
            lcout => \c0.n17836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i109_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19540\,
            in1 => \N__36463\,
            in2 => \_gnd_net_\,
            in3 => \N__32820\,
            lcout => data_out_frame2_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i142_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32818\,
            in1 => \N__35602\,
            in2 => \_gnd_net_\,
            in3 => \N__17117\,
            lcout => data_out_frame2_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16056_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__17614\,
            in1 => \N__30986\,
            in2 => \N__20849\,
            in3 => \N__30670\,
            lcout => OPEN,
            ltout => \c0.n18534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18534_bdd_4_lut_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30987\,
            in1 => \N__17170\,
            in2 => \N__17120\,
            in3 => \N__17116\,
            lcout => OPEN,
            ltout => \c0.n18537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26782\,
            in1 => \N__19025\,
            in2 => \N__17105\,
            in3 => \N__26942\,
            lcout => \c0.n22_adj_2523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15950_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__17621\,
            in1 => \N__26783\,
            in2 => \N__26667\,
            in3 => \N__17102\,
            lcout => OPEN,
            ltout => \c0.n18384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18384_bdd_4_lut_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__26624\,
            in1 => \N__17096\,
            in2 => \N__17087\,
            in3 => \N__18134\,
            lcout => OPEN,
            ltout => \c0.n18387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17084\,
            in1 => \N__26625\,
            in2 => \N__17183\,
            in3 => \N__26476\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50285\,
            ce => \N__26400\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__30988\,
            in1 => \N__17180\,
            in2 => \N__17846\,
            in3 => \N__30672\,
            lcout => \c0.n6_adj_2466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15824_3_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__30673\,
            in1 => \_gnd_net_\,
            in2 => \N__23249\,
            in3 => \N__30989\,
            lcout => \c0.n18084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i46_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36409\,
            in1 => \N__18148\,
            in2 => \_gnd_net_\,
            in3 => \N__32651\,
            lcout => data_out_frame2_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i62_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32648\,
            in1 => \N__35595\,
            in2 => \_gnd_net_\,
            in3 => \N__17197\,
            lcout => data_out_frame2_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i134_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35099\,
            in1 => \N__17171\,
            in2 => \_gnd_net_\,
            in3 => \N__32650\,
            lcout => data_out_frame2_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i78_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32649\,
            in1 => \N__36410\,
            in2 => \_gnd_net_\,
            in3 => \N__17158\,
            lcout => data_out_frame2_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1128_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36547\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \c0.n6_adj_2550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i51_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32647\,
            in1 => \N__35306\,
            in2 => \_gnd_net_\,
            in3 => \N__17140\,
            lcout => data_out_frame2_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16016_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__20816\,
            in1 => \N__31033\,
            in2 => \N__29156\,
            in3 => \N__30671\,
            lcout => OPEN,
            ltout => \c0.n18486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18486_bdd_4_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31034\,
            in1 => \N__17246\,
            in2 => \N__17231\,
            in3 => \N__19208\,
            lcout => OPEN,
            ltout => \c0.n18489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26843\,
            in1 => \N__20861\,
            in2 => \N__17228\,
            in3 => \N__26906\,
            lcout => \c0.n22_adj_2529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15921_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__19352\,
            in1 => \N__17768\,
            in2 => \N__26662\,
            in3 => \N__26844\,
            lcout => OPEN,
            ltout => \c0.n18366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18366_bdd_4_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__26626\,
            in1 => \N__17225\,
            in2 => \N__17219\,
            in3 => \N__17216\,
            lcout => OPEN,
            ltout => \c0.n18369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17207\,
            in1 => \N__26627\,
            in2 => \N__17201\,
            in3 => \N__26500\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50298\,
            ce => \N__26409\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30766\,
            in1 => \_gnd_net_\,
            in2 => \N__19181\,
            in3 => \N__17198\,
            lcout => \c0.n5_adj_2495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20996\,
            in1 => \N__30761\,
            in2 => \_gnd_net_\,
            in3 => \N__17938\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16026_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__30760\,
            in1 => \N__17281\,
            in2 => \N__17828\,
            in3 => \N__30965\,
            lcout => \c0.n18492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19310\,
            in1 => \N__30764\,
            in2 => \_gnd_net_\,
            in3 => \N__19229\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__30765\,
            in1 => \N__18262\,
            in2 => \N__17285\,
            in3 => \N__30968\,
            lcout => \c0.n6_adj_2504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16046_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__30967\,
            in1 => \N__30763\,
            in2 => \N__18122\,
            in3 => \N__17950\,
            lcout => \c0.n18522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16110_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__30762\,
            in1 => \N__30966\,
            in2 => \N__19484\,
            in3 => \N__17962\,
            lcout => \c0.n18600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i115_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17282\,
            in1 => \N__35298\,
            in2 => \_gnd_net_\,
            in3 => \N__32796\,
            lcout => data_out_frame2_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__20834\,
            in1 => \N__30981\,
            in2 => \N__17810\,
            in3 => \N__30738\,
            lcout => OPEN,
            ltout => \c0.n18606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18606_bdd_4_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30982\,
            in1 => \N__18211\,
            in2 => \N__17273\,
            in3 => \N__30047\,
            lcout => \c0.n17779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16086_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18079\,
            in1 => \N__30983\,
            in2 => \N__17711\,
            in3 => \N__30739\,
            lcout => OPEN,
            ltout => \c0.n18570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18570_bdd_4_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__30984\,
            in1 => \N__20945\,
            in2 => \N__17270\,
            in3 => \N__19082\,
            lcout => OPEN,
            ltout => \c0.n17773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__17267\,
            in1 => \N__26619\,
            in2 => \N__17261\,
            in3 => \N__26784\,
            lcout => OPEN,
            ltout => \c0.n18432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18432_bdd_4_lut_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__17258\,
            in1 => \N__26661\,
            in2 => \N__17249\,
            in3 => \N__18293\,
            lcout => OPEN,
            ltout => \c0.n18435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__19454\,
            in1 => \N__26620\,
            in2 => \N__17336\,
            in3 => \N__26501\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50314\,
            ce => \N__26405\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15916_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19241\,
            in1 => \N__26616\,
            in2 => \N__17333\,
            in3 => \N__26780\,
            lcout => OPEN,
            ltout => \c0.n18360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18360_bdd_4_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__26617\,
            in1 => \N__30488\,
            in2 => \N__17318\,
            in3 => \N__17315\,
            lcout => \c0.n18363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18468_bdd_4_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__17981\,
            in1 => \N__18269\,
            in2 => \N__18002\,
            in3 => \N__30990\,
            lcout => OPEN,
            ltout => \c0.n18471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26781\,
            in1 => \N__21044\,
            in2 => \N__17306\,
            in3 => \N__26933\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17303\,
            in1 => \N__26618\,
            in2 => \N__17297\,
            in3 => \N__26518\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50323\,
            ce => \N__26378\,
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_2_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18605\,
            in2 => \_gnd_net_\,
            in3 => \N__17294\,
            lcout => n321,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => \c0.tx2.n16372\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_3_lut_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18397\,
            in2 => \_gnd_net_\,
            in3 => \N__17291\,
            lcout => n320,
            ltout => OPEN,
            carryin => \c0.tx2.n16372\,
            carryout => \c0.tx2.n16373\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_4_lut_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18589\,
            in2 => \_gnd_net_\,
            in3 => \N__17288\,
            lcout => n319,
            ltout => OPEN,
            carryin => \c0.tx2.n16373\,
            carryout => \c0.tx2.n16374\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_5_lut_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18554\,
            in2 => \_gnd_net_\,
            in3 => \N__17372\,
            lcout => n318,
            ltout => OPEN,
            carryin => \c0.tx2.n16374\,
            carryout => \c0.tx2.n16375\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_6_lut_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18571\,
            in2 => \_gnd_net_\,
            in3 => \N__17369\,
            lcout => n317,
            ltout => OPEN,
            carryin => \c0.tx2.n16375\,
            carryout => \c0.tx2.n16376\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_7_lut_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18538\,
            in2 => \_gnd_net_\,
            in3 => \N__17366\,
            lcout => n316,
            ltout => OPEN,
            carryin => \c0.tx2.n16376\,
            carryout => \c0.tx2.n16377\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_8_lut_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18440\,
            in1 => \N__18499\,
            in2 => \_gnd_net_\,
            in3 => \N__17363\,
            lcout => \c0.tx2.n18013\,
            ltout => OPEN,
            carryin => \c0.tx2.n16377\,
            carryout => \c0.tx2.n16378\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_9_lut_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18438\,
            in1 => \N__18517\,
            in2 => \_gnd_net_\,
            in3 => \N__17360\,
            lcout => \c0.tx2.n17953\,
            ltout => OPEN,
            carryin => \c0.tx2.n16378\,
            carryout => \c0.tx2.n16379\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.add_59_10_lut_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18439\,
            in1 => \N__18477\,
            in2 => \_gnd_net_\,
            in3 => \N__17357\,
            lcout => \c0.tx2.n17939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i7_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17354\,
            in1 => \N__21416\,
            in2 => \_gnd_net_\,
            in3 => \N__18518\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i6_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21415\,
            in1 => \N__18500\,
            in2 => \_gnd_net_\,
            in3 => \N__17348\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i8_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18478\,
            in1 => \N__21417\,
            in2 => \_gnd_net_\,
            in3 => \N__17342\,
            lcout => \c0.tx2.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i5_LC_1_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__17405\,
            in1 => \N__18539\,
            in2 => \N__21432\,
            in3 => \N__18445\,
            lcout => \r_Clock_Count_5_adj_2629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_4_lut_4_lut_LC_1_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__21340\,
            in1 => \N__21266\,
            in2 => \N__21431\,
            in3 => \N__21470\,
            lcout => n10244,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16081_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__31030\,
            in1 => \N__17729\,
            in2 => \N__17879\,
            in3 => \N__30645\,
            lcout => \c0.n18564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_991_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17391\,
            in1 => \N__21858\,
            in2 => \_gnd_net_\,
            in3 => \N__20426\,
            lcout => \c0.n17507\,
            ltout => \c0.n17507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_914_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21772\,
            in1 => \N__19784\,
            in2 => \N__17399\,
            in3 => \N__18735\,
            lcout => \c0.n8687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17927\,
            in1 => \N__17690\,
            in2 => \_gnd_net_\,
            in3 => \N__30644\,
            lcout => \c0.n5_adj_2515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i36_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__20427\,
            in1 => \N__24218\,
            in2 => \N__27578\,
            in3 => \N__31979\,
            lcout => \c0.data_in_frame_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50252\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1047_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17390\,
            in2 => \_gnd_net_\,
            in3 => \N__21857\,
            lcout => \c0.n20_adj_2427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16076_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__30643\,
            in1 => \N__17747\,
            in2 => \N__31084\,
            in3 => \N__17861\,
            lcout => \c0.n18558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1098_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22548\,
            in1 => \N__21895\,
            in2 => \_gnd_net_\,
            in3 => \N__22637\,
            lcout => \c0.n2839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_964_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17423\,
            in1 => \N__20611\,
            in2 => \N__20689\,
            in3 => \N__18789\,
            lcout => \c0.n12_adj_2492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_973_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21907\,
            in1 => \N__18679\,
            in2 => \_gnd_net_\,
            in3 => \N__21839\,
            lcout => \c0.n9058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_962_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28217\,
            in1 => \N__20668\,
            in2 => \_gnd_net_\,
            in3 => \N__19937\,
            lcout => \c0.n17476\,
            ltout => \c0.n17476_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_977_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25445\,
            in1 => \N__24884\,
            in2 => \N__17417\,
            in3 => \N__23773\,
            lcout => OPEN,
            ltout => \c0.n17478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_983_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__17414\,
            in2 => \N__17408\,
            in3 => \N__20178\,
            lcout => \c0.n9_adj_2507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i17_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__27122\,
            in1 => \N__24246\,
            in2 => \N__18662\,
            in3 => \N__31950\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i8_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24245\,
            in1 => \N__18680\,
            in2 => \N__31981\,
            in3 => \N__21653\,
            lcout => \c0.data_in_frame_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i22_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__26996\,
            in1 => \N__17500\,
            in2 => \N__24278\,
            in3 => \N__31951\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1076_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23794\,
            in1 => \N__22952\,
            in2 => \N__18938\,
            in3 => \N__22839\,
            lcout => \c0.n17629\,
            ltout => \c0.n17629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17519\,
            in3 => \N__20402\,
            lcout => \c0.n16_adj_2546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1020_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22670\,
            in1 => \N__22627\,
            in2 => \_gnd_net_\,
            in3 => \N__20099\,
            lcout => \c0.n9254\,
            ltout => \c0.n9254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1002_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20437\,
            in1 => \N__20481\,
            in2 => \N__17504\,
            in3 => \N__17499\,
            lcout => \c0.n17522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i20_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__21723\,
            in2 => \N__31980\,
            in3 => \N__37573\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_939_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24931\,
            in1 => \N__20144\,
            in2 => \_gnd_net_\,
            in3 => \N__17471\,
            lcout => \c0.n8886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i12_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24275\,
            in1 => \N__27643\,
            in2 => \N__17459\,
            in3 => \N__31808\,
            lcout => \c0.data_in_frame_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i50_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31806\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20186\,
            lcout => \c0.data_in_frame_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i65_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__28767\,
            in1 => \N__31804\,
            in2 => \N__23918\,
            in3 => \N__20261\,
            lcout => data_in_frame_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__30758\,
            in1 => \N__20798\,
            in2 => \N__17438\,
            in3 => \N__31031\,
            lcout => \c0.n6_adj_2506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i38_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24276\,
            in1 => \N__21905\,
            in2 => \N__27215\,
            in3 => \N__31809\,
            lcout => \c0.data_in_frame_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i49_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31805\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23777\,
            lcout => \c0.data_in_frame_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i42_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24277\,
            in1 => \N__24963\,
            in2 => \N__39899\,
            in3 => \N__31807\,
            lcout => data_in_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_913_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21773\,
            in1 => \N__22172\,
            in2 => \N__18743\,
            in3 => \N__22480\,
            lcout => \c0.n17467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3963_3_lut_4_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__34673\,
            in2 => \N__22102\,
            in3 => \N__28062\,
            lcout => \c0.n2607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3953_3_lut_4_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__34674\,
            in1 => \N__29563\,
            in2 => \N__28067\,
            in3 => \N__18767\,
            lcout => \c0.n2602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i6_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__33166\,
            in1 => \N__17549\,
            in2 => \N__33697\,
            in3 => \N__23866\,
            lcout => \c0.data_out_frame2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i28_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24259\,
            in1 => \N__27548\,
            in2 => \N__17537\,
            in3 => \N__31817\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i13_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__19963\,
            in1 => \N__37661\,
            in2 => \N__31923\,
            in3 => \N__24261\,
            lcout => \c0.data_in_frame_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i41_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24260\,
            in1 => \N__22098\,
            in2 => \N__21605\,
            in3 => \N__31816\,
            lcout => data_in_frame_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i46_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__29564\,
            in1 => \N__18768\,
            in2 => \N__31922\,
            in3 => \N__24262\,
            lcout => data_in_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_972_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__24556\,
            in1 => \N__17603\,
            in2 => \N__17597\,
            in3 => \N__17588\,
            lcout => \c0.n9_adj_2500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i64_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20033\,
            lcout => \c0.data_in_frame_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i48_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24264\,
            in1 => \N__28315\,
            in2 => \N__36923\,
            in3 => \N__31838\,
            lcout => data_in_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i52_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22280\,
            lcout => \c0.data_in_frame_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i56_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__36962\,
            in2 => \N__25107\,
            in3 => \N__31840\,
            lcout => \c0.data_in_frame_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i27_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__37523\,
            in2 => \N__31926\,
            in3 => \N__24266\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i63_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22736\,
            in2 => \_gnd_net_\,
            in3 => \N__31839\,
            lcout => \c0.data_in_frame_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i25_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__22580\,
            in1 => \N__27839\,
            in2 => \N__31925\,
            in3 => \N__24265\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_982_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22241\,
            in1 => \N__22190\,
            in2 => \N__17558\,
            in3 => \N__17645\,
            lcout => OPEN,
            ltout => \c0.n17325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_984_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17666\,
            in1 => \N__24806\,
            in2 => \N__17657\,
            in3 => \N__18953\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_970_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22767\,
            in1 => \N__20306\,
            in2 => \N__18907\,
            in3 => \N__22379\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__18863\,
            in1 => \N__19997\,
            in2 => \N__17654\,
            in3 => \N__17651\,
            lcout => \c0.n11_adj_2460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15860_3_lut_4_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__23198\,
            in1 => \N__33522\,
            in2 => \N__33379\,
            in3 => \N__33242\,
            lcout => \c0.n9605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1086_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33241\,
            in1 => \N__33363\,
            in2 => \N__33529\,
            in3 => \N__23199\,
            lcout => \c0.n9900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i107_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35828\,
            in2 => \N__17792\,
            in3 => \N__32764\,
            lcout => data_out_frame2_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18540_bdd_4_lut_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__30963\,
            in1 => \N__17758\,
            in2 => \N__19100\,
            in3 => \N__23627\,
            lcout => \c0.n17806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i57_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24575\,
            lcout => data_in_frame_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i150_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17615\,
            in2 => \N__32825\,
            in3 => \N__35098\,
            lcout => data_out_frame2_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18492_bdd_4_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__17788\,
            in1 => \N__30962\,
            in2 => \N__19013\,
            in3 => \N__17780\,
            lcout => \c0.n17827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i102_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17759\,
            in2 => \N__32824\,
            in3 => \N__35097\,
            lcout => data_out_frame2_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_853_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25062\,
            in1 => \N__23050\,
            in2 => \_gnd_net_\,
            in3 => \N__19058\,
            lcout => \c0.n9043\,
            ltout => \c0.n9043_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1120_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22893\,
            in1 => \N__28316\,
            in2 => \N__17750\,
            in3 => \N__25073\,
            lcout => \c0.n17562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i119_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36042\,
            in1 => \N__17743\,
            in2 => \_gnd_net_\,
            in3 => \N__32620\,
            lcout => data_out_frame2_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i41_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__35951\,
            in2 => \_gnd_net_\,
            in3 => \N__18310\,
            lcout => data_out_frame2_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i87_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36044\,
            in1 => \N__17725\,
            in2 => \_gnd_net_\,
            in3 => \N__32623\,
            lcout => data_out_frame2_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i89_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32619\,
            in1 => \N__34886\,
            in2 => \_gnd_net_\,
            in3 => \N__17704\,
            lcout => data_out_frame2_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i55_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36043\,
            in1 => \N__17680\,
            in2 => \_gnd_net_\,
            in3 => \N__32621\,
            lcout => data_out_frame2_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i63_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32618\,
            in1 => \N__35534\,
            in2 => \_gnd_net_\,
            in3 => \N__17920\,
            lcout => data_out_frame2_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i70_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17906\,
            in1 => \N__35093\,
            in2 => \_gnd_net_\,
            in3 => \N__32622\,
            lcout => data_out_frame2_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i122_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32616\,
            in1 => \N__34829\,
            in2 => \_gnd_net_\,
            in3 => \N__17893\,
            lcout => data_out_frame2_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i95_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32757\,
            in1 => \N__35533\,
            in2 => \_gnd_net_\,
            in3 => \N__17875\,
            lcout => data_out_frame2_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i127_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35532\,
            in1 => \N__17860\,
            in2 => \_gnd_net_\,
            in3 => \N__32760\,
            lcout => data_out_frame2_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i43_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32754\,
            in1 => \N__35821\,
            in2 => \_gnd_net_\,
            in3 => \N__17842\,
            lcout => data_out_frame2_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i123_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34764\,
            in1 => \N__17824\,
            in2 => \_gnd_net_\,
            in3 => \N__32759\,
            lcout => data_out_frame2_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i71_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32755\,
            in1 => \N__35042\,
            in2 => \_gnd_net_\,
            in3 => \N__18025\,
            lcout => data_out_frame2_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i121_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34885\,
            in1 => \N__17806\,
            in2 => \_gnd_net_\,
            in3 => \N__32758\,
            lcout => data_out_frame2_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i83_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32756\,
            in1 => \N__35305\,
            in2 => \_gnd_net_\,
            in3 => \N__18250\,
            lcout => data_out_frame2_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18564_bdd_4_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__23378\,
            in1 => \N__31032\,
            in2 => \N__18026\,
            in3 => \N__18014\,
            lcout => \c0.n17794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i146_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32626\,
            in1 => \N__34165\,
            in2 => \_gnd_net_\,
            in3 => \N__18283\,
            lcout => data_out_frame2_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i130_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34164\,
            in1 => \N__17998\,
            in2 => \_gnd_net_\,
            in3 => \N__32629\,
            lcout => data_out_frame2_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i137_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32625\,
            in1 => \N__34880\,
            in2 => \_gnd_net_\,
            in3 => \N__18064\,
            lcout => data_out_frame2_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i138_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34825\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \N__32630\,
            lcout => data_out_frame2_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i129_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32624\,
            in1 => \N__34220\,
            in2 => \_gnd_net_\,
            in3 => \N__18046\,
            lcout => data_out_frame2_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i145_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34219\,
            in1 => \N__17963\,
            in2 => \_gnd_net_\,
            in3 => \N__32631\,
            lcout => data_out_frame2_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i84_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32627\,
            in1 => \N__35260\,
            in2 => \_gnd_net_\,
            in3 => \N__17951\,
            lcout => data_out_frame2_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i117_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__17939\,
            in2 => \_gnd_net_\,
            in3 => \N__32628\,
            lcout => data_out_frame2_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__18161\,
            in1 => \N__30768\,
            in2 => \N__18155\,
            in3 => \N__31122\,
            lcout => \c0.n6_adj_2496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i92_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35706\,
            in1 => \N__18121\,
            in2 => \_gnd_net_\,
            in3 => \N__32723\,
            lcout => data_out_frame2_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_954_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20461\,
            in1 => \N__18107\,
            in2 => \_gnd_net_\,
            in3 => \N__18098\,
            lcout => \c0.n8890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i64_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45291\,
            in1 => \N__29800\,
            in2 => \_gnd_net_\,
            in3 => \N__32140\,
            lcout => data_in_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_993_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30767\,
            in2 => \_gnd_net_\,
            in3 => \N__31118\,
            lcout => \c0.n134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i81_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35407\,
            in1 => \N__18080\,
            in2 => \_gnd_net_\,
            in3 => \N__32722\,
            lcout => data_out_frame2_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i53_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32721\,
            in1 => \N__36151\,
            in2 => \_gnd_net_\,
            in3 => \N__30214\,
            lcout => data_out_frame2_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__20327\,
            in1 => \N__19192\,
            in2 => \N__31142\,
            in3 => \N__30769\,
            lcout => \c0.n6_adj_2464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18600_bdd_4_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__31132\,
            in1 => \N__18068\,
            in2 => \N__18050\,
            in3 => \N__18032\,
            lcout => \c0.n18603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__30735\,
            in1 => \_gnd_net_\,
            in2 => \N__19328\,
            in3 => \N__19139\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__31134\,
            in1 => \N__18314\,
            in2 => \N__18296\,
            in3 => \N__30737\,
            lcout => \c0.n6_adj_2436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i151_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35029\,
            in1 => \N__18377\,
            in2 => \_gnd_net_\,
            in3 => \N__32810\,
            lcout => data_out_frame2_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16001_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__31133\,
            in1 => \N__18284\,
            in2 => \N__21032\,
            in3 => \N__30736\,
            lcout => \c0.n18468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i42_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35886\,
            in1 => \N__18263\,
            in2 => \_gnd_net_\,
            in3 => \N__32811\,
            lcout => data_out_frame2_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16031_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__31131\,
            in1 => \N__18251\,
            in2 => \N__18236\,
            in3 => \N__30734\,
            lcout => \c0.n18504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i97_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34213\,
            in1 => \N__18212\,
            in2 => \_gnd_net_\,
            in3 => \N__32812\,
            lcout => data_out_frame2_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15960_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18200\,
            in1 => \N__26675\,
            in2 => \N__18815\,
            in3 => \N__26827\,
            lcout => OPEN,
            ltout => \c0.n18408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18408_bdd_4_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__26676\,
            in1 => \N__18191\,
            in2 => \N__18176\,
            in3 => \N__18173\,
            lcout => OPEN,
            ltout => \c0.n18411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__18359\,
            in1 => \N__26677\,
            in2 => \N__18380\,
            in3 => \N__26508\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50333\,
            ce => \N__26377\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16071_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__31140\,
            in1 => \N__18376\,
            in2 => \N__21101\,
            in3 => \N__30733\,
            lcout => OPEN,
            ltout => \c0.n18552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18552_bdd_4_lut_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__19555\,
            in1 => \N__19295\,
            in2 => \N__18365\,
            in3 => \N__31141\,
            lcout => OPEN,
            ltout => \c0.n18555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26826\,
            in1 => \N__20636\,
            in2 => \N__18362\,
            in3 => \N__26929\,
            lcout => \c0.n22_adj_2521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i4_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__21411\,
            in1 => \N__18570\,
            in2 => \N__18353\,
            in3 => \N__18444\,
            lcout => \r_Clock_Count_4_adj_2630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i3_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__18441\,
            in1 => \N__21413\,
            in2 => \N__18344\,
            in3 => \N__18553\,
            lcout => \r_Clock_Count_3_adj_2631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i2_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__21412\,
            in1 => \N__18590\,
            in2 => \N__18335\,
            in3 => \N__18443\,
            lcout => \r_Clock_Count_2_adj_2632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21505\,
            in1 => \N__21347\,
            in2 => \N__21294\,
            in3 => \N__21409\,
            lcout => \c0.tx2.n7727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__21410\,
            in1 => \N__18442\,
            in2 => \N__18323\,
            in3 => \N__18604\,
            lcout => \r_Clock_Count_0_adj_2634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4_4_lut_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18603\,
            in1 => \N__18588\,
            in2 => \N__18572\,
            in3 => \N__18552\,
            lcout => OPEN,
            ltout => \c0.tx2.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5_3_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__18537\,
            in1 => \_gnd_net_\,
            in2 => \N__18521\,
            in3 => \N__18396\,
            lcout => \c0.tx2.n16452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11588211_i1_3_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25889\,
            in1 => \N__19568\,
            in2 => \_gnd_net_\,
            in3 => \N__19490\,
            lcout => \c0.tx2.o_Tx_Serial_N_2354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15730_2_lut_3_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25884\,
            in1 => \N__26181\,
            in2 => \_gnd_net_\,
            in3 => \N__21465\,
            lcout => \c0.tx2.n17990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_4_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18516\,
            in1 => \N__18498\,
            in2 => \N__18482\,
            in3 => \N__18461\,
            lcout => \c0.tx2.r_SM_Main_2_N_2323_1\,
            ltout => \c0.tx2.r_SM_Main_2_N_2323_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__21284\,
            in1 => \N__21342\,
            in2 => \N__18455\,
            in3 => \N__21425\,
            lcout => \c0.tx2.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21343\,
            in1 => \N__21466\,
            in2 => \N__21433\,
            in3 => \N__21283\,
            lcout => \r_SM_Main_2_adj_2628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i1_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__18452\,
            in1 => \N__21421\,
            in2 => \N__18401\,
            in3 => \N__18446\,
            lcout => \r_Clock_Count_1_adj_2633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i9901_3_lut_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__18614\,
            in1 => \N__21279\,
            in2 => \_gnd_net_\,
            in3 => \N__21341\,
            lcout => OPEN,
            ltout => \c0.tx2.n12306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21414\,
            in2 => \N__18608\,
            in3 => \N__21135\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \N__33378\,
            in1 => \N__33515\,
            in2 => \N__33698\,
            in3 => \N__33229\,
            lcout => \c0.FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50254\,
            ce => 'H',
            sr => \N__33413\
        );

    \c0.i3945_3_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39932\,
            in1 => \N__22009\,
            in2 => \_gnd_net_\,
            in3 => \N__24217\,
            lcout => n2598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_859_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47648\,
            in2 => \_gnd_net_\,
            in3 => \N__41807\,
            lcout => \c0.n8600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_894_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21552\,
            in2 => \_gnd_net_\,
            in3 => \N__22046\,
            lcout => \c0.n17424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_986_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19753\,
            in2 => \_gnd_net_\,
            in3 => \N__18640\,
            lcout => \c0.n17614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_100_i4_2_lut_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__39241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39313\,
            lcout => n4_adj_2582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_102_i4_2_lut_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__39314\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39240\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i62_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20729\,
            in1 => \N__45482\,
            in2 => \_gnd_net_\,
            in3 => \N__36210\,
            lcout => data_in_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_965_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19807\,
            in1 => \N__18686\,
            in2 => \N__29133\,
            in3 => \N__20528\,
            lcout => \c0.n9334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i6_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__37616\,
            in1 => \N__24270\,
            in2 => \N__21868\,
            in3 => \N__31876\,
            lcout => \c0.data_in_frame_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_961_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18678\,
            in1 => \N__18731\,
            in2 => \_gnd_net_\,
            in3 => \N__18657\,
            lcout => \c0.n9349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i15_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__27797\,
            in1 => \N__24269\,
            in2 => \N__19904\,
            in3 => \N__31875\,
            lcout => \c0.data_in_frame_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i32_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24268\,
            in1 => \N__18641\,
            in2 => \N__31943\,
            in3 => \N__23954\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1026_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18638\,
            lcout => \c0.n17553\,
            ltout => \c0.n17553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_994_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22134\,
            in1 => \N__29122\,
            in2 => \N__18644\,
            in3 => \N__19898\,
            lcout => \c0.n8658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1033_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21685\,
            in1 => \N__19754\,
            in2 => \N__21764\,
            in3 => \N__18639\,
            lcout => \c0.n25_adj_2491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_933_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22485\,
            in2 => \_gnd_net_\,
            in3 => \N__22669\,
            lcout => \c0.n17406\,
            ltout => \c0.n17406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_936_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18855\,
            in1 => \N__22591\,
            in2 => \N__18617\,
            in3 => \N__21837\,
            lcout => \c0.n17656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i2_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24240\,
            in1 => \N__29126\,
            in2 => \N__31941\,
            in3 => \N__27077\,
            lcout => \c0.data_in_frame_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i1_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__23984\,
            in1 => \N__24242\,
            in2 => \N__18883\,
            in3 => \N__31870\,
            lcout => \c0.data_in_frame_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_846_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18876\,
            in2 => \_gnd_net_\,
            in3 => \N__18769\,
            lcout => \c0.n23_adj_2426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i21_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__27325\,
            in1 => \N__24243\,
            in2 => \N__18739\,
            in3 => \N__31871\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i35_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__24241\,
            in1 => \N__29858\,
            in2 => \N__31942\,
            in3 => \N__21754\,
            lcout => \c0.data_in_frame_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i14_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__18705\,
            in1 => \N__36259\,
            in2 => \N__31850\,
            in3 => \N__24213\,
            lcout => \c0.data_in_frame_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_942_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__34660\,
            in1 => \N__34452\,
            in2 => \_gnd_net_\,
            in3 => \N__31712\,
            lcout => n9419,
            ltout => \n9419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i67_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__31713\,
            in1 => \N__33941\,
            in2 => \N__18689\,
            in3 => \N__22953\,
            lcout => data_in_frame_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i47_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24212\,
            in1 => \N__31271\,
            in2 => \N__24677\,
            in3 => \N__31723\,
            lcout => data_in_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i23_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__22484\,
            in1 => \N__27718\,
            in2 => \N__31851\,
            in3 => \N__24214\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1087_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29056\,
            in1 => \N__18793\,
            in2 => \N__20570\,
            in3 => \N__21722\,
            lcout => \c0.n17569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i39_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__28384\,
            in1 => \N__22628\,
            in2 => \N__31852\,
            in3 => \N__24215\,
            lcout => \c0.data_in_frame_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12308_3_lut_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33508\,
            in1 => \N__25133\,
            in2 => \_gnd_net_\,
            in3 => \N__23263\,
            lcout => \c0.n81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i70_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__31790\,
            in1 => \N__20728\,
            in2 => \N__20276\,
            in3 => \N__19053\,
            lcout => data_in_frame_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i61_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27473\,
            in2 => \_gnd_net_\,
            in3 => \N__31796\,
            lcout => \c0.data_in_frame_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i30_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__25385\,
            in1 => \N__27182\,
            in2 => \N__31920\,
            in3 => \N__24267\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i71_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__28438\,
            in1 => \N__31791\,
            in2 => \N__38768\,
            in3 => \N__20273\,
            lcout => data_in_frame_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i69_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__31789\,
            in1 => \N__38384\,
            in2 => \N__20275\,
            in3 => \N__25052\,
            lcout => data_in_frame_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1017_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__33387\,
            in1 => \N__33217\,
            in2 => \N__32826\,
            in3 => \N__23859\,
            lcout => n1396,
            ltout => \n1396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i88_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18839\,
            in3 => \N__23156\,
            lcout => \c0.data_in_frame_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i53_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18908\,
            in2 => \_gnd_net_\,
            in3 => \N__31795\,
            lcout => \c0.data_in_frame_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3927_3_lut_4_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__33764\,
            in1 => \N__34675\,
            in2 => \N__28631\,
            in3 => \N__28058\,
            lcout => n2589,
            ltout => \n2589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_899_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25502\,
            in1 => \N__24782\,
            in2 => \N__18836\,
            in3 => \N__18903\,
            lcout => \c0.n23_adj_2462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i74_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28826\,
            in2 => \_gnd_net_\,
            in3 => \N__31822\,
            lcout => \c0.data_in_frame_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i54_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27947\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i59_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18833\,
            in2 => \_gnd_net_\,
            in3 => \N__31821\,
            lcout => \c0.data_in_frame_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i62_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__31819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22352\,
            lcout => \c0.data_in_frame_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i51_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24908\,
            in2 => \_gnd_net_\,
            in3 => \N__31820\,
            lcout => \c0.data_in_frame_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18558_bdd_4_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__30991\,
            in2 => \N__20759\,
            in3 => \N__18827\,
            lcout => \c0.n17797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1095_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28477\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22832\,
            lcout => \c0.n9028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_979_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__18980\,
            in1 => \N__25232\,
            in2 => \N__18965\,
            in3 => \N__27946\,
            lcout => \c0.n10_adj_2505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1092_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28340\,
            in1 => \N__25345\,
            in2 => \_gnd_net_\,
            in3 => \N__20136\,
            lcout => \c0.n8061\,
            ltout => \c0.n8061_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1099_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18947\,
            in1 => \N__28621\,
            in2 => \N__18941\,
            in3 => \N__20579\,
            lcout => \c0.n17538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3939_3_lut_4_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__18937\,
            in1 => \N__34672\,
            in2 => \N__27437\,
            in3 => \N__28052\,
            lcout => n2595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_896_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29084\,
            in2 => \_gnd_net_\,
            in3 => \N__18884\,
            lcout => \c0.n9039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_967_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28432\,
            in1 => \N__28476\,
            in2 => \_gnd_net_\,
            in3 => \N__25461\,
            lcout => \c0.n9279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i164_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24315\,
            in1 => \N__32985\,
            in2 => \N__36557\,
            in3 => \N__25207\,
            lcout => \c0.data_out_frame2_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__32771\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_903_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19996\,
            in1 => \N__21608\,
            in2 => \_gnd_net_\,
            in3 => \N__18862\,
            lcout => \c0.n9151\,
            ltout => \c0.n9151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_850_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19031\,
            in1 => \N__25106\,
            in2 => \N__19064\,
            in3 => \N__22805\,
            lcout => \c0.n17588\,
            ltout => \c0.n17588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i156_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32984\,
            in2 => \N__19061\,
            in3 => \N__32213\,
            lcout => \c0.data_out_frame2_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__32771\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_849_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28433\,
            in2 => \_gnd_net_\,
            in3 => \N__19057\,
            lcout => \c0.n6_adj_2429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i166_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__36556\,
            in1 => \N__32256\,
            in2 => \_gnd_net_\,
            in3 => \N__25175\,
            lcout => \c0.data_out_frame2_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__32771\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i157_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28808\,
            in1 => \N__29197\,
            in2 => \_gnd_net_\,
            in3 => \N__24316\,
            lcout => \c0.data_out_frame2_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50292\,
            ce => \N__32771\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i99_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34108\,
            in1 => \N__32607\,
            in2 => \_gnd_net_\,
            in3 => \N__19012\,
            lcout => data_out_frame2_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i120_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32601\,
            in1 => \N__36003\,
            in2 => \_gnd_net_\,
            in3 => \N__19444\,
            lcout => data_out_frame2_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i106_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18994\,
            in1 => \N__32605\,
            in2 => \_gnd_net_\,
            in3 => \N__35888\,
            lcout => data_out_frame2_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i56_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32603\,
            in1 => \N__36004\,
            in2 => \_gnd_net_\,
            in3 => \N__20341\,
            lcout => data_out_frame2_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i126_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__32606\,
            in2 => \_gnd_net_\,
            in3 => \N__23641\,
            lcout => data_out_frame2_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i128_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32602\,
            in1 => \N__35467\,
            in2 => \_gnd_net_\,
            in3 => \N__19429\,
            lcout => data_out_frame2_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i8_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__33149\,
            in1 => \N__23464\,
            in2 => \N__33677\,
            in3 => \N__23877\,
            lcout => \c0.data_out_frame2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i98_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32604\,
            in1 => \N__34166\,
            in2 => \_gnd_net_\,
            in3 => \N__19153\,
            lcout => data_out_frame2_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i57_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34884\,
            in1 => \N__19135\,
            in2 => \_gnd_net_\,
            in3 => \N__32762\,
            lcout => data_out_frame2_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1038_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33345\,
            in1 => \N__33230\,
            in2 => \N__33530\,
            in3 => \N__23206\,
            lcout => n9606,
            ltout => \n9606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i86_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36104\,
            in2 => \N__19121\,
            in3 => \N__19117\,
            lcout => data_out_frame2_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i110_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32598\,
            in1 => \N__36408\,
            in2 => \_gnd_net_\,
            in3 => \N__19096\,
            lcout => data_out_frame2_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i73_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35950\,
            in1 => \N__19078\,
            in2 => \_gnd_net_\,
            in3 => \N__32763\,
            lcout => data_out_frame2_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i141_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32599\,
            in1 => \_gnd_net_\,
            in2 => \N__35663\,
            in3 => \N__26200\,
            lcout => data_out_frame2_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i108_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35774\,
            in1 => \N__23329\,
            in2 => \_gnd_net_\,
            in3 => \N__32761\,
            lcout => data_out_frame2_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i74_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32600\,
            in1 => \N__35887\,
            in2 => \_gnd_net_\,
            in3 => \N__19267\,
            lcout => data_out_frame2_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i50_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19228\,
            in1 => \N__32614\,
            in2 => \_gnd_net_\,
            in3 => \N__35355\,
            lcout => data_out_frame2_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i139_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32608\,
            in1 => \N__34757\,
            in2 => \_gnd_net_\,
            in3 => \N__19207\,
            lcout => data_out_frame2_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i48_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36308\,
            in1 => \N__32613\,
            in2 => \_gnd_net_\,
            in3 => \N__19193\,
            lcout => data_out_frame2_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i67_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32611\,
            in1 => \N__34101\,
            in2 => \_gnd_net_\,
            in3 => \N__19372\,
            lcout => data_out_frame2_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i112_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36307\,
            in1 => \N__32612\,
            in2 => \_gnd_net_\,
            in3 => \N__19402\,
            lcout => data_out_frame2_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i54_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32610\,
            in1 => \N__36100\,
            in2 => \_gnd_net_\,
            in3 => \N__19174\,
            lcout => data_out_frame2_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i60_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35715\,
            in1 => \N__32615\,
            in2 => \_gnd_net_\,
            in3 => \N__19717\,
            lcout => data_out_frame2_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i49_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32609\,
            in1 => \N__35408\,
            in2 => \_gnd_net_\,
            in3 => \N__19324\,
            lcout => data_out_frame2_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i58_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32715\,
            in1 => \N__34824\,
            in2 => \_gnd_net_\,
            in3 => \N__19309\,
            lcout => data_out_frame2_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i135_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35040\,
            in1 => \N__19291\,
            in2 => \_gnd_net_\,
            in3 => \N__32718\,
            lcout => data_out_frame2_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16105_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__19276\,
            in1 => \N__20923\,
            in2 => \N__31130\,
            in3 => \N__30759\,
            lcout => \c0.n18588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i96_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35460\,
            in1 => \N__19277\,
            in2 => \_gnd_net_\,
            in3 => \N__32720\,
            lcout => data_out_frame2_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i76_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32716\,
            in1 => \_gnd_net_\,
            in2 => \N__23510\,
            in3 => \N__35770\,
            lcout => data_out_frame2_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i66_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34160\,
            in1 => \N__19252\,
            in2 => \_gnd_net_\,
            in3 => \N__32719\,
            lcout => data_out_frame2_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18480_bdd_4_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__31100\,
            in1 => \N__19268\,
            in2 => \N__19253\,
            in3 => \N__23288\,
            lcout => \c0.n17833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i132_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35210\,
            in1 => \N__25999\,
            in2 => \_gnd_net_\,
            in3 => \N__32717\,
            lcout => data_out_frame2_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i75_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35809\,
            in1 => \N__19388\,
            in2 => \_gnd_net_\,
            in3 => \N__32800\,
            lcout => data_out_frame2_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i153_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32798\,
            in1 => \N__19474\,
            in2 => \_gnd_net_\,
            in3 => \N__25831\,
            lcout => data_out_frame2_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39778\,
            in2 => \_gnd_net_\,
            in3 => \N__30182\,
            lcout => \c0.rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i152_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32797\,
            in1 => \N__34956\,
            in2 => \_gnd_net_\,
            in3 => \N__21233\,
            lcout => data_out_frame2_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i104_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19415\,
            in1 => \N__34955\,
            in2 => \_gnd_net_\,
            in3 => \N__32799\,
            lcout => data_out_frame2_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__26834\,
            in1 => \N__19460\,
            in2 => \N__20879\,
            in3 => \N__26905\,
            lcout => \c0.n22_adj_2510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16096_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__30754\,
            in2 => \N__31143\,
            in3 => \N__19430\,
            lcout => OPEN,
            ltout => \c0.n18582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18582_bdd_4_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31128\,
            in1 => \N__19414\,
            in2 => \N__19406\,
            in3 => \N__19403\,
            lcout => \c0.n17788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18504_bdd_4_lut_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__19387\,
            in1 => \N__31129\,
            in2 => \N__19376\,
            in3 => \N__19358\,
            lcout => \c0.n17824\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__26118\,
            in1 => \N__26051\,
            in2 => \N__26180\,
            in3 => \N__19340\,
            lcout => OPEN,
            ltout => \c0.tx2.n18612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18612_bdd_4_lut_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__19592\,
            in1 => \N__19580\,
            in2 => \N__19571\,
            in3 => \N__26168\,
            lcout => \c0.tx2.n18615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_16115_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__21005\,
            in1 => \N__19562\,
            in2 => \N__26129\,
            in3 => \N__26167\,
            lcout => \c0.tx2.n18450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__26119\,
            in1 => \N__25935\,
            in2 => \_gnd_net_\,
            in3 => \N__25905\,
            lcout => \r_Bit_Index_0_adj_2637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__25906\,
            in1 => \N__26169\,
            in2 => \N__25942\,
            in3 => \N__26120\,
            lcout => \r_Bit_Index_1_adj_2636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i143_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19556\,
            in1 => \N__35523\,
            in2 => \_gnd_net_\,
            in3 => \N__32809\,
            lcout => data_out_frame2_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__30773\,
            in1 => \N__19703\,
            in2 => \N__19730\,
            in3 => \N__31043\,
            lcout => \c0.n6_adj_2432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20981\,
            in1 => \N__19544\,
            in2 => \_gnd_net_\,
            in3 => \N__30771\,
            lcout => OPEN,
            ltout => \c0.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_15987_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__31035\,
            in1 => \N__19526\,
            in2 => \N__19514\,
            in3 => \N__26833\,
            lcout => \c0.n18444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18450_bdd_4_lut_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__19511\,
            in1 => \N__26170\,
            in2 => \N__26432\,
            in3 => \N__19496\,
            lcout => \c0.tx2.n18453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i44_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19729\,
            in1 => \N__35769\,
            in2 => \_gnd_net_\,
            in3 => \N__32813\,
            lcout => data_out_frame2_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19718\,
            in1 => \N__20777\,
            in2 => \_gnd_net_\,
            in3 => \N__30772\,
            lcout => \c0.n5_adj_2509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1100_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__26519\,
            in2 => \_gnd_net_\,
            in3 => \N__26785\,
            lcout => OPEN,
            ltout => \c0.n18_adj_2544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1102_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19697\,
            in1 => \N__19673\,
            in2 => \N__19649\,
            in3 => \N__19646\,
            lcout => \c0.n19_adj_2540\,
            ltout => \c0.n19_adj_2540_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15867_2_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19622\,
            in3 => \N__19822\,
            lcout => \c0.tx2_transmit_N_2287\,
            ltout => \c0.tx2_transmit_N_2287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_3602_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33251\,
            in1 => \N__33322\,
            in2 => \N__19607\,
            in3 => \N__33518\,
            lcout => \c0.r_SM_Main_2_N_2326_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50365\,
            ce => 'H',
            sr => \N__33633\
        );

    \c0.i3_3_lut_adj_1105_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__33517\,
            in1 => \N__33249\,
            in2 => \_gnd_net_\,
            in3 => \N__33320\,
            lcout => OPEN,
            ltout => \c0.n67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1071_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__19823\,
            in1 => \N__19604\,
            in2 => \N__19595\,
            in3 => \N__32643\,
            lcout => \c0.n4_adj_2480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11145_2_lut_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21500\,
            in2 => \_gnd_net_\,
            in3 => \N__21523\,
            lcout => \c0.n13530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15907_2_lut_3_lut_LC_3_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__33250\,
            in1 => \N__33321\,
            in2 => \_gnd_net_\,
            in3 => \N__33516\,
            lcout => \c0.n142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1018_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20290\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25273\,
            lcout => \c0.n8062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_938_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19814\,
            in2 => \_gnd_net_\,
            in3 => \N__28716\,
            lcout => \c0.n17529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_847_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29134\,
            in1 => \N__19922\,
            in2 => \N__20135\,
            in3 => \N__19796\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_848_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \N__19787\,
            in3 => \N__20289\,
            lcout => \c0.n9324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1050_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21684\,
            in1 => \N__20527\,
            in2 => \_gnd_net_\,
            in3 => \N__19748\,
            lcout => \c0.n17442\,
            ltout => \c0.n17442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_948_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29089\,
            in1 => \N__19775\,
            in2 => \N__19766\,
            in3 => \N__19763\,
            lcout => \c0.n8674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i10_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__31382\,
            in2 => \N__28723\,
            in3 => \N__31937\,
            lcout => data_in_frame_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i33_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__19749\,
            in1 => \N__27865\,
            in2 => \N__31978\,
            in3 => \N__24257\,
            lcout => \c0.data_in_frame_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1079_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28714\,
            in1 => \N__20093\,
            in2 => \N__22041\,
            in3 => \N__19851\,
            lcout => \c0.n8874\,
            ltout => \c0.n8874_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_963_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19902\,
            in1 => \N__19967\,
            in2 => \N__19940\,
            in3 => \N__19936\,
            lcout => \c0.n9368\,
            ltout => \c0.n9368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1093_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21906\,
            in1 => \N__21606\,
            in2 => \N__19925\,
            in3 => \N__19918\,
            lcout => \c0.n12_adj_2542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_3_lut_4_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22595\,
            in1 => \N__22635\,
            in2 => \N__28261\,
            in3 => \N__22542\,
            lcout => \c0.n9306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1031_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22138\,
            in2 => \_gnd_net_\,
            in3 => \N__19903\,
            lcout => \c0.n17632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_865_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20094\,
            in1 => \N__22033\,
            in2 => \_gnd_net_\,
            in3 => \N__28715\,
            lcout => \c0.n17485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i40_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__22543\,
            in1 => \N__24258\,
            in2 => \N__27245\,
            in3 => \N__31877\,
            lcout => \c0.data_in_frame_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i26_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24237\,
            in1 => \N__27689\,
            in2 => \N__19858\,
            in3 => \N__31994\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_884_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19832\,
            in1 => \N__21553\,
            in2 => \N__24764\,
            in3 => \N__22183\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24838\,
            in1 => \N__22973\,
            in2 => \N__20189\,
            in3 => \N__20182\,
            lcout => OPEN,
            ltout => \c0.n24_adj_2454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22358\,
            in1 => \N__20159\,
            in2 => \N__20147\,
            in3 => \N__20003\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i73_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29351\,
            in2 => \_gnd_net_\,
            in3 => \N__31993\,
            lcout => \c0.data_in_frame_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i44_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24238\,
            in1 => \N__20122\,
            in2 => \N__23698\,
            in3 => \N__31992\,
            lcout => data_in_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i24_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20098\,
            in1 => \N__27284\,
            in2 => \N__31997\,
            in3 => \N__24239\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3917_3_lut_4_lut_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__20075\,
            in1 => \N__34659\,
            in2 => \N__32161\,
            in3 => \N__28045\,
            lcout => n2584,
            ltout => \n2584_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_901_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__20021\,
            in1 => \N__22783\,
            in2 => \N__20006\,
            in3 => \N__22273\,
            lcout => \c0.n21_adj_2465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i68_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__25555\,
            in1 => \N__31798\,
            in2 => \N__29747\,
            in3 => \N__20265\,
            lcout => data_in_frame_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i66_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__31797\,
            in1 => \N__37042\,
            in2 => \N__20274\,
            in3 => \N__22925\,
            lcout => data_in_frame_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i72_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__20375\,
            in1 => \N__31799\,
            in2 => \N__29807\,
            in3 => \N__20266\,
            lcout => data_in_frame_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i16_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__25432\,
            in1 => \N__27041\,
            in2 => \N__31921\,
            in3 => \N__24216\,
            lcout => \c0.data_in_frame_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i55_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22375\,
            in2 => \_gnd_net_\,
            in3 => \N__31803\,
            lcout => \c0.data_in_frame_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_909_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__27942\,
            in2 => \N__20237\,
            in3 => \N__22201\,
            lcout => \c0.n18_adj_2468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i60_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22202\,
            in1 => \_gnd_net_\,
            in2 => \N__31924\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_910_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__22345\,
            in1 => \N__23753\,
            in2 => \N__20225\,
            in3 => \N__20312\,
            lcout => OPEN,
            ltout => \c0.n26_adj_2469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_916_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20207\,
            in1 => \N__22718\,
            in2 => \N__20201\,
            in3 => \N__20198\,
            lcout => \c0.n1_adj_2443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i87_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31824\,
            in2 => \_gnd_net_\,
            in3 => \N__29450\,
            lcout => data_in_frame_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i85_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__31829\,
            in1 => \N__28658\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i80_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31823\,
            in2 => \_gnd_net_\,
            in3 => \N__25220\,
            lcout => \c0.data_in_frame_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i79_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__31828\,
            in1 => \N__28894\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => data_in_frame_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i9_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24251\,
            in1 => \N__24014\,
            in2 => \N__22668\,
            in3 => \N__31849\,
            lcout => \c0.data_in_frame_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30674\,
            in1 => \N__32285\,
            in2 => \_gnd_net_\,
            in3 => \N__20345\,
            lcout => \c0.n5_adj_2501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i34_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24250\,
            in1 => \N__21683\,
            in2 => \N__38513\,
            in3 => \N__31848\,
            lcout => \c0.data_in_frame_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_887_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24523\,
            in1 => \_gnd_net_\,
            in2 => \N__20599\,
            in3 => \N__22310\,
            lcout => \c0.n17534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i76_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31847\,
            lcout => \c0.data_in_frame_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i31_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__29088\,
            in1 => \N__28190\,
            in2 => \N__31927\,
            in3 => \N__24252\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_978_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28565\,
            in1 => \N__25270\,
            in2 => \_gnd_net_\,
            in3 => \N__20305\,
            lcout => \c0.n17591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i37_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__27371\,
            in1 => \N__21829\,
            in2 => \N__31928\,
            in3 => \N__24253\,
            lcout => \c0.data_in_frame_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1045_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20491\,
            in1 => \N__20621\,
            in2 => \N__25272\,
            in3 => \N__24995\,
            lcout => \c0.n17470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_842_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22706\,
            in2 => \_gnd_net_\,
            in3 => \N__20376\,
            lcout => n9148,
            ltout => \n9148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25021\,
            in1 => \N__21929\,
            in2 => \N__20573\,
            in3 => \N__25582\,
            lcout => n17585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i45_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__24255\,
            in1 => \N__25263\,
            in2 => \N__27407\,
            in3 => \N__31892\,
            lcout => data_in_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1111_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20566\,
            in1 => \N__20513\,
            in2 => \N__25271\,
            in3 => \N__20537\,
            lcout => \c0.n17605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i19_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__24383\,
            in2 => \N__20523\,
            in3 => \N__31893\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1036_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20492\,
            in1 => \N__20462\,
            in2 => \_gnd_net_\,
            in3 => \N__20441\,
            lcout => \c0.n8751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i77_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31219\,
            in1 => \_gnd_net_\,
            in2 => \N__36470\,
            in3 => \N__32678\,
            lcout => data_out_frame2_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1127_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23024\,
            in1 => \N__20401\,
            in2 => \N__20381\,
            in3 => \N__20735\,
            lcout => \c0.n17647\,
            ltout => \c0.n17647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_854_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28530\,
            in2 => \N__20738\,
            in3 => \N__24416\,
            lcout => \c0.n17648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1125_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24693\,
            in1 => \N__20648\,
            in2 => \N__22405\,
            in3 => \N__24499\,
            lcout => \c0.n12_adj_2549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i70_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45385\,
            in1 => \N__20712\,
            in2 => \_gnd_net_\,
            in3 => \N__32909\,
            lcout => data_in_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1035_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21976\,
            in1 => \N__22511\,
            in2 => \N__20696\,
            in3 => \N__20669\,
            lcout => \c0.n9345\,
            ltout => \c0.n9345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_906_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28342\,
            in2 => \N__20642\,
            in3 => \N__24694\,
            lcout => \c0.n17532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25193\,
            in1 => \N__32983\,
            in2 => \N__20905\,
            in3 => \N__32064\,
            lcout => OPEN,
            ltout => \c0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i160_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23099\,
            in2 => \N__20639\,
            in3 => \N__21073\,
            lcout => \c0.data_out_frame2_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => \N__32828\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i167_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29506\,
            lcout => \c0.data_out_frame2_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => \N__32828\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_837_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29389\,
            lcout => \c0.n8995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i161_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20912\,
            in1 => \N__32214\,
            in2 => \N__20906\,
            in3 => \N__20891\,
            lcout => \c0.data_out_frame2_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => \N__32828\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_975_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24320\,
            in1 => \N__28693\,
            in2 => \_gnd_net_\,
            in3 => \N__29390\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i163_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23528\,
            in1 => \N__29279\,
            in2 => \N__20864\,
            in3 => \N__28850\,
            lcout => \c0.data_out_frame2_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => \N__32828\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i158_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__29391\,
            in2 => \N__36806\,
            in3 => \N__23126\,
            lcout => \c0.data_out_frame2_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50309\,
            ce => \N__32828\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i113_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35406\,
            in1 => \N__32751\,
            in2 => \_gnd_net_\,
            in3 => \N__20830\,
            lcout => data_out_frame2_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i147_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32747\,
            in1 => \N__34100\,
            in2 => \_gnd_net_\,
            in3 => \N__20812\,
            lcout => data_out_frame2_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i47_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36356\,
            in1 => \N__32752\,
            in2 => \_gnd_net_\,
            in3 => \N__20791\,
            lcout => data_out_frame2_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i52_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32748\,
            in1 => \N__35261\,
            in2 => \_gnd_net_\,
            in3 => \N__20773\,
            lcout => data_out_frame2_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i103_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35041\,
            in1 => \N__32750\,
            in2 => \_gnd_net_\,
            in3 => \N__20752\,
            lcout => data_out_frame2_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i93_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32749\,
            in1 => \N__35658\,
            in2 => \_gnd_net_\,
            in3 => \N__25670\,
            lcout => data_out_frame2_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i82_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35357\,
            in1 => \N__32753\,
            in2 => \_gnd_net_\,
            in3 => \N__23300\,
            lcout => data_out_frame2_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i111_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32746\,
            in1 => \N__36355\,
            in2 => \_gnd_net_\,
            in3 => \N__20959\,
            lcout => data_out_frame2_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i65_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__34212\,
            in2 => \_gnd_net_\,
            in3 => \N__20938\,
            lcout => data_out_frame2_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i148_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35209\,
            in1 => \N__26035\,
            in2 => \_gnd_net_\,
            in3 => \N__32638\,
            lcout => data_out_frame2_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i144_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32632\,
            in1 => \N__35459\,
            in2 => \_gnd_net_\,
            in3 => \N__21205\,
            lcout => data_out_frame2_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i124_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__23363\,
            in2 => \_gnd_net_\,
            in3 => \N__32636\,
            lcout => data_out_frame2_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i88_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32634\,
            in1 => \N__36005\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => data_out_frame2_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i72_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34963\,
            in1 => \N__23419\,
            in2 => \_gnd_net_\,
            in3 => \N__32639\,
            lcout => data_out_frame2_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i90_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__32635\,
            in1 => \N__34817\,
            in2 => \N__23315\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i140_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35717\,
            in1 => \N__25978\,
            in2 => \_gnd_net_\,
            in3 => \N__32637\,
            lcout => data_out_frame2_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i125_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35647\,
            in1 => \N__20995\,
            in2 => \_gnd_net_\,
            in3 => \N__32790\,
            lcout => data_out_frame2_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i39_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45292\,
            in1 => \N__28365\,
            in2 => \_gnd_net_\,
            in3 => \N__31270\,
            lcout => \c0.data_in_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i149_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35138\,
            in1 => \N__26260\,
            in2 => \_gnd_net_\,
            in3 => \N__32791\,
            lcout => data_out_frame2_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i85_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32788\,
            in1 => \N__36143\,
            in2 => \_gnd_net_\,
            in3 => \N__25687\,
            lcout => data_out_frame2_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i80_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__32787\,
            in1 => \N__36306\,
            in2 => \N__23435\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i101_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35137\,
            in1 => \N__20980\,
            in2 => \_gnd_net_\,
            in3 => \N__32789\,
            lcout => data_out_frame2_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1096_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29392\,
            in1 => \N__28645\,
            in2 => \_gnd_net_\,
            in3 => \N__24318\,
            lcout => \c0.n17504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_838_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28974\,
            in2 => \_gnd_net_\,
            in3 => \N__28937\,
            lcout => OPEN,
            ltout => \c0.n17535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i159_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29323\,
            in1 => \N__21086\,
            in2 => \N__21104\,
            in3 => \N__36743\,
            lcout => \c0.data_out_frame2_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50345\,
            ce => \N__32792\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_852_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28694\,
            in2 => \_gnd_net_\,
            in3 => \N__32066\,
            lcout => \c0.n9240\,
            ltout => \c0.n9240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1117_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21064\,
            in1 => \N__29393\,
            in2 => \N__21077\,
            in3 => \N__29479\,
            lcout => \c0.n10_adj_2470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1110_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__29257\,
            in2 => \N__31520\,
            in3 => \N__25637\,
            lcout => \c0.n9131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1121_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36742\,
            in2 => \_gnd_net_\,
            in3 => \N__36692\,
            lcout => OPEN,
            ltout => \c0.n17409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i162_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36632\,
            in1 => \N__32216\,
            in2 => \N__21053\,
            in3 => \N__21050\,
            lcout => \c0.data_out_frame2_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50345\,
            ce => \N__32792\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i154_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32215\,
            in1 => \N__36631\,
            in2 => \_gnd_net_\,
            in3 => \N__28880\,
            lcout => \c0.data_out_frame2_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50345\,
            ce => \N__32792\,
            sr => \_gnd_net_\
        );

    \c0.n18420_bdd_4_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__26673\,
            in1 => \N__21020\,
            in2 => \N__23450\,
            in3 => \N__21173\,
            lcout => OPEN,
            ltout => \c0.n18423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21188\,
            in1 => \N__26674\,
            in2 => \N__21008\,
            in3 => \N__26520\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50355\,
            ce => \N__26417\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16091_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21232\,
            in1 => \N__31094\,
            in2 => \N__21221\,
            in3 => \N__30791\,
            lcout => OPEN,
            ltout => \c0.n18576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18576_bdd_4_lut_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31095\,
            in1 => \N__22427\,
            in2 => \N__21209\,
            in3 => \N__21206\,
            lcout => OPEN,
            ltout => \c0.n18579_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26841\,
            in1 => \N__23171\,
            in2 => \N__21191\,
            in3 => \N__26941\,
            lcout => \c0.n22_adj_2520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15970_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23396\,
            in1 => \N__26672\,
            in2 => \N__21182\,
            in3 => \N__26840\,
            lcout => \c0.n18420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__33326\,
            in2 => \_gnd_net_\,
            in3 => \N__33265\,
            lcout => \c0.FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50366\,
            ce => 'H',
            sr => \N__21167\
        );

    \c0.rx.i1_2_lut_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39656\,
            in2 => \_gnd_net_\,
            in3 => \N__39565\,
            lcout => \c0.rx.n79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_adj_824_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21326\,
            in2 => \_gnd_net_\,
            in3 => \N__21501\,
            lcout => \c0.tx2.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__21288\,
            in1 => \N__21533\,
            in2 => \N__21434\,
            in3 => \N__21512\,
            lcout => OPEN,
            ltout => \c0.tx2.n9568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21292\,
            in2 => \N__21527\,
            in3 => \N__21524\,
            lcout => \c0.tx2.tx2_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_4_lut_adj_823_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__21323\,
            in1 => \N__21426\,
            in2 => \N__21295\,
            in3 => \N__21467\,
            lcout => n9652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21324\,
            lcout => \c0.tx2.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i29_4_lut_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__26131\,
            in1 => \N__21506\,
            in2 => \N__21296\,
            in3 => \N__21479\,
            lcout => OPEN,
            ltout => \c0.tx2.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__21469\,
            in1 => \N__21325\,
            in2 => \N__21437\,
            in3 => \N__21430\,
            lcout => \c0.tx2.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4452_2_lut_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26185\,
            lcout => OPEN,
            ltout => \c0.tx2.n6812_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7506_4_lut_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__21293\,
            in1 => \N__26130\,
            in2 => \N__21236\,
            in3 => \N__25926\,
            lcout => n9922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i44_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45496\,
            in1 => \N__23678\,
            in2 => \_gnd_net_\,
            in3 => \N__22297\,
            lcout => data_in_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i52_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45497\,
            in1 => \N__25727\,
            in2 => \_gnd_net_\,
            in3 => \N__22296\,
            lcout => data_in_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21646\,
            in1 => \N__45488\,
            in2 => \_gnd_net_\,
            in3 => \N__27037\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15249_2_lut_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21645\,
            in2 => \_gnd_net_\,
            in3 => \N__27629\,
            lcout => OPEN,
            ltout => \c0.n17697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15315_4_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24002\,
            in1 => \N__21624\,
            in2 => \N__21632\,
            in3 => \N__36242\,
            lcout => \c0.n17765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45487\,
            in1 => \N__37566\,
            in2 => \_gnd_net_\,
            in3 => \N__27630\,
            lcout => \c0.data_in_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21628\,
            in1 => \N__37660\,
            in2 => \_gnd_net_\,
            in3 => \N__45493\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36243\,
            in1 => \_gnd_net_\,
            in2 => \N__45505\,
            in3 => \N__26989\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24003\,
            in1 => \N__45489\,
            in2 => \_gnd_net_\,
            in3 => \N__27115\,
            lcout => \c0.data_in_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1057_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24970\,
            in1 => \N__21607\,
            in2 => \N__21554\,
            in3 => \N__22034\,
            lcout => n9054,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__24378\,
            in1 => \N__28142\,
            in2 => \N__45503\,
            in3 => \_gnd_net_\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28143\,
            in1 => \N__45474\,
            in2 => \_gnd_net_\,
            in3 => \N__23737\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i11_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__24125\,
            in1 => \N__28144\,
            in2 => \N__22042\,
            in3 => \N__31974\,
            lcout => \c0.data_in_frame_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_951_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22010\,
            in1 => \N__27509\,
            in2 => \_gnd_net_\,
            in3 => \N__28773\,
            lcout => \c0.n9208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1113_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24759\,
            in1 => \N__21977\,
            in2 => \N__21953\,
            in3 => \N__22544\,
            lcout => n9100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_969_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22451\,
            in1 => \N__21908\,
            in2 => \N__28979\,
            in3 => \N__21833\,
            lcout => n6_adj_2583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37518\,
            in1 => \N__24377\,
            in2 => \N__45504\,
            in3 => \_gnd_net_\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_861_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22155\,
            in1 => \N__21869\,
            in2 => \N__21838\,
            in3 => \N__21785\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_959_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21768\,
            in1 => \N__21727\,
            in2 => \N__21689\,
            in3 => \N__21686\,
            lcout => \c0.n8695\,
            ltout => \c0.n8695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_886_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22193\,
            in3 => \N__28335\,
            lcout => \c0.n8064\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1049_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000111100"
        )
    port map (
            in0 => \N__25112\,
            in1 => \N__23065\,
            in2 => \N__36961\,
            in3 => \N__24069\,
            lcout => \c0.n8867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i7_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24071\,
            in1 => \N__22161\,
            in2 => \N__31996\,
            in3 => \N__27749\,
            lcout => \c0.data_in_frame_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i29_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__27908\,
            in1 => \N__24072\,
            in2 => \N__22133\,
            in3 => \N__31988\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i3_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__24070\,
            in1 => \N__29001\,
            in2 => \N__31995\,
            in3 => \N__23741\,
            lcout => \c0.data_in_frame_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i41_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45460\,
            in1 => \N__22086\,
            in2 => \_gnd_net_\,
            in3 => \N__23830\,
            lcout => data_in_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3919_3_lut_4_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__22856\,
            in1 => \N__34553\,
            in2 => \N__22063\,
            in3 => \N__28008\,
            lcout => n2585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i63_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__38761\,
            in2 => \_gnd_net_\,
            in3 => \N__22059\,
            lcout => data_in_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i55_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__31287\,
            in1 => \N__45456\,
            in2 => \N__22064\,
            in3 => \_gnd_net_\,
            lcout => data_in_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i57_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45454\,
            in1 => \N__23905\,
            in2 => \_gnd_net_\,
            in3 => \N__24598\,
            lcout => data_in_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3935_3_lut_4_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__23043\,
            in1 => \N__34552\,
            in2 => \N__31291\,
            in3 => \N__28007\,
            lcout => n2593,
            ltout => \n2593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__28920\,
            in1 => \N__22261\,
            in2 => \N__22361\,
            in3 => \N__24901\,
            lcout => \c0.n22_adj_2461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3921_3_lut_4_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__28492\,
            in1 => \N__34554\,
            in2 => \N__36223\,
            in3 => \N__28009\,
            lcout => n2586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1103_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27516\,
            in1 => \N__22334\,
            in2 => \N__22705\,
            in3 => \N__24781\,
            lcout => \c0.n17412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3929_3_lut_4_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__37016\,
            in1 => \N__34569\,
            in2 => \N__22695\,
            in3 => \N__28004\,
            lcout => n2590,
            ltout => \n2590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_885_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22768\,
            in1 => \N__22496\,
            in2 => \N__22313\,
            in3 => \N__24758\,
            lcout => \c0.n10_adj_2450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3941_3_lut_4_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__22902\,
            in1 => \N__34570\,
            in2 => \N__22304\,
            in3 => \N__28005\,
            lcout => n2596,
            ltout => \n2596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_971_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111001111101"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__25346\,
            in2 => \N__22244\,
            in3 => \N__24476\,
            lcout => \c0.n10_adj_2498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3925_3_lut_4_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__22224\,
            in1 => \N__34571\,
            in2 => \N__25723\,
            in3 => \N__28006\,
            lcout => n2588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1053_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101001"
        )
    port map (
            in0 => \N__22769\,
            in1 => \N__22729\,
            in2 => \N__24698\,
            in3 => \N__24482\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i58_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22712\,
            in2 => \_gnd_net_\,
            in3 => \N__31906\,
            lcout => \c0.data_in_frame_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1106_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22653\,
            in1 => \N__22636\,
            in2 => \N__22590\,
            in3 => \N__22552\,
            lcout => \c0.n17403\,
            ltout => \c0.n17403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_985_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24438\,
            in1 => \N__22926\,
            in2 => \N__22499\,
            in3 => \N__22492\,
            lcout => n9283,
            ltout => \n9283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_3_lut_4_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25587\,
            in1 => \N__25064\,
            in2 => \N__22430\,
            in3 => \N__28094\,
            lcout => n16_adj_2656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i136_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34964\,
            in1 => \N__22420\,
            in2 => \_gnd_net_\,
            in3 => \N__32833\,
            lcout => data_out_frame2_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13614_3_lut_4_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__38801\,
            in1 => \N__34605\,
            in2 => \N__29245\,
            in3 => \N__34446\,
            lcout => \c0.n15927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_974_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22927\,
            in1 => \N__24439\,
            in2 => \_gnd_net_\,
            in3 => \N__28481\,
            lcout => \c0.n9219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_829_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28339\,
            in2 => \_gnd_net_\,
            in3 => \N__25331\,
            lcout => \c0.n17519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28254\,
            in1 => \N__28563\,
            in2 => \N__24614\,
            in3 => \N__23066\,
            lcout => OPEN,
            ltout => \c0.n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23051\,
            in1 => \N__23023\,
            in2 => \N__22991\,
            in3 => \N__22988\,
            lcout => OPEN,
            ltout => \c0.n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28397\,
            in1 => \N__22982\,
            in2 => \N__22976\,
            in3 => \N__22862\,
            lcout => \c0.n9355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i86_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32936\,
            in2 => \_gnd_net_\,
            in3 => \N__31973\,
            lcout => \c0.data_in_frame_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_adj_907_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__28341\,
            in2 => \N__24691\,
            in3 => \N__22871\,
            lcout => \c0.n11_adj_2453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22961\,
            in1 => \N__22903\,
            in2 => \_gnd_net_\,
            in3 => \N__22928\,
            lcout => \c0.n9144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22904\,
            in1 => \N__25525\,
            in2 => \_gnd_net_\,
            in3 => \N__22870\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_980_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22846\,
            in1 => \N__28491\,
            in2 => \N__22801\,
            in3 => \N__22784\,
            lcout => \c0.n17582\,
            ltout => \c0.n17582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i168_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23174\,
            in3 => \N__23098\,
            lcout => \c0.data_out_frame2_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50310\,
            ce => \N__32814\,
            sr => \_gnd_net_\
        );

    \c0.i3869_3_lut_4_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__34628\,
            in1 => \N__30473\,
            in2 => \N__36685\,
            in3 => \N__34445\,
            lcout => n2560,
            ltout => \n2560_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_860_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23144\,
            in1 => \N__23135\,
            in2 => \N__23129\,
            in3 => \N__23083\,
            lcout => OPEN,
            ltout => \c0.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_867_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111011"
        )
    port map (
            in0 => \N__23125\,
            in1 => \N__23108\,
            in2 => \N__23102\,
            in3 => \N__24470\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_928_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36872\,
            in1 => \N__32264\,
            in2 => \N__36625\,
            in3 => \N__36579\,
            lcout => \c0.n17418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3893_3_lut_4_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__34627\,
            in1 => \N__29681\,
            in2 => \N__36581\,
            in3 => \N__34444\,
            lcout => n2572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29700\,
            in1 => \N__29659\,
            in2 => \_gnd_net_\,
            in3 => \N__23072\,
            lcout => n18104,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => \c0.tx.n16357\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29712\,
            in1 => \N__29582\,
            in2 => \_gnd_net_\,
            in3 => \N__23069\,
            lcout => n18101,
            ltout => OPEN,
            carryin => \c0.tx.n16357\,
            carryout => \c0.tx.n16358\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29699\,
            in1 => \N__33794\,
            in2 => \_gnd_net_\,
            in3 => \N__23228\,
            lcout => n18102,
            ltout => OPEN,
            carryin => \c0.tx.n16358\,
            carryout => \c0.tx.n16359\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29713\,
            in1 => \N__29620\,
            in2 => \_gnd_net_\,
            in3 => \N__23225\,
            lcout => n18103,
            ltout => OPEN,
            carryin => \c0.tx.n16359\,
            carryout => \c0.tx.n16360\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29701\,
            in1 => \N__29602\,
            in2 => \_gnd_net_\,
            in3 => \N__23222\,
            lcout => n18097,
            ltout => OPEN,
            carryin => \c0.tx.n16360\,
            carryout => \c0.tx.n16361\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29714\,
            in1 => \N__29640\,
            in2 => \_gnd_net_\,
            in3 => \N__23219\,
            lcout => n18054,
            ltout => OPEN,
            carryin => \c0.tx.n16361\,
            carryout => \c0.tx.n16362\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__33832\,
            in1 => \N__37265\,
            in2 => \_gnd_net_\,
            in3 => \N__23216\,
            lcout => n18010,
            ltout => OPEN,
            carryin => \c0.tx.n16362\,
            carryout => \c0.tx.n16363\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__33831\,
            in1 => \N__37229\,
            in2 => \_gnd_net_\,
            in3 => \N__23213\,
            lcout => n17952,
            ltout => OPEN,
            carryin => \c0.tx.n16363\,
            carryout => \c0.tx.n16364\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__37325\,
            in1 => \N__33833\,
            in2 => \_gnd_net_\,
            in3 => \N__23210\,
            lcout => n17950,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i133_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32743\,
            in1 => \_gnd_net_\,
            in2 => \N__35149\,
            in3 => \N__26221\,
            lcout => data_out_frame2_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1081_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25636\,
            in1 => \N__28692\,
            in2 => \_gnd_net_\,
            in3 => \N__32045\,
            lcout => n9051,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_870_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__33272\,
            in1 => \N__25132\,
            in2 => \N__33367\,
            in3 => \N__23207\,
            lcout => \c0.n136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i79_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32744\,
            in1 => \N__36354\,
            in2 => \_gnd_net_\,
            in3 => \N__23377\,
            lcout => data_out_frame2_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i116_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35250\,
            in1 => \N__23350\,
            in2 => \_gnd_net_\,
            in3 => \N__32745\,
            lcout => data_out_frame2_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16041_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__30695\,
            in1 => \N__23362\,
            in2 => \N__23351\,
            in3 => \N__31052\,
            lcout => OPEN,
            ltout => \c0.n18516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18516_bdd_4_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31053\,
            in1 => \N__25777\,
            in2 => \N__23336\,
            in3 => \N__23333\,
            lcout => \c0.n17818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16011_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__23311\,
            in1 => \N__23299\,
            in2 => \N__31096\,
            in3 => \N__30694\,
            lcout => \c0.n18480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12304_4_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110010"
        )
    port map (
            in0 => \N__33514\,
            in1 => \N__23276\,
            in2 => \N__33148\,
            in3 => \N__23270\,
            lcout => \c0.n14631\,
            ltout => \c0.n14631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i5_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__33666\,
            in1 => \_gnd_net_\,
            in2 => \N__23252\,
            in3 => \N__26710\,
            lcout => \c0.data_out_frame2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i3_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__23242\,
            in1 => \N__33667\,
            in2 => \_gnd_net_\,
            in3 => \N__25789\,
            lcout => \c0.data_out_frame2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i45_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__36459\,
            in1 => \N__26863\,
            in2 => \N__32842\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i68_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32834\,
            in2 => \N__23492\,
            in3 => \N__35194\,
            lcout => data_out_frame2_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_843_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32987\,
            in2 => \_gnd_net_\,
            in3 => \N__36686\,
            lcout => \c0.n17482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18522_bdd_4_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__31075\,
            in1 => \N__23509\,
            in2 => \N__23491\,
            in3 => \N__23477\,
            lcout => \c0.n17815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15819_3_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__30722\,
            in1 => \N__23468\,
            in2 => \_gnd_net_\,
            in3 => \N__31074\,
            lcout => \c0.n18076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18588_bdd_4_lut_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__31073\,
            in1 => \N__23431\,
            in2 => \N__23420\,
            in3 => \N__23405\,
            lcout => \c0.n17785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i0_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34201\,
            in2 => \_gnd_net_\,
            in3 => \N__23387\,
            lcout => rand_data_0,
            ltout => OPEN,
            carryin => \bfn_5_29_0_\,
            carryout => n16319,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i1_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34139\,
            in2 => \_gnd_net_\,
            in3 => \N__23384\,
            lcout => rand_data_1,
            ltout => OPEN,
            carryin => n16319,
            carryout => n16320,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i2_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34078\,
            in2 => \_gnd_net_\,
            in3 => \N__23381\,
            lcout => rand_data_2,
            ltout => OPEN,
            carryin => n16320,
            carryout => n16321,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i3_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35190\,
            in2 => \_gnd_net_\,
            in3 => \N__23555\,
            lcout => rand_data_3,
            ltout => OPEN,
            carryin => n16321,
            carryout => n16322,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i4_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35133\,
            in2 => \_gnd_net_\,
            in3 => \N__23552\,
            lcout => rand_data_4,
            ltout => OPEN,
            carryin => n16322,
            carryout => n16323,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i5_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35071\,
            in2 => \_gnd_net_\,
            in3 => \N__23549\,
            lcout => rand_data_5,
            ltout => OPEN,
            carryin => n16323,
            carryout => n16324,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i6_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35013\,
            in2 => \_gnd_net_\,
            in3 => \N__23546\,
            lcout => rand_data_6,
            ltout => OPEN,
            carryin => n16324,
            carryout => n16325,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i7_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34938\,
            in2 => \_gnd_net_\,
            in3 => \N__23543\,
            lcout => rand_data_7,
            ltout => OPEN,
            carryin => n16325,
            carryout => n16326,
            clk => \N__50356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i8_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34856\,
            in2 => \_gnd_net_\,
            in3 => \N__23540\,
            lcout => rand_data_8,
            ltout => OPEN,
            carryin => \bfn_5_30_0_\,
            carryout => n16327,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i9_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34801\,
            in2 => \_gnd_net_\,
            in3 => \N__23537\,
            lcout => rand_data_9,
            ltout => OPEN,
            carryin => n16327,
            carryout => n16328,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i10_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34736\,
            in2 => \_gnd_net_\,
            in3 => \N__23534\,
            lcout => rand_data_10,
            ltout => OPEN,
            carryin => n16328,
            carryout => n16329,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i11_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35685\,
            in2 => \_gnd_net_\,
            in3 => \N__23531\,
            lcout => rand_data_11,
            ltout => OPEN,
            carryin => n16329,
            carryout => n16330,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i12_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35632\,
            in2 => \_gnd_net_\,
            in3 => \N__23585\,
            lcout => rand_data_12,
            ltout => OPEN,
            carryin => n16330,
            carryout => n16331,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i13_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35563\,
            in2 => \_gnd_net_\,
            in3 => \N__23582\,
            lcout => rand_data_13,
            ltout => OPEN,
            carryin => n16331,
            carryout => n16332,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i14_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35503\,
            in2 => \_gnd_net_\,
            in3 => \N__23579\,
            lcout => rand_data_14,
            ltout => OPEN,
            carryin => n16332,
            carryout => n16333,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i15_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35437\,
            in2 => \_gnd_net_\,
            in3 => \N__23576\,
            lcout => rand_data_15,
            ltout => OPEN,
            carryin => n16333,
            carryout => n16334,
            clk => \N__50367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i16_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35386\,
            in2 => \_gnd_net_\,
            in3 => \N__23573\,
            lcout => rand_data_16,
            ltout => OPEN,
            carryin => \bfn_5_31_0_\,
            carryout => n16335,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i17_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35335\,
            in2 => \_gnd_net_\,
            in3 => \N__23570\,
            lcout => rand_data_17,
            ltout => OPEN,
            carryin => n16335,
            carryout => n16336,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i18_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35283\,
            in2 => \_gnd_net_\,
            in3 => \N__23567\,
            lcout => rand_data_18,
            ltout => OPEN,
            carryin => n16336,
            carryout => n16337,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i19_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35239\,
            in2 => \_gnd_net_\,
            in3 => \N__23564\,
            lcout => rand_data_19,
            ltout => OPEN,
            carryin => n16337,
            carryout => n16338,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i20_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36131\,
            in2 => \_gnd_net_\,
            in3 => \N__23561\,
            lcout => rand_data_20,
            ltout => OPEN,
            carryin => n16338,
            carryout => n16339,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i21_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36076\,
            in2 => \_gnd_net_\,
            in3 => \N__23558\,
            lcout => rand_data_21,
            ltout => OPEN,
            carryin => n16339,
            carryout => n16340,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i22_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36027\,
            in2 => \_gnd_net_\,
            in3 => \N__23612\,
            lcout => rand_data_22,
            ltout => OPEN,
            carryin => n16340,
            carryout => n16341,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i23_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35978\,
            in2 => \_gnd_net_\,
            in3 => \N__23609\,
            lcout => rand_data_23,
            ltout => OPEN,
            carryin => n16341,
            carryout => n16342,
            clk => \N__50375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i24_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35920\,
            in2 => \_gnd_net_\,
            in3 => \N__23606\,
            lcout => rand_data_24,
            ltout => OPEN,
            carryin => \bfn_5_32_0_\,
            carryout => n16343,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i25_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35860\,
            in2 => \_gnd_net_\,
            in3 => \N__23603\,
            lcout => rand_data_25,
            ltout => OPEN,
            carryin => n16343,
            carryout => n16344,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i26_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35796\,
            in2 => \_gnd_net_\,
            in3 => \N__23600\,
            lcout => rand_data_26,
            ltout => OPEN,
            carryin => n16344,
            carryout => n16345,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i27_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35749\,
            in2 => \_gnd_net_\,
            in3 => \N__23597\,
            lcout => rand_data_27,
            ltout => OPEN,
            carryin => n16345,
            carryout => n16346,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i28_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36437\,
            in2 => \_gnd_net_\,
            in3 => \N__23594\,
            lcout => rand_data_28,
            ltout => OPEN,
            carryin => n16346,
            carryout => n16347,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i29_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36383\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => rand_data_29,
            ltout => OPEN,
            carryin => n16347,
            carryout => n16348,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i30_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36335\,
            in2 => \_gnd_net_\,
            in3 => \N__23588\,
            lcout => rand_data_30,
            ltout => OPEN,
            carryin => n16348,
            carryout => n16349,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2269__i31_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36287\,
            in2 => \_gnd_net_\,
            in3 => \N__23705\,
            lcout => rand_data_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45501\,
            in1 => \N__27275\,
            in2 => \_gnd_net_\,
            in3 => \N__23947\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i36_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45502\,
            in1 => \N__27564\,
            in2 => \_gnd_net_\,
            in3 => \N__23679\,
            lcout => data_in_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15296_4_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23945\,
            in1 => \N__27173\,
            in2 => \N__23977\,
            in3 => \N__27782\,
            lcout => \c0.n17745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27174\,
            in1 => \N__45418\,
            in2 => \_gnd_net_\,
            in3 => \N__27199\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15266_3_lut_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27271\,
            in1 => \N__26977\,
            in2 => \_gnd_net_\,
            in3 => \N__27062\,
            lcout => OPEN,
            ltout => \c0.n17715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_941_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__27103\,
            in2 => \N__23654\,
            in3 => \N__23924\,
            lcout => \c0.n8_adj_2474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16061_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__30770\,
            in1 => \N__25655\,
            in2 => \N__23651\,
            in3 => \N__31124\,
            lcout => \c0.n18540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27232\,
            in1 => \N__45419\,
            in2 => \_gnd_net_\,
            in3 => \N__23946\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23973\,
            in1 => \_gnd_net_\,
            in2 => \N__45484\,
            in3 => \N__24007\,
            lcout => \c0.data_in_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_940_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23969\,
            in2 => \_gnd_net_\,
            in3 => \N__23944\,
            lcout => \c0.n6_adj_2473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i53_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27454\,
            in1 => \_gnd_net_\,
            in2 => \N__45485\,
            in3 => \N__27426\,
            lcout => \c0.data_in_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i65_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29419\,
            in1 => \_gnd_net_\,
            in2 => \N__45486\,
            in3 => \N__23893\,
            lcout => data_in_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i2_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__33158\,
            in1 => \N__31171\,
            in2 => \N__33693\,
            in3 => \N__23882\,
            lcout => \c0.data_out_frame2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3947_3_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23831\,
            in1 => \N__23804\,
            in2 => \_gnd_net_\,
            in3 => \N__24118\,
            lcout => n2599,
            ltout => \n2599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_893_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001111011"
        )
    port map (
            in0 => \N__24560\,
            in1 => \N__28591\,
            in2 => \N__23756\,
            in3 => \N__27466\,
            lcout => \c0.n20_adj_2452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_934_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27315\,
            in1 => \N__27536\,
            in2 => \N__31410\,
            in3 => \N__27707\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_937_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27680\,
            in1 => \N__23736\,
            in2 => \N__23720\,
            in3 => \N__23717\,
            lcout => \c0.n8556\,
            ltout => \c0.n8556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_944_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24395\,
            in3 => \N__27740\,
            lcout => \c0.n6_adj_2478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27133\,
            in2 => \_gnd_net_\,
            in3 => \N__24343\,
            lcout => OPEN,
            ltout => \c0.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_947_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__28141\,
            in1 => \N__28183\,
            in2 => \N__24392\,
            in3 => \N__31378\,
            lcout => n63,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_946_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__27872\,
            in2 => \N__37553\,
            in3 => \N__24389\,
            lcout => \c0.n8460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_956_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24379\,
            in1 => \N__27280\,
            in2 => \N__28117\,
            in3 => \N__24344\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1010_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__27604\,
            in1 => \N__24332\,
            in2 => \N__24323\,
            in3 => \N__26951\,
            lcout => n63_adj_2642,
            ltout => \n63_adj_2642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10279_3_lut_4_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__34550\,
            in1 => \N__24317\,
            in2 => \N__24281\,
            in3 => \N__39845\,
            lcout => n2561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1009_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__34307\,
            in1 => \_gnd_net_\,
            in2 => \N__34408\,
            in3 => \N__34548\,
            lcout => n16468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1011_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34308\,
            in2 => \_gnd_net_\,
            in3 => \N__34367\,
            lcout => \c0.n4_adj_2512\,
            ltout => \c0.n4_adj_2512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10772_3_lut_4_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__24594\,
            in1 => \N__25472\,
            in2 => \N__24578\,
            in3 => \N__34549\,
            lcout => n2591,
            ltout => \n2591_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_902_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24555\,
            in1 => \N__24524\,
            in2 => \N__24506\,
            in3 => \N__24503\,
            lcout => \c0.n17533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3959_3_lut_4_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__24763\,
            in1 => \N__34551\,
            in2 => \N__33037\,
            in3 => \N__28035\,
            lcout => \c0.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3889_3_lut_4_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__34394\,
            in1 => \N__36597\,
            in2 => \N__34642\,
            in3 => \N__32908\,
            lcout => n2570,
            ltout => \n2570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i78_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24458\,
            in3 => \N__31907\,
            lcout => \c0.data_in_frame_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1013_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24455\,
            in1 => \N__27904\,
            in2 => \N__28118\,
            in3 => \N__27140\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1014_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__27741\,
            in1 => \N__27824\,
            in2 => \N__24446\,
            in3 => \N__37472\,
            lcout => \FRAME_MATCHER_next_state_31_N_2026_1\,
            ltout => \FRAME_MATCHER_next_state_31_N_2026_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3943_3_lut_4_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__24443\,
            in2 => \N__24419\,
            in3 => \N__28033\,
            lcout => n2597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3883_3_lut_4_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__29926\,
            in1 => \N__34594\,
            in2 => \N__25631\,
            in3 => \N__34393\,
            lcout => n2567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_898_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25389\,
            in1 => \N__24879\,
            in2 => \_gnd_net_\,
            in3 => \N__24994\,
            lcout => \c0.n17575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3961_3_lut_4_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__28043\,
            in1 => \N__24971\,
            in2 => \N__39892\,
            in3 => \N__34575\,
            lcout => \c0.n2606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3951_3_lut_4_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34574\,
            in1 => \N__28042\,
            in2 => \N__24692\,
            in3 => \N__31263\,
            lcout => OPEN,
            ltout => \c0.n2601_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_968_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24791\,
            in1 => \N__24935\,
            in2 => \N__24911\,
            in3 => \N__24900\,
            lcout => \c0.n11_adj_2494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1043_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25444\,
            in1 => \N__24883\,
            in2 => \N__25403\,
            in3 => \N__28196\,
            lcout => OPEN,
            ltout => \c0.n17428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_981_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__24848\,
            in1 => \N__24821\,
            in2 => \N__24815\,
            in3 => \N__24812\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1058_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__24753\,
            in2 => \_gnd_net_\,
            in3 => \N__24790\,
            lcout => \c0.n9103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_900_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24682\,
            lcout => \c0.n17430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3955_3_lut_4_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34576\,
            in1 => \N__28044\,
            in2 => \N__27403\,
            in3 => \N__25277\,
            lcout => \c0.n2603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3885_3_lut_4_lut_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__29828\,
            in1 => \N__34640\,
            in2 => \N__32263\,
            in3 => \N__34434\,
            lcout => n2568,
            ltout => \n2568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111001111101"
        )
    port map (
            in0 => \N__25208\,
            in1 => \N__25189\,
            in2 => \N__25178\,
            in3 => \N__31450\,
            lcout => OPEN,
            ltout => \c0.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_866_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__25174\,
            in1 => \N__27914\,
            in2 => \N__25145\,
            in3 => \N__32935\,
            lcout => OPEN,
            ltout => \c0.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28781\,
            in1 => \N__25142\,
            in2 => \N__25136\,
            in3 => \N__28499\,
            lcout => \c0.n5_adj_2438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3897_3_lut_4_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__27657\,
            in1 => \N__34641\,
            in2 => \N__36741\,
            in3 => \N__34433\,
            lcout => n2574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i74_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45344\,
            in1 => \N__29531\,
            in2 => \_gnd_net_\,
            in3 => \N__27658\,
            lcout => data_in_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50311\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1119_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28098\,
            in2 => \_gnd_net_\,
            in3 => \N__25108\,
            lcout => \c0.n4_adj_2548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_1131_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25063\,
            lcout => n19_adj_2651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i35_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45280\,
            in1 => \N__29844\,
            in2 => \_gnd_net_\,
            in3 => \N__33027\,
            lcout => data_in_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25588\,
            in2 => \_gnd_net_\,
            in3 => \N__28439\,
            lcout => OPEN,
            ltout => \n6_adj_2604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25529\,
            in1 => \N__25501\,
            in2 => \N__25475\,
            in3 => \N__25471\,
            lcout => n17547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1046_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25443\,
            in1 => \N__29762\,
            in2 => \N__25399\,
            in3 => \N__25361\,
            lcout => \c0.n8666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i114_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35356\,
            in1 => \N__25309\,
            in2 => \_gnd_net_\,
            in3 => \N__32815\,
            lcout => data_out_frame2_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40371\,
            in1 => \N__25295\,
            in2 => \_gnd_net_\,
            in3 => \N__29660\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27326\,
            in1 => \N__37648\,
            in2 => \_gnd_net_\,
            in3 => \N__45245\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40372\,
            in1 => \N__29603\,
            in2 => \_gnd_net_\,
            in3 => \N__25289\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29621\,
            in1 => \N__25283\,
            in2 => \_gnd_net_\,
            in3 => \N__40374\,
            lcout => \r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i60_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25710\,
            in1 => \N__29734\,
            in2 => \_gnd_net_\,
            in3 => \N__45246\,
            lcout => data_in_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40373\,
            in1 => \N__25694\,
            in2 => \_gnd_net_\,
            in3 => \N__29641\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25688\,
            in1 => \N__25669\,
            in2 => \_gnd_net_\,
            in3 => \N__30753\,
            lcout => \c0.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i123_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34049\,
            in1 => \_gnd_net_\,
            in2 => \N__45347\,
            in3 => \N__29881\,
            lcout => data_in_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i61_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30235\,
            in1 => \N__35662\,
            in2 => \_gnd_net_\,
            in3 => \N__32823\,
            lcout => data_out_frame2_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i80_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45238\,
            in1 => \N__29826\,
            in2 => \_gnd_net_\,
            in3 => \N__30472\,
            lcout => data_in_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i118_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36099\,
            in1 => \N__25651\,
            in2 => \_gnd_net_\,
            in3 => \N__32822\,
            lcout => data_out_frame2_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i165_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__38443\,
            in1 => \_gnd_net_\,
            in2 => \N__45348\,
            in3 => \N__29896\,
            lcout => data_in_20_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_953_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29258\,
            in2 => \_gnd_net_\,
            in3 => \N__25635\,
            lcout => \c0.n17559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11212_2_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39245\,
            in2 => \_gnd_net_\,
            in3 => \N__39307\,
            lcout => n13597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i107_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45226\,
            in1 => \N__34705\,
            in2 => \_gnd_net_\,
            in3 => \N__29870\,
            lcout => data_in_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i4_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__33645\,
            in1 => \N__25810\,
            in2 => \_gnd_net_\,
            in3 => \N__25790\,
            lcout => \c0.data_out_frame2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i100_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25778\,
            in1 => \N__35204\,
            in2 => \_gnd_net_\,
            in3 => \N__32832\,
            lcout => data_out_frame2_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i51_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33060\,
            in1 => \N__33763\,
            in2 => \_gnd_net_\,
            in3 => \N__45231\,
            lcout => data_in_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i155_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25766\,
            in1 => \_gnd_net_\,
            in2 => \N__45345\,
            in3 => \N__38464\,
            lcout => data_in_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i163_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30014\,
            in1 => \N__45227\,
            in2 => \_gnd_net_\,
            in3 => \N__25765\,
            lcout => data_in_20_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15930_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__26663\,
            in1 => \N__25757\,
            in2 => \N__25751\,
            in3 => \N__26846\,
            lcout => OPEN,
            ltout => \c0.n18372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18372_bdd_4_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__25796\,
            in1 => \N__25742\,
            in2 => \N__25730\,
            in3 => \N__26664\,
            lcout => OPEN,
            ltout => \c0.n18375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26665\,
            in1 => \N__25949\,
            in2 => \N__26054\,
            in3 => \N__26521\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50357\,
            ce => \N__26416\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16036_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__26039\,
            in1 => \N__31076\,
            in2 => \N__26021\,
            in3 => \N__30789\,
            lcout => OPEN,
            ltout => \c0.n18510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18510_bdd_4_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31077\,
            in1 => \N__26003\,
            in2 => \N__25985\,
            in3 => \N__25982\,
            lcout => OPEN,
            ltout => \c0.n18513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26845\,
            in1 => \N__25964\,
            in2 => \N__25952\,
            in3 => \N__26925\,
            lcout => \c0.n22_adj_2527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__25871\,
            in1 => \N__25943\,
            in2 => \N__26093\,
            in3 => \N__25910\,
            lcout => \r_Bit_Index_2_adj_2635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i153_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45232\,
            in1 => \N__37823\,
            in2 => \_gnd_net_\,
            in3 => \N__29938\,
            lcout => data_in_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26081\,
            in1 => \N__30375\,
            in2 => \N__29969\,
            in3 => \N__30316\,
            lcout => \r_Clock_Count_1_adj_2623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_955_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31516\,
            in1 => \N__32065\,
            in2 => \N__25847\,
            in3 => \N__28534\,
            lcout => n9135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15817_3_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__30790\,
            in1 => \N__25811\,
            in2 => \_gnd_net_\,
            in3 => \N__31123\,
            lcout => \c0.n18082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2450_2_lut_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26135\,
            lcout => n4980,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29988\,
            in2 => \_gnd_net_\,
            in3 => \N__26084\,
            lcout => n226,
            ltout => OPEN,
            carryin => \bfn_6_30_0_\,
            carryout => \c0.rx.n16365\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29965\,
            in3 => \N__26075\,
            lcout => n225,
            ltout => OPEN,
            carryin => \c0.rx.n16365\,
            carryout => \c0.rx.n16366\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30110\,
            in2 => \_gnd_net_\,
            in3 => \N__26072\,
            lcout => n224,
            ltout => OPEN,
            carryin => \c0.rx.n16366\,
            carryout => \c0.rx.n16367\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30070\,
            in2 => \_gnd_net_\,
            in3 => \N__26069\,
            lcout => n223,
            ltout => OPEN,
            carryin => \c0.rx.n16367\,
            carryout => \c0.rx.n16368\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30334\,
            in2 => \_gnd_net_\,
            in3 => \N__26066\,
            lcout => n222,
            ltout => OPEN,
            carryin => \c0.rx.n16368\,
            carryout => \c0.rx.n16369\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38101\,
            in2 => \_gnd_net_\,
            in3 => \N__26063\,
            lcout => n221,
            ltout => OPEN,
            carryin => \c0.rx.n16369\,
            carryout => \c0.rx.n16370\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__30119\,
            in1 => \N__37998\,
            in2 => \_gnd_net_\,
            in3 => \N__26060\,
            lcout => \c0.rx.n18001\,
            ltout => OPEN,
            carryin => \c0.rx.n16370\,
            carryout => \c0.rx.n16371\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__38055\,
            in1 => \N__30118\,
            in2 => \_gnd_net_\,
            in3 => \N__26057\,
            lcout => \c0.rx.n17999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__30108\,
            in1 => \N__26318\,
            in2 => \N__30317\,
            in3 => \N__30376\,
            lcout => \r_Clock_Count_2_adj_2622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26306\,
            in1 => \N__30373\,
            in2 => \N__29993\,
            in3 => \N__30310\,
            lcout => \r_Clock_Count_0_adj_2624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__30315\,
            in1 => \N__30377\,
            in2 => \N__38110\,
            in3 => \N__26300\,
            lcout => \r_Clock_Count_5_adj_2619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__26294\,
            in1 => \N__30374\,
            in2 => \N__30074\,
            in3 => \N__30314\,
            lcout => \r_Clock_Count_3_adj_2621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11152_2_lut_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30107\,
            in2 => \_gnd_net_\,
            in3 => \N__30068\,
            lcout => \c0.rx.n13537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30309\,
            in1 => \N__38056\,
            in2 => \_gnd_net_\,
            in3 => \N__26288\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18444_bdd_4_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__26273\,
            in2 => \N__31190\,
            in3 => \N__26842\,
            lcout => \c0.n18447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_16051_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__30795\,
            in1 => \N__26264\,
            in2 => \N__26243\,
            in3 => \N__31155\,
            lcout => OPEN,
            ltout => \c0.n18528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18528_bdd_4_lut_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31156\,
            in1 => \N__26225\,
            in2 => \N__26207\,
            in3 => \N__26204\,
            lcout => OPEN,
            ltout => \c0.n18531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__29294\,
            in1 => \N__26934\,
            in2 => \N__26870\,
            in3 => \N__26798\,
            lcout => \c0.n22_adj_2525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15709_2_lut_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26867\,
            in2 => \_gnd_net_\,
            in3 => \N__30796\,
            lcout => OPEN,
            ltout => \c0.n17955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_1__bdd_4_lut_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__30200\,
            in1 => \N__31157\,
            in2 => \N__26849\,
            in3 => \N__26799\,
            lcout => OPEN,
            ltout => \c0.n18456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18456_bdd_4_lut_4_lut_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100100"
        )
    port map (
            in0 => \N__26800\,
            in1 => \N__26714\,
            in2 => \N__26696\,
            in3 => \N__30797\,
            lcout => OPEN,
            ltout => \c0.n18459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11600217_i1_3_lut_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26693\,
            in2 => \N__26687\,
            in3 => \N__26666\,
            lcout => OPEN,
            ltout => \c0.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_6_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__26684\,
            in1 => \N__26678\,
            in2 => \N__26528\,
            in3 => \N__26525\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50391\,
            ce => \N__26404\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27364\,
            in1 => \_gnd_net_\,
            in2 => \N__45483\,
            in3 => \N__27895\,
            lcout => \c0.data_in_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27073\,
            in1 => \N__31377\,
            in2 => \_gnd_net_\,
            in3 => \N__45416\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45410\,
            in1 => \N__27175\,
            in2 => \_gnd_net_\,
            in3 => \N__26985\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27111\,
            in1 => \N__27835\,
            in2 => \_gnd_net_\,
            in3 => \N__45415\,
            lcout => \c0.data_in_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45409\,
            in1 => \N__27032\,
            in2 => \_gnd_net_\,
            in3 => \N__27276\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i40_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36916\,
            in1 => \N__27231\,
            in2 => \_gnd_net_\,
            in3 => \N__45417\,
            lcout => data_in_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i38_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__45411\,
            in2 => \_gnd_net_\,
            in3 => \N__27198\,
            lcout => data_in_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i46_2_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27596\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => OPEN,
            ltout => \c0.n28_adj_2475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_943_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27789\,
            in1 => \N__27172\,
            in2 => \N__27149\,
            in3 => \N__27146\,
            lcout => \c0.n8559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_957_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27104\,
            in1 => \N__27063\,
            in2 => \N__27033\,
            in3 => \N__26978\,
            lcout => \c0.n17_adj_2486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37552\,
            in1 => \N__45430\,
            in2 => \_gnd_net_\,
            in3 => \N__27538\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i82_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45429\,
            in1 => \N__31316\,
            in2 => \_gnd_net_\,
            in3 => \N__29523\,
            lcout => data_in_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__45432\,
            in2 => \_gnd_net_\,
            in3 => \N__27644\,
            lcout => \c0.data_in_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27571\,
            in1 => \N__45431\,
            in2 => \_gnd_net_\,
            in3 => \N__27537\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3923_3_lut_4_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__27517\,
            in1 => \N__34643\,
            in2 => \N__27455\,
            in3 => \N__28034\,
            lcout => n2587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i61_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45329\,
            in1 => \N__38377\,
            in2 => \_gnd_net_\,
            in3 => \N__27453\,
            lcout => \c0.data_in_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i45_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27427\,
            in1 => \N__45295\,
            in2 => \_gnd_net_\,
            in3 => \N__27390\,
            lcout => data_in_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i37_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27389\,
            in1 => \N__45330\,
            in2 => \_gnd_net_\,
            in3 => \N__27357\,
            lcout => \c0.data_in_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40375\,
            in1 => \N__27341\,
            in2 => \_gnd_net_\,
            in3 => \N__37199\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45294\,
            in1 => \N__27897\,
            in2 => \_gnd_net_\,
            in3 => \N__27314\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15294_4_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27896\,
            in1 => \N__27823\,
            in2 => \N__37612\,
            in3 => \N__37508\,
            lcout => \c0.n17743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27831\,
            in1 => \N__27866\,
            in2 => \_gnd_net_\,
            in3 => \N__45452\,
            lcout => \c0.data_in_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27796\,
            in1 => \_gnd_net_\,
            in2 => \N__45494\,
            in3 => \N__27742\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27714\,
            in1 => \N__28182\,
            in2 => \_gnd_net_\,
            in3 => \N__45451\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13622_3_lut_4_lut_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__38348\,
            in1 => \N__34606\,
            in2 => \N__31505\,
            in3 => \N__34426\,
            lcout => n2571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i73_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29927\,
            in1 => \N__29412\,
            in2 => \_gnd_net_\,
            in3 => \N__45453\,
            lcout => data_in_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45445\,
            in1 => \N__38506\,
            in2 => \_gnd_net_\,
            in3 => \N__27681\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27682\,
            in1 => \N__45447\,
            in2 => \_gnd_net_\,
            in3 => \N__31409\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i66_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45446\,
            in1 => \N__37032\,
            in2 => \_gnd_net_\,
            in3 => \N__27662\,
            lcout => data_in_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_828_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28493\,
            in2 => \_gnd_net_\,
            in3 => \N__28434\,
            lcout => \c0.n17473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45346\,
            in2 => \N__28385\,
            in3 => \N__28181\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3949_3_lut_4_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__28343\,
            in1 => \N__34572\,
            in2 => \N__36912\,
            in3 => \N__28023\,
            lcout => OPEN,
            ltout => \c0.n2600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_966_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28274\,
            in1 => \N__28262\,
            in2 => \N__28220\,
            in3 => \N__28216\,
            lcout => \c0.n10_adj_2493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_932_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__28174\,
            in1 => \N__31376\,
            in2 => \_gnd_net_\,
            in3 => \N__28148\,
            lcout => \c0.n8572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3937_3_lut_4_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__28100\,
            in1 => \N__34573\,
            in2 => \N__36190\,
            in3 => \N__28024\,
            lcout => n2594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i84_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31451\,
            in2 => \_gnd_net_\,
            in3 => \N__31972\,
            lcout => \c0.data_in_frame_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10244_3_lut_4_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__34436\,
            in1 => \N__36493\,
            in2 => \N__34644\,
            in3 => \N__32106\,
            lcout => n2573,
            ltout => \n2573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_1156_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29173\,
            in1 => \N__28774\,
            in2 => \N__27917\,
            in3 => \N__28732\,
            lcout => n17481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1122_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28978\,
            in1 => \N__28933\,
            in2 => \N__28646\,
            in3 => \N__28895\,
            lcout => \c0.n17536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3879_3_lut_4_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__36524\,
            in1 => \N__34601\,
            in2 => \N__32057\,
            in3 => \N__34435\,
            lcout => n2565,
            ltout => \n2565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__28873\,
            in1 => \N__28849\,
            in2 => \N__28829\,
            in3 => \N__28819\,
            lcout => OPEN,
            ltout => \c0.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_862_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111111111"
        )
    port map (
            in0 => \N__28807\,
            in1 => \N__31537\,
            in2 => \N__28790\,
            in3 => \N__28787\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_1130_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28775\,
            in2 => \_gnd_net_\,
            in3 => \N__28733\,
            lcout => n17479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3875_3_lut_4_lut_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__28679\,
            in2 => \N__34661\,
            in3 => \N__38330\,
            lcout => n2563,
            ltout => \n2563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1118_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28641\,
            in1 => \N__28595\,
            in2 => \N__28568\,
            in3 => \N__28564\,
            lcout => OPEN,
            ltout => \c0.n17592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__28535\,
            in1 => \N__29344\,
            in2 => \N__28502\,
            in3 => \N__29429\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3881_3_lut_4_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__29530\,
            in1 => \N__34622\,
            in2 => \N__36871\,
            in3 => \N__34454\,
            lcout => n2566,
            ltout => \n2566_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_841_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__29507\,
            in1 => \N__29480\,
            in2 => \N__29453\,
            in3 => \N__29446\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3899_3_lut_4_lut_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__29423\,
            in1 => \N__34626\,
            in2 => \N__29388\,
            in3 => \N__34456\,
            lcout => n2575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1091_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29246\,
            in2 => \_gnd_net_\,
            in3 => \N__36691\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i165_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29333\,
            in1 => \N__29269\,
            in2 => \N__29312\,
            in3 => \N__29309\,
            lcout => \c0.data_out_frame2_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50329\,
            ce => \N__32841\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31512\,
            lcout => \c0.n17488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i155_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29247\,
            in1 => \N__29210\,
            in2 => \N__29201\,
            in3 => \N__29177\,
            lcout => \c0.data_out_frame2_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50329\,
            ce => \N__32841\,
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1059_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29138\,
            in1 => \N__29093\,
            in2 => \N__29060\,
            in3 => \N__29012\,
            lcout => \c0.n10_adj_2536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29578\,
            in1 => \_gnd_net_\,
            in2 => \N__40370\,
            in3 => \N__29756\,
            lcout => \r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i68_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45250\,
            in1 => \N__29733\,
            in2 => \_gnd_net_\,
            in3 => \N__29677\,
            lcout => data_in_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40155\,
            in2 => \_gnd_net_\,
            in3 => \N__40350\,
            lcout => OPEN,
            ltout => \n8517_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1138_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__33086\,
            in1 => \N__37346\,
            in2 => \N__29717\,
            in3 => \N__33852\,
            lcout => n17366,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i76_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45251\,
            in1 => \_gnd_net_\,
            in2 => \N__36989\,
            in3 => \N__29676\,
            lcout => data_in_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33789\,
            in1 => \N__29658\,
            in2 => \N__29642\,
            in3 => \N__29619\,
            lcout => OPEN,
            ltout => \c0.tx.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5_3_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29601\,
            in2 => \N__29585\,
            in3 => \N__29577\,
            lcout => n16466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i46_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29553\,
            in1 => \N__36191\,
            in2 => \_gnd_net_\,
            in3 => \N__45248\,
            lcout => data_in_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i69_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35153\,
            in1 => \N__31204\,
            in2 => \_gnd_net_\,
            in3 => \N__32652\,
            lcout => data_out_frame2_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__33724\,
            in1 => \N__37909\,
            in2 => \N__37946\,
            in3 => \N__33709\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i145_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45247\,
            in1 => \N__37453\,
            in2 => \_gnd_net_\,
            in3 => \N__29942\,
            lcout => data_in_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i81_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29919\,
            in1 => \N__36785\,
            in2 => \_gnd_net_\,
            in3 => \N__45249\,
            lcout => data_in_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__33976\,
            in1 => \N__37941\,
            in2 => \N__29897\,
            in3 => \N__37910\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i115_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45066\,
            in1 => \N__29869\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => data_in_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i136_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__30406\,
            in2 => \_gnd_net_\,
            in3 => \N__31472\,
            lcout => data_in_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45067\,
            in1 => \N__29851\,
            in2 => \_gnd_net_\,
            in3 => \N__37507\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i72_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29827\,
            in1 => \N__29784\,
            in2 => \_gnd_net_\,
            in3 => \N__45068\,
            lcout => data_in_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__30139\,
            in1 => \N__39654\,
            in2 => \N__40459\,
            in3 => \N__39584\,
            lcout => n8567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i105_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35949\,
            in1 => \N__30040\,
            in2 => \_gnd_net_\,
            in3 => \N__32843\,
            lcout => data_out_frame2_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i150_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45233\,
            in1 => \N__30025\,
            in2 => \_gnd_net_\,
            in3 => \N__37721\,
            lcout => data_in_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i142_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30026\,
            in1 => \N__45234\,
            in2 => \_gnd_net_\,
            in3 => \N__34264\,
            lcout => data_in_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_4_lut_adj_820_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30140\,
            in1 => \N__39655\,
            in2 => \N__40460\,
            in3 => \N__39585\,
            lcout => n8562,
            ltout => \n8562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__34033\,
            in1 => \N__30013\,
            in2 => \N__30017\,
            in3 => \N__37894\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__39687\,
            in1 => \N__39556\,
            in2 => \N__37895\,
            in3 => \N__34245\,
            lcout => \c0.rx.n2\,
            ltout => \c0.rx.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_818_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__39521\,
            in1 => \N__39752\,
            in2 => \N__30002\,
            in3 => \N__30383\,
            lcout => \c0.rx.n4_adj_2424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_819_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__39754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29999\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30333\,
            in1 => \N__29992\,
            in2 => \_gnd_net_\,
            in3 => \N__29958\,
            lcout => \c0.rx.n124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__39690\,
            in1 => \N__34232\,
            in2 => \N__39771\,
            in3 => \N__30194\,
            lcout => \c0.rx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.n18594_bdd_4_lut_4_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100011"
        )
    port map (
            in0 => \N__34246\,
            in1 => \N__37876\,
            in2 => \N__38297\,
            in3 => \N__39689\,
            lcout => \c0.rx.n18597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30173\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_816_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39753\,
            in2 => \_gnd_net_\,
            in3 => \N__39688\,
            lcout => \c0.rx.n17381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__30085\,
            in2 => \N__38106\,
            in3 => \N__30157\,
            lcout => \c0.rx.r_SM_Main_2_N_2386_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15740_4_lut_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30158\,
            in1 => \N__38096\,
            in2 => \N__30089\,
            in3 => \N__30148\,
            lcout => OPEN,
            ltout => \c0.rx.n18003_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i57_4_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__30149\,
            in1 => \N__30138\,
            in2 => \N__30125\,
            in3 => \N__30251\,
            lcout => n13880,
            ltout => \n13880_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i7678_1_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30122\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.n10193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_813_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30109\,
            in1 => \N__30084\,
            in2 => \_gnd_net_\,
            in3 => \N__30069\,
            lcout => \c0.rx.n97\,
            ltout => \c0.rx.n97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_817_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38100\,
            in1 => \N__38054\,
            in2 => \N__30386\,
            in3 => \N__37997\,
            lcout => \c0.rx.n17345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__30294\,
            in1 => \N__30372\,
            in2 => \N__30341\,
            in3 => \N__30347\,
            lcout => \r_Clock_Count_4_adj_2620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37999\,
            in1 => \N__30293\,
            in2 => \_gnd_net_\,
            in3 => \N__30278\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15405_4_lut_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000110000"
        )
    port map (
            in0 => \N__49063\,
            in1 => \N__49039\,
            in2 => \N__49112\,
            in3 => \N__49087\,
            lcout => n17855,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15406_4_lut_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111001000"
        )
    port map (
            in0 => \N__49088\,
            in1 => \N__49111\,
            in2 => \N__49043\,
            in3 => \N__49064\,
            lcout => OPEN,
            ltout => \n17856_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15407_3_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__50459\,
            in1 => \_gnd_net_\,
            in2 => \N__30272\,
            in3 => \N__30269\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__38102\,
            in1 => \N__38050\,
            in2 => \N__38020\,
            in3 => \N__37993\,
            lcout => \c0.rx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50392\,
            ce => 'H',
            sr => \N__39608\
        );

    \c0.rx.i1_2_lut_adj_814_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38049\,
            in2 => \_gnd_net_\,
            in3 => \N__37992\,
            lcout => \c0.rx.n112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30239\,
            in1 => \N__30221\,
            in2 => \_gnd_net_\,
            in3 => \N__30794\,
            lcout => \c0.n5_adj_2425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30793\,
            in1 => \N__31226\,
            in2 => \_gnd_net_\,
            in3 => \N__31205\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15708_3_lut_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__31181\,
            in1 => \N__31154\,
            in2 => \_gnd_net_\,
            in3 => \N__30792\,
            lcout => \c0.n18086\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i88_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30446\,
            in1 => \N__44937\,
            in2 => \_gnd_net_\,
            in3 => \N__30462\,
            lcout => data_in_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i96_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30437\,
            in1 => \_gnd_net_\,
            in2 => \N__45153\,
            in3 => \N__30445\,
            lcout => data_in_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i104_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30428\,
            in1 => \N__44935\,
            in2 => \_gnd_net_\,
            in3 => \N__30436\,
            lcout => data_in_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i112_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30419\,
            in1 => \_gnd_net_\,
            in2 => \N__45152\,
            in3 => \N__30427\,
            lcout => data_in_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i120_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30395\,
            in1 => \N__44936\,
            in2 => \_gnd_net_\,
            in3 => \N__30418\,
            lcout => data_in_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i128_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44934\,
            in1 => \N__30394\,
            in2 => \_gnd_net_\,
            in3 => \N__30410\,
            lcout => data_in_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i114_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45433\,
            in1 => \N__31429\,
            in2 => \_gnd_net_\,
            in3 => \N__36761\,
            lcout => data_in_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_next_state_i1_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__34683\,
            in1 => \N__34453\,
            in2 => \N__33548\,
            in3 => \N__34318\,
            lcout => \FRAME_MATCHER_next_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3877_3_lut_4_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__36978\,
            in1 => \N__34662\,
            in2 => \N__36836\,
            in3 => \N__34447\,
            lcout => n2564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i106_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31333\,
            in1 => \N__31433\,
            in2 => \_gnd_net_\,
            in3 => \N__45350\,
            lcout => data_in_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31414\,
            in1 => \N__31363\,
            in2 => \_gnd_net_\,
            in3 => \N__45351\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i102_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45349\,
            in1 => \N__38615\,
            in2 => \_gnd_net_\,
            in3 => \N__32869\,
            lcout => data_in_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i98_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31334\,
            in1 => \N__31324\,
            in2 => \_gnd_net_\,
            in3 => \N__45352\,
            lcout => data_in_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i90_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31325\,
            in1 => \N__45353\,
            in2 => \_gnd_net_\,
            in3 => \N__31309\,
            lcout => data_in_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i47_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45253\,
            in1 => \N__31247\,
            in2 => \_gnd_net_\,
            in3 => \N__31298\,
            lcout => data_in_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i64_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35474\,
            in1 => \N__32278\,
            in2 => \_gnd_net_\,
            in3 => \N__32827\,
            lcout => data_out_frame2_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_935_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36857\,
            in1 => \N__32246\,
            in2 => \_gnd_net_\,
            in3 => \N__36831\,
            lcout => \c0.n17433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i56_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36948\,
            in1 => \N__32165\,
            in2 => \_gnd_net_\,
            in3 => \N__45254\,
            lcout => data_in_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i75_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31969\,
            in2 => \_gnd_net_\,
            in3 => \N__32126\,
            lcout => \c0.data_in_frame_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i83_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__31971\,
            in1 => \N__32078\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i82_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31968\,
            in2 => \_gnd_net_\,
            in3 => \N__32009\,
            lcout => \c0.data_in_frame_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i77_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__31970\,
            in1 => \N__31541\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i164_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45155\,
            in1 => \N__33998\,
            in2 => \_gnd_net_\,
            in3 => \N__38626\,
            lcout => data_in_20_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i144_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45154\,
            in1 => \N__31462\,
            in2 => \_gnd_net_\,
            in3 => \N__37133\,
            lcout => data_in_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Done_44_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110111000"
        )
    port map (
            in0 => \N__33077\,
            in1 => \N__36767\,
            in2 => \N__40369\,
            in3 => \N__32849\,
            lcout => n7364,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i43_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45156\,
            in1 => \_gnd_net_\,
            in2 => \N__33071\,
            in3 => \N__33014\,
            lcout => data_in_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3873_3_lut_4_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__34679\,
            in1 => \N__32919\,
            in2 => \N__32986\,
            in3 => \N__34448\,
            lcout => n2562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i79_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39844\,
            in1 => \N__38790\,
            in2 => \_gnd_net_\,
            in3 => \N__45163\,
            lcout => data_in_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i86_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45160\,
            in1 => \N__32858\,
            in2 => \_gnd_net_\,
            in3 => \N__32920\,
            lcout => data_in_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i78_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32921\,
            in1 => \N__45162\,
            in2 => \_gnd_net_\,
            in3 => \N__32892\,
            lcout => data_in_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i94_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45161\,
            in1 => \N__32857\,
            in2 => \_gnd_net_\,
            in3 => \N__32873\,
            lcout => data_in_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15809_2_lut_3_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40159\,
            in1 => \N__40403\,
            in2 => \_gnd_net_\,
            in3 => \N__40215\,
            lcout => n18098,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4717_4_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__42979\,
            in1 => \N__37280\,
            in2 => \N__40163\,
            in3 => \N__40402\,
            lcout => n7080,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_220_Select_0_i1_2_lut_4_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__34289\,
            in2 => \N__33388\,
            in3 => \N__33460\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => \c0.FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50349\,
            ce => 'H',
            sr => \N__33560\
        );

    \c0.select_220_Select_1_i1_2_lut_4_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33268\,
            in1 => \N__33547\,
            in2 => \N__33389\,
            in3 => \N__33459\,
            lcout => \c0.n1_adj_2437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_4_lut_adj_826_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37321\,
            in1 => \N__37215\,
            in2 => \N__37261\,
            in3 => \N__33860\,
            lcout => \r_SM_Main_2_N_2323_1\,
            ltout => \r_SM_Main_2_N_2323_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15308_4_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__40145\,
            in1 => \N__40339\,
            in2 => \N__33395\,
            in3 => \N__40213\,
            lcout => n17757,
            ltout => \n17757_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9716_4_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000001000"
        )
    port map (
            in0 => \N__39126\,
            in1 => \N__37442\,
            in2 => \N__33392\,
            in3 => \N__37395\,
            lcout => n12123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1048_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33380\,
            in2 => \_gnd_net_\,
            in3 => \N__33266\,
            lcout => \c0.n157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40325\,
            in1 => \N__33098\,
            in2 => \_gnd_net_\,
            in3 => \N__37254\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_4_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37253\,
            in1 => \N__37315\,
            in2 => \N__40237\,
            in3 => \N__37222\,
            lcout => n9390,
            ltout => \n9390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15234_3_lut_4_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111011"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__40102\,
            in2 => \N__33866\,
            in3 => \N__37362\,
            lcout => OPEN,
            ltout => \n17681_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15277_4_lut_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101111"
        )
    port map (
            in0 => \N__37363\,
            in1 => \N__33770\,
            in2 => \N__33863\,
            in3 => \N__33859\,
            lcout => n17356,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33803\,
            in1 => \N__40289\,
            in2 => \_gnd_net_\,
            in3 => \N__33793\,
            lcout => \r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i83_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45117\,
            in1 => \N__33881\,
            in2 => \_gnd_net_\,
            in3 => \N__36516\,
            lcout => data_in_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i11216_2_lut_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40101\,
            in2 => \_gnd_net_\,
            in3 => \N__40288\,
            lcout => n13601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i59_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45116\,
            in1 => \N__33931\,
            in2 => \_gnd_net_\,
            in3 => \N__33750\,
            lcout => data_in_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__37917\,
            in1 => \N__37117\,
            in2 => \N__33911\,
            in3 => \N__33731\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i167_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33953\,
            in1 => \N__33713\,
            in2 => \_gnd_net_\,
            in3 => \N__45141\,
            lcout => data_in_20_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000101000"
        )
    port map (
            in0 => \N__37440\,
            in1 => \N__39122\,
            in2 => \N__38925\,
            in3 => \N__38950\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i131_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38405\,
            in1 => \N__34045\,
            in2 => \_gnd_net_\,
            in3 => \N__45140\,
            lcout => data_in_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__34034\,
            in1 => \N__33903\,
            in2 => \N__33997\,
            in3 => \N__37918\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__37916\,
            in1 => \N__37702\,
            in2 => \N__33910\,
            in3 => \N__33980\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__7__3526_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46049\,
            in1 => \N__34907\,
            in2 => \_gnd_net_\,
            in3 => \N__45899\,
            lcout => data_out_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i159_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33952\,
            in1 => \N__45105\,
            in2 => \_gnd_net_\,
            in3 => \N__37774\,
            lcout => data_in_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__6__3527_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46048\,
            in1 => \N__34982\,
            in2 => \_gnd_net_\,
            in3 => \N__46134\,
            lcout => data_out_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i67_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36497\,
            in1 => \N__33924\,
            in2 => \_gnd_net_\,
            in3 => \N__45110\,
            lcout => data_in_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37952\,
            in1 => \N__33902\,
            in2 => \N__37754\,
            in3 => \N__37919\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i91_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34694\,
            in1 => \_gnd_net_\,
            in2 => \N__45252\,
            in3 => \N__33877\,
            lcout => data_in_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i99_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34709\,
            in1 => \N__45106\,
            in2 => \_gnd_net_\,
            in3 => \N__34693\,
            lcout => data_in_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15728_2_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43650\,
            in2 => \_gnd_net_\,
            in3 => \N__48420\,
            lcout => \c0.n17911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_next_state_i0_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101110111"
        )
    port map (
            in0 => \N__34685\,
            in1 => \N__34457\,
            in2 => \N__34288\,
            in3 => \N__34325\,
            lcout => \FRAME_MATCHER_next_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41476\,
            in1 => \N__41825\,
            in2 => \_gnd_net_\,
            in3 => \N__48421\,
            lcout => \c0.n5_adj_2488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i134_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45142\,
            in1 => \N__38725\,
            in2 => \_gnd_net_\,
            in3 => \N__34268\,
            lcout => data_in_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15793_2_lut_3_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__37914\,
            in1 => \N__39571\,
            in2 => \_gnd_net_\,
            in3 => \N__34253\,
            lcout => \c0.rx.n18066\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i0_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34211\,
            in2 => \N__39436\,
            in3 => \_gnd_net_\,
            lcout => rand_setpoint_0,
            ltout => OPEN,
            carryin => \bfn_9_29_0_\,
            carryout => n16412,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i1_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34148\,
            in2 => \N__39160\,
            in3 => \N__34115\,
            lcout => rand_setpoint_1,
            ltout => OPEN,
            carryin => n16412,
            carryout => n16413,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i2_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34088\,
            in2 => \N__37738\,
            in3 => \N__34052\,
            lcout => rand_setpoint_2,
            ltout => OPEN,
            carryin => n16413,
            carryout => n16414,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i3_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35205\,
            in2 => \N__43351\,
            in3 => \N__35156\,
            lcout => rand_setpoint_3,
            ltout => OPEN,
            carryin => n16414,
            carryout => n16415,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i4_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35139\,
            in2 => \N__38216\,
            in3 => \N__35102\,
            lcout => rand_setpoint_4,
            ltout => OPEN,
            carryin => n16415,
            carryout => n16416,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i5_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35087\,
            in2 => \N__39412\,
            in3 => \N__35045\,
            lcout => rand_setpoint_5,
            ltout => OPEN,
            carryin => n16416,
            carryout => n16417,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i6_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34978\,
            in2 => \N__35039\,
            in3 => \N__34967\,
            lcout => rand_setpoint_6,
            ltout => OPEN,
            carryin => n16417,
            carryout => n16418,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i7_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34951\,
            in2 => \N__34906\,
            in3 => \N__34889\,
            lcout => rand_setpoint_7,
            ltout => OPEN,
            carryin => n16418,
            carryout => n16419,
            clk => \N__50393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i8_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34867\,
            in2 => \N__41500\,
            in3 => \N__34832\,
            lcout => rand_setpoint_8,
            ltout => OPEN,
            carryin => \bfn_9_30_0_\,
            carryout => n16420,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i9_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34813\,
            in2 => \N__44209\,
            in3 => \N__34772\,
            lcout => rand_setpoint_9,
            ltout => OPEN,
            carryin => n16420,
            carryout => n16421,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i10_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34745\,
            in2 => \N__38126\,
            in3 => \N__34712\,
            lcout => rand_setpoint_10,
            ltout => OPEN,
            carryin => n16421,
            carryout => n16422,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i11_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35689\,
            in2 => \N__38192\,
            in3 => \N__35666\,
            lcout => rand_setpoint_11,
            ltout => OPEN,
            carryin => n16422,
            carryout => n16423,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i12_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35657\,
            in2 => \N__41716\,
            in3 => \N__35606\,
            lcout => rand_setpoint_12,
            ltout => OPEN,
            carryin => n16423,
            carryout => n16424,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i13_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35585\,
            in2 => \N__41410\,
            in3 => \N__35537\,
            lcout => rand_setpoint_13,
            ltout => OPEN,
            carryin => n16424,
            carryout => n16425,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i14_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40561\,
            in2 => \N__35522\,
            in3 => \N__35477\,
            lcout => rand_setpoint_14,
            ltout => OPEN,
            carryin => n16425,
            carryout => n16426,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i15_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35458\,
            in2 => \N__40588\,
            in3 => \N__35411\,
            lcout => rand_setpoint_15,
            ltout => OPEN,
            carryin => n16426,
            carryout => n16427,
            clk => \N__50398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i16_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35396\,
            in2 => \N__41845\,
            in3 => \N__35360\,
            lcout => rand_setpoint_16,
            ltout => OPEN,
            carryin => \bfn_9_31_0_\,
            carryout => n16428,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i17_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35345\,
            in2 => \N__43858\,
            in3 => \N__35309\,
            lcout => rand_setpoint_17,
            ltout => OPEN,
            carryin => n16428,
            carryout => n16429,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i18_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35289\,
            in2 => \N__39505\,
            in3 => \N__35264\,
            lcout => rand_setpoint_18,
            ltout => OPEN,
            carryin => n16429,
            carryout => n16430,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i19_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35249\,
            in2 => \N__40765\,
            in3 => \N__35213\,
            lcout => rand_setpoint_19,
            ltout => OPEN,
            carryin => n16430,
            carryout => n16431,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i20_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36144\,
            in2 => \N__40615\,
            in3 => \N__36107\,
            lcout => rand_setpoint_20,
            ltout => OPEN,
            carryin => n16431,
            carryout => n16432,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i21_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43879\,
            in2 => \N__36098\,
            in3 => \N__36047\,
            lcout => rand_setpoint_21,
            ltout => OPEN,
            carryin => n16432,
            carryout => n16433,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i22_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38227\,
            in2 => \N__36034\,
            in3 => \N__36008\,
            lcout => rand_setpoint_22,
            ltout => OPEN,
            carryin => n16433,
            carryout => n16434,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i23_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35991\,
            in2 => \N__41881\,
            in3 => \N__35954\,
            lcout => rand_setpoint_23,
            ltout => OPEN,
            carryin => n16434,
            carryout => n16435,
            clk => \N__50404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i24_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35939\,
            in2 => \N__38249\,
            in3 => \N__35891\,
            lcout => rand_setpoint_24,
            ltout => OPEN,
            carryin => \bfn_9_32_0_\,
            carryout => n16436,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i25_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35867\,
            in2 => \N__38176\,
            in3 => \N__35831\,
            lcout => rand_setpoint_25,
            ltout => OPEN,
            carryin => n16436,
            carryout => n16437,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i26_LC_9_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35802\,
            in2 => \N__39463\,
            in3 => \N__35777\,
            lcout => rand_setpoint_26,
            ltout => OPEN,
            carryin => n16437,
            carryout => n16438,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i27_LC_9_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35759\,
            in2 => \N__38282\,
            in3 => \N__35720\,
            lcout => rand_setpoint_27,
            ltout => OPEN,
            carryin => n16438,
            carryout => n16439,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i28_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36458\,
            in2 => \N__41587\,
            in3 => \N__36413\,
            lcout => rand_setpoint_28,
            ltout => OPEN,
            carryin => n16439,
            carryout => n16440,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i29_LC_9_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38264\,
            in2 => \N__36399\,
            in3 => \N__36359\,
            lcout => rand_setpoint_29,
            ltout => OPEN,
            carryin => n16440,
            carryout => n16441,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i30_LC_9_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38155\,
            in2 => \N__36353\,
            in3 => \N__36311\,
            lcout => rand_setpoint_30,
            ltout => OPEN,
            carryin => n16441,
            carryout => n16442,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2270__i31_LC_9_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36297\,
            in1 => \N__38140\,
            in2 => \_gnd_net_\,
            in3 => \N__36263\,
            lcout => rand_setpoint_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45340\,
            in1 => \N__37604\,
            in2 => \_gnd_net_\,
            in3 => \N__36260\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37417\,
            in1 => \N__48683\,
            in2 => \_gnd_net_\,
            in3 => \N__38690\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i54_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36177\,
            in1 => \N__36224\,
            in2 => \_gnd_net_\,
            in3 => \N__45202\,
            lcout => data_in_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i124_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45200\,
            in1 => \N__37106\,
            in2 => \_gnd_net_\,
            in3 => \N__37087\,
            lcout => data_in_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i50_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37015\,
            in1 => \N__39918\,
            in2 => \_gnd_net_\,
            in3 => \N__45201\,
            lcout => \c0.data_in_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i58_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37043\,
            in1 => \N__45198\,
            in2 => \_gnd_net_\,
            in3 => \N__37008\,
            lcout => \c0.data_in_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i84_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36982\,
            in1 => \N__38570\,
            in2 => \_gnd_net_\,
            in3 => \N__45199\,
            lcout => data_in_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i48_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45197\,
            in1 => \N__36947\,
            in2 => \_gnd_net_\,
            in3 => \N__36902\,
            lcout => data_in_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_844_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36858\,
            in2 => \_gnd_net_\,
            in3 => \N__36832\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i89_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38843\,
            in1 => \N__45208\,
            in2 => \_gnd_net_\,
            in3 => \N__36778\,
            lcout => data_in_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4723_2_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__40214\,
            in1 => \N__40160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n7086,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i122_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36754\,
            in1 => \N__45206\,
            in2 => \_gnd_net_\,
            in3 => \N__38972\,
            lcout => data_in_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_976_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36729\,
            in1 => \N__36690\,
            in2 => \N__36624\,
            in3 => \N__36580\,
            lcout => \c0.n8989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i75_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45205\,
            in1 => \N__36492\,
            in2 => \_gnd_net_\,
            in3 => \N__36523\,
            lcout => data_in_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i152_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37132\,
            in1 => \N__45207\,
            in2 => \_gnd_net_\,
            in3 => \N__37067\,
            lcout => data_in_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i168_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44948\,
            in1 => \N__37121\,
            in2 => \_gnd_net_\,
            in3 => \N__37075\,
            lcout => data_in_20_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i132_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45164\,
            in1 => \N__37102\,
            in2 => \_gnd_net_\,
            in3 => \N__38672\,
            lcout => data_in_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__7__3566_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__46412\,
            in1 => \N__46880\,
            in2 => \N__47143\,
            in3 => \N__47297\,
            lcout => \data_out_5__7__N_931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i116_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44947\,
            in1 => \N__38713\,
            in2 => \_gnd_net_\,
            in3 => \N__37091\,
            lcout => data_in_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i160_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37076\,
            in1 => \N__44949\,
            in2 => \_gnd_net_\,
            in3 => \N__37066\,
            lcout => data_in_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__37396\,
            in1 => \N__37286\,
            in2 => \N__38927\,
            in3 => \N__37055\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001010"
        )
    port map (
            in0 => \N__37049\,
            in1 => \N__40404\,
            in2 => \N__40376\,
            in3 => \N__40221\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37274\,
            in1 => \N__48674\,
            in2 => \_gnd_net_\,
            in3 => \N__38639\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15317_2_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37441\,
            in2 => \_gnd_net_\,
            in3 => \N__38943\,
            lcout => n17767,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__39125\,
            in1 => \N__37402\,
            in2 => \_gnd_net_\,
            in3 => \N__38918\,
            lcout => \c0.tx.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__48614\,
            in1 => \N__37273\,
            in2 => \N__37403\,
            in3 => \N__39124\,
            lcout => n18462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_4_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37252\,
            in1 => \N__37320\,
            in2 => \N__40222\,
            in3 => \N__37209\,
            lcout => n12_adj_2618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11594214_i1_3_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39077\,
            in1 => \_gnd_net_\,
            in2 => \N__38926\,
            in3 => \N__38807\,
            lcout => OPEN,
            ltout => \n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010101"
        )
    port map (
            in0 => \N__40206\,
            in1 => \_gnd_net_\,
            in2 => \N__37181\,
            in3 => \N__40146\,
            lcout => OPEN,
            ltout => \n3_adj_2650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37144\,
            in2 => \N__37178\,
            in3 => \N__40346\,
            lcout => tx_o_adj_2584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_831_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46148\,
            in2 => \_gnd_net_\,
            in3 => \N__41480\,
            lcout => \c0.n9087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_881_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44489\,
            in1 => \N__43274\,
            in2 => \_gnd_net_\,
            in3 => \N__43332\,
            lcout => \c0.n17556\,
            ltout => \c0.n17556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__3__3522_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46149\,
            in1 => \N__37784\,
            in2 => \N__37664\,
            in3 => \N__43532\,
            lcout => \c0.data_out_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50360\,
            ce => \N__46034\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1012_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__37656\,
            in1 => \N__37608\,
            in2 => \N__37574\,
            in3 => \N__37519\,
            lcout => \c0.n16_adj_2513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i137_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37457\,
            in1 => \N__45111\,
            in2 => \_gnd_net_\,
            in3 => \N__39019\,
            lcout => data_in_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7381_2_lut_4_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__37398\,
            in1 => \N__38906\,
            in2 => \N__40133\,
            in3 => \N__39107\,
            lcout => n9796,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_15992_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__37418\,
            in1 => \N__37397\,
            in2 => \N__39123\,
            in3 => \N__39052\,
            lcout => n18438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__40103\,
            in1 => \N__40290\,
            in2 => \_gnd_net_\,
            in3 => \N__37364\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40291\,
            in1 => \N__37334\,
            in2 => \_gnd_net_\,
            in3 => \N__37319\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__40107\,
            in1 => \N__40414\,
            in2 => \N__40240\,
            in3 => \N__40292\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46366\,
            in1 => \N__39485\,
            in2 => \_gnd_net_\,
            in3 => \N__48314\,
            lcout => \c0.n5_adj_2499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__40108\,
            in1 => \N__40415\,
            in2 => \N__40241\,
            in3 => \N__40293\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1072_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40793\,
            in1 => \N__49706\,
            in2 => \_gnd_net_\,
            in3 => \N__43649\,
            lcout => \c0.n6_adj_2448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i143_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37763\,
            in1 => \N__44792\,
            in2 => \_gnd_net_\,
            in3 => \N__37804\,
            lcout => data_in_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i151_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44791\,
            in1 => \N__37762\,
            in2 => \_gnd_net_\,
            in3 => \N__37775\,
            lcout => data_in_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i162_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37753\,
            in1 => \_gnd_net_\,
            in2 => \N__44968\,
            in3 => \N__39041\,
            lcout => data_in_20_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__2__3531_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46041\,
            in1 => \N__37739\,
            in2 => \_gnd_net_\,
            in3 => \N__43328\,
            lcout => data_out_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i158_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37691\,
            in1 => \N__44866\,
            in2 => \_gnd_net_\,
            in3 => \N__37717\,
            lcout => data_in_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i166_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44865\,
            in1 => \N__37706\,
            in2 => \_gnd_net_\,
            in3 => \N__37690\,
            lcout => data_in_20_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__37682\,
            in1 => \N__48110\,
            in2 => \N__37673\,
            in3 => \N__47984\,
            lcout => \c0.n18498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40701\,
            in1 => \N__44141\,
            in2 => \_gnd_net_\,
            in3 => \N__48425\,
            lcout => OPEN,
            ltout => \c0.n2_adj_2487_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18498_bdd_4_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__41336\,
            in1 => \N__37961\,
            in2 => \N__37955\,
            in3 => \N__48111\,
            lcout => \c0.n18501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_104_i4_2_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39230\,
            in2 => \_gnd_net_\,
            in3 => \N__39286\,
            lcout => n4_adj_2649,
            ltout => \n4_adj_2649_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__37834\,
            in1 => \N__37945\,
            in2 => \N__37922\,
            in3 => \N__37915\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__0__3597_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__47561\,
            in1 => \N__47400\,
            in2 => \N__46879\,
            in3 => \N__47079\,
            lcout => data_out_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i161_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37838\,
            in1 => \N__44890\,
            in2 => \_gnd_net_\,
            in3 => \N__37819\,
            lcout => data_in_20_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i135_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37808\,
            in1 => \_gnd_net_\,
            in2 => \N__45112\,
            in3 => \N__37792\,
            lcout => data_in_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i127_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44888\,
            in1 => \N__38200\,
            in2 => \_gnd_net_\,
            in3 => \N__37793\,
            lcout => data_in_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__3__3594_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001110"
        )
    port map (
            in0 => \N__47399\,
            in1 => \N__47670\,
            in2 => \N__47111\,
            in3 => \N__46793\,
            lcout => data_out_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__4__3529_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46033\,
            in1 => \N__38215\,
            in2 => \_gnd_net_\,
            in3 => \N__49603\,
            lcout => data_out_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i119_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38201\,
            in1 => \N__44889\,
            in2 => \_gnd_net_\,
            in3 => \N__44551\,
            lcout => data_in_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__3__3538_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__47448\,
            in1 => \N__45677\,
            in2 => \N__46917\,
            in3 => \N__38191\,
            lcout => \c0.data_out_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50399\,
            ce => \N__44192\,
            sr => \_gnd_net_\
        );

    \c0.i15710_2_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47445\,
            lcout => \c0.n17962\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15722_2_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38159\,
            lcout => \c0.n17972\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15723_2_lut_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38141\,
            in2 => \_gnd_net_\,
            in3 => \N__47446\,
            lcout => \c0.n17974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15760_2_lut_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47444\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38125\,
            lcout => \c0.n17921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i130_3_lut_4_lut_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__38111\,
            in1 => \N__38060\,
            in2 => \N__38021\,
            in3 => \N__38000\,
            lcout => \c0.rx.r_SM_Main_2_N_2380_2\,
            ltout => \c0.rx.r_SM_Main_2_N_2380_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15739_2_lut_3_lut_4_lut_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40452\,
            in1 => \N__39236\,
            in2 => \N__37964\,
            in3 => \N__39300\,
            lcout => OPEN,
            ltout => \c0.rx.n18000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111000000"
        )
    port map (
            in0 => \N__39631\,
            in1 => \N__39711\,
            in2 => \N__38300\,
            in3 => \N__39590\,
            lcout => \c0.rx.n18594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15874_4_lut_4_lut_4_lut_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47106\,
            in2 => \_gnd_net_\,
            in3 => \N__47439\,
            lcout => n9519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15714_2_lut_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38281\,
            lcout => OPEN,
            ltout => \c0.n17966_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__3__3554_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__40792\,
            in1 => \N__49443\,
            in2 => \N__38267\,
            in3 => \N__46891\,
            lcout => \c0.data_out_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50405\,
            ce => \N__46516\,
            sr => \_gnd_net_\
        );

    \c0.i15717_2_lut_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38263\,
            lcout => OPEN,
            ltout => \c0.n17970_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__5__3552_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111100100"
        )
    port map (
            in0 => \N__46892\,
            in1 => \N__49444\,
            in2 => \N__38252\,
            in3 => \N__49853\,
            lcout => \c0.data_out_7__5__N_543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50405\,
            ce => \N__46516\,
            sr => \_gnd_net_\
        );

    \c0.i15705_2_lut_LC_10_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38248\,
            lcout => OPEN,
            ltout => \c0.n17957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__0__3557_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011101"
        )
    port map (
            in0 => \N__47771\,
            in1 => \N__49442\,
            in2 => \N__38234\,
            in3 => \N__46890\,
            lcout => \c0.data_out_6__3__N_788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50405\,
            ce => \N__46516\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6__3543_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__47443\,
            in1 => \N__40631\,
            in2 => \N__38231\,
            in3 => \N__46893\,
            lcout => \c0.data_out_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50405\,
            ce => \N__46516\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i147_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44649\,
            in1 => \N__38413\,
            in2 => \_gnd_net_\,
            in3 => \N__38474\,
            lcout => data_in_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i149_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38432\,
            in1 => \N__44652\,
            in2 => \_gnd_net_\,
            in3 => \N__38422\,
            lcout => data_in_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i157_LC_10_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44651\,
            in1 => \N__38453\,
            in2 => \_gnd_net_\,
            in3 => \N__38431\,
            lcout => data_in_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i141_LC_10_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44648\,
            in1 => \N__38536\,
            in2 => \_gnd_net_\,
            in3 => \N__38423\,
            lcout => data_in_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i139_LC_10_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38414\,
            in1 => \N__44650\,
            in2 => \_gnd_net_\,
            in3 => \N__38398\,
            lcout => data_in_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i69_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38347\,
            in1 => \N__45212\,
            in2 => \_gnd_net_\,
            in3 => \N__38364\,
            lcout => data_in_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i77_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38326\,
            in1 => \_gnd_net_\,
            in2 => \N__45342\,
            in3 => \N__38346\,
            lcout => data_in_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i85_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__45213\,
            in2 => \_gnd_net_\,
            in3 => \N__38325\,
            lcout => data_in_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i93_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38597\,
            in1 => \_gnd_net_\,
            in2 => \N__45343\,
            in3 => \N__38308\,
            lcout => data_in_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i101_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38588\,
            in1 => \N__45210\,
            in2 => \_gnd_net_\,
            in3 => \N__38596\,
            lcout => data_in_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i109_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38579\,
            in1 => \_gnd_net_\,
            in2 => \N__45341\,
            in3 => \N__38587\,
            lcout => data_in_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i117_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38558\,
            in1 => \N__45211\,
            in2 => \_gnd_net_\,
            in3 => \N__38578\,
            lcout => data_in_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i92_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45196\,
            in1 => \N__38569\,
            in2 => \_gnd_net_\,
            in3 => \N__38828\,
            lcout => data_in_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i125_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45209\,
            in1 => \N__38557\,
            in2 => \_gnd_net_\,
            in3 => \N__38525\,
            lcout => data_in_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i133_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45158\,
            in1 => \N__38524\,
            in2 => \_gnd_net_\,
            in3 => \N__38546\,
            lcout => data_in_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i34_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39885\,
            in1 => \N__38493\,
            in2 => \_gnd_net_\,
            in3 => \N__45159\,
            lcout => data_in_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15747_2_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41797\,
            in2 => \_gnd_net_\,
            in3 => \N__48397\,
            lcout => OPEN,
            ltout => \c0.n18089_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18426_bdd_4_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__43973\,
            in1 => \N__38678\,
            in2 => \N__38477\,
            in3 => \N__48109\,
            lcout => OPEN,
            ltout => \c0.n18429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11402_4_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__44063\,
            in1 => \N__48845\,
            in2 => \N__38693\,
            in3 => \N__48754\,
            lcout => \tx_data_7_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15753_2_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45662\,
            in2 => \_gnd_net_\,
            in3 => \N__48396\,
            lcout => OPEN,
            ltout => \c0.n18017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_16021_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__39395\,
            in1 => \N__48108\,
            in2 => \N__38681\,
            in3 => \N__47981\,
            lcout => \c0.n18426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i140_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44950\,
            in1 => \N__38671\,
            in2 => \_gnd_net_\,
            in3 => \N__38852\,
            lcout => data_in_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15935_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__40874\,
            in1 => \N__48080\,
            in2 => \N__38660\,
            in3 => \N__47982\,
            lcout => OPEN,
            ltout => \c0.n18378_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18378_bdd_4_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48081\,
            in1 => \N__41351\,
            in2 => \N__38645\,
            in3 => \N__40655\,
            lcout => OPEN,
            ltout => \c0.n18381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11425_4_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__43157\,
            in1 => \N__48844\,
            in2 => \N__38642\,
            in3 => \N__48759\,
            lcout => \tx_data_2_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i156_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44952\,
            in1 => \N__38633\,
            in2 => \_gnd_net_\,
            in3 => \N__38860\,
            lcout => data_in_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i110_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45204\,
            in1 => \N__38608\,
            in2 => \_gnd_net_\,
            in3 => \N__39335\,
            lcout => data_in_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i148_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44951\,
            in1 => \N__38851\,
            in2 => \_gnd_net_\,
            in3 => \N__38861\,
            lcout => data_in_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i97_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45051\,
            in1 => \N__38842\,
            in2 => \_gnd_net_\,
            in3 => \N__39068\,
            lcout => data_in_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i100_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38824\,
            in1 => \N__45052\,
            in2 => \_gnd_net_\,
            in3 => \N__38702\,
            lcout => data_in_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n18462_bdd_4_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__42206\,
            in1 => \N__39368\,
            in2 => \N__39137\,
            in3 => \N__38813\,
            lcout => n18465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i71_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__38743\,
            in2 => \_gnd_net_\,
            in3 => \N__45053\,
            lcout => data_in_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i126_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45050\,
            in1 => \N__39349\,
            in2 => \_gnd_net_\,
            in3 => \N__38732\,
            lcout => data_in_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i9_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__42438\,
            in1 => \N__40019\,
            in2 => \N__41936\,
            in3 => \N__42579\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i6_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__41964\,
            in1 => \N__39941\,
            in2 => \N__42581\,
            in3 => \N__42437\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i108_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45054\,
            in1 => \N__38701\,
            in2 => \_gnd_net_\,
            in3 => \N__38714\,
            lcout => data_in_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i138_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45115\,
            in1 => \N__38983\,
            in2 => \_gnd_net_\,
            in3 => \N__38873\,
            lcout => data_in_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_924_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__41900\,
            in2 => \_gnd_net_\,
            in3 => \N__38996\,
            lcout => \c0.n17349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15288_2_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41018\,
            in2 => \_gnd_net_\,
            in3 => \N__41048\,
            lcout => OPEN,
            ltout => \n17737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_1137_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40981\,
            in1 => \N__42884\,
            in2 => \N__38999\,
            in3 => \N__41159\,
            lcout => n17312,
            ltout => \n17312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_1144_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38990\,
            in3 => \N__42263\,
            lcout => n14_adj_2615,
            ltout => \n14_adj_2615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__42697\,
            in1 => \N__41320\,
            in2 => \N__38987\,
            in3 => \N__41306\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43034\,
            in1 => \N__42696\,
            in2 => \N__48164\,
            in3 => \N__42729\,
            lcout => byte_transmit_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i130_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38984\,
            in1 => \N__45056\,
            in2 => \_gnd_net_\,
            in3 => \N__38965\,
            lcout => data_in_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001000100"
        )
    port map (
            in0 => \N__38905\,
            in1 => \N__40154\,
            in2 => \_gnd_net_\,
            in3 => \N__38954\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i146_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45113\,
            in1 => \N__38872\,
            in2 => \_gnd_net_\,
            in3 => \N__39029\,
            lcout => data_in_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n18438_bdd_4_lut_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__39143\,
            in1 => \N__43181\,
            in2 => \N__42797\,
            in3 => \N__39130\,
            lcout => n18441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i105_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39064\,
            in1 => \N__45055\,
            in2 => \_gnd_net_\,
            in3 => \N__39179\,
            lcout => data_in_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48642\,
            in1 => \N__39053\,
            in2 => \_gnd_net_\,
            in3 => \N__40514\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i154_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45114\,
            in1 => \N__39040\,
            in2 => \_gnd_net_\,
            in3 => \N__39028\,
            lcout => data_in_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__43073\,
            in1 => \N__48377\,
            in2 => \N__42708\,
            in3 => \N__40054\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i121_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39008\,
            in1 => \N__44946\,
            in2 => \_gnd_net_\,
            in3 => \N__39190\,
            lcout => data_in_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15801_2_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45713\,
            in2 => \_gnd_net_\,
            in3 => \N__48306\,
            lcout => \c0.n17937\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__39290\,
            in1 => \N__39320\,
            in2 => \N__40502\,
            in3 => \N__40472\,
            lcout => \r_Bit_Index_2_adj_2625\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i129_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44945\,
            in1 => \N__39007\,
            in2 => \_gnd_net_\,
            in3 => \N__39020\,
            lcout => data_in_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11225_4_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__39377\,
            in1 => \N__48837\,
            in2 => \N__48761\,
            in3 => \N__43202\,
            lcout => OPEN,
            ltout => \tx_data_0_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48648\,
            in2 => \N__39371\,
            in3 => \N__39367\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i118_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44767\,
            in1 => \N__39353\,
            in2 => \_gnd_net_\,
            in3 => \N__39331\,
            lcout => data_in_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_868_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40741\,
            in1 => \N__48592\,
            in2 => \_gnd_net_\,
            in3 => \N__43940\,
            lcout => \c0.n17465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2428_2_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40444\,
            in2 => \_gnd_net_\,
            in3 => \N__39228\,
            lcout => n4958,
            ltout => \n4958_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i7504_3_lut_4_lut_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011001100"
        )
    port map (
            in0 => \N__39285\,
            in1 => \N__40496\,
            in2 => \N__39251\,
            in3 => \N__39718\,
            lcout => n9920,
            ltout => \n9920_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__40497\,
            in1 => \N__40445\,
            in2 => \N__39248\,
            in3 => \N__39229\,
            lcout => \r_Bit_Index_1_adj_2626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i113_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44902\,
            in1 => \N__39175\,
            in2 => \_gnd_net_\,
            in3 => \N__39194\,
            lcout => data_in_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__1__3532_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46031\,
            in1 => \_gnd_net_\,
            in2 => \N__39164\,
            in3 => \N__44481\,
            lcout => data_out_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__0__3533_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47826\,
            in1 => \N__46030\,
            in2 => \_gnd_net_\,
            in3 => \N__39437\,
            lcout => data_out_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1062_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44474\,
            in1 => \N__47825\,
            in2 => \_gnd_net_\,
            in3 => \N__39484\,
            lcout => \c0.n8953\,
            ltout => \c0.n8953_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1044_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41657\,
            in2 => \N__39419\,
            in3 => \N__45597\,
            lcout => \c0.n17626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__5__3528_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46032\,
            in1 => \N__39416\,
            in2 => \_gnd_net_\,
            in3 => \N__49697\,
            lcout => data_out_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48394\,
            in1 => \N__43527\,
            in2 => \_gnd_net_\,
            in3 => \N__47800\,
            lcout => \c0.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_882_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40693\,
            in1 => \N__47669\,
            in2 => \_gnd_net_\,
            in3 => \N__40740\,
            lcout => \c0.n17400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__6__3551_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001011"
        )
    port map (
            in0 => \N__49446\,
            in1 => \N__40643\,
            in2 => \N__46916\,
            in3 => \N__39383\,
            lcout => \c0.data_out_7__6__N_530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50406\,
            ce => \N__46546\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__7__I_0_3654_2_lut_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48569\,
            in2 => \_gnd_net_\,
            in3 => \N__45653\,
            lcout => \c0.data_out_7__1__N_626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1003_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45914\,
            lcout => \c0.n17665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__39773\,
            in1 => \N__39641\,
            in2 => \N__39719\,
            in3 => \N__39588\,
            lcout => \c0.rx.n9553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_4_lut_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__39587\,
            in1 => \N__39772\,
            in2 => \N__39650\,
            in3 => \N__39713\,
            lcout => n9646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15891_2_lut_3_lut_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__39589\,
            in1 => \N__39774\,
            in2 => \_gnd_net_\,
            in3 => \N__39712\,
            lcout => \c0.rx.n17351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_815_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39710\,
            in2 => \_gnd_net_\,
            in3 => \N__39586\,
            lcout => \c0.rx.n17376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2__I_596_2_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43803\,
            lcout => \c0.data_out_6__2__N_803\,
            ltout => \c0.data_out_6__2__N_803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_832_i1_4_lut_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__49790\,
            in1 => \N__43132\,
            in2 => \N__39509\,
            in3 => \N__49447\,
            lcout => OPEN,
            ltout => \c0.n2216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2__3547_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47415\,
            in1 => \N__39506\,
            in2 => \N__39488\,
            in3 => \N__46889\,
            lcout => \c0.data_out_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50412\,
            ce => \N__46538\,
            sr => \_gnd_net_\
        );

    \c0.i15712_2_lut_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39467\,
            in2 => \_gnd_net_\,
            in3 => \N__47414\,
            lcout => OPEN,
            ltout => \c0.n17964_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2__3555_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__49448\,
            in1 => \N__39446\,
            in2 => \N__39440\,
            in3 => \N__46888\,
            lcout => \c0.data_out_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50412\,
            ce => \N__46538\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_855_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41237\,
            lcout => \c0.n17525\,
            ltout => \c0.n17525_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_856_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40702\,
            in1 => \N__47644\,
            in2 => \N__39791\,
            in3 => \N__47579\,
            lcout => \c0.n17644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_904_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46954\,
            in1 => \N__49846\,
            in2 => \_gnd_net_\,
            in3 => \N__43561\,
            lcout => \c0.n6_adj_2467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__4__3585_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__49450\,
            in1 => \N__49867\,
            in2 => \N__46502\,
            in3 => \N__46884\,
            lcout => \c0.data_out_5__5__N_950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__2__3587_LC_11_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__46882\,
            in1 => \N__46484\,
            in2 => \N__43770\,
            in3 => \N__49451\,
            lcout => data_out_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__7__3582_LC_11_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110010"
        )
    port map (
            in0 => \N__47453\,
            in1 => \N__46883\,
            in2 => \N__41793\,
            in3 => \N__47136\,
            lcout => data_out_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1061_LC_11_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__49615\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49651\,
            lcout => \c0.n8970\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__4__3569_LC_11_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__47137\,
            in1 => \N__41244\,
            in2 => \N__47498\,
            in3 => \N__47454\,
            lcout => data_out_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__5__3592_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__47452\,
            in1 => \N__47135\,
            in2 => \N__43946\,
            in3 => \N__47494\,
            lcout => data_out_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__39788\,
            in1 => \N__39779\,
            in2 => \N__44768\,
            in3 => \N__39717\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i42_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45293\,
            in1 => \N__39878\,
            in2 => \_gnd_net_\,
            in3 => \N__39931\,
            lcout => data_in_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i87_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45157\,
            in1 => \N__39812\,
            in2 => \_gnd_net_\,
            in3 => \N__39834\,
            lcout => data_in_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i43_4_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111010"
        )
    port map (
            in0 => \N__46795\,
            in1 => \N__40928\,
            in2 => \N__49308\,
            in3 => \N__42155\,
            lcout => \c0.n25_adj_2517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__49244\,
            in1 => \N__46794\,
            in2 => \_gnd_net_\,
            in3 => \N__47342\,
            lcout => n9631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i8_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40031\,
            in1 => \N__42329\,
            in2 => \_gnd_net_\,
            in3 => \N__42429\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i95_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45203\,
            in1 => \N__39811\,
            in2 => \_gnd_net_\,
            in3 => \N__40943\,
            lcout => data_in_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15306_4_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42300\,
            in1 => \N__42083\,
            in2 => \N__42334\,
            in3 => \N__41738\,
            lcout => \c0.n17755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i10_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__41739\,
            in1 => \N__42562\,
            in2 => \N__40010\,
            in3 => \N__42427\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i3_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__42428\,
            in1 => \N__41123\,
            in2 => \N__39959\,
            in3 => \N__42569\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1021_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__42656\,
            in1 => \N__39983\,
            in2 => \_gnd_net_\,
            in3 => \N__47283\,
            lcout => \c0.n1314\,
            ltout => \c0.n1314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i2_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__42561\,
            in1 => \N__39968\,
            in2 => \N__39977\,
            in3 => \N__41086\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_2_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41043\,
            in2 => \_gnd_net_\,
            in3 => \N__39974\,
            lcout => \c0.n7275\,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \c0.n16305\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_3_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41102\,
            in2 => \_gnd_net_\,
            in3 => \N__39971\,
            lcout => \c0.n7274\,
            ltout => OPEN,
            carryin => \c0.n16305\,
            carryout => \c0.n16306\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_4_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41085\,
            in2 => \_gnd_net_\,
            in3 => \N__39962\,
            lcout => \c0.n7273\,
            ltout => OPEN,
            carryin => \c0.n16306\,
            carryout => \c0.n16307\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_5_lut_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41121\,
            in2 => \_gnd_net_\,
            in3 => \N__39950\,
            lcout => \c0.n7272\,
            ltout => OPEN,
            carryin => \c0.n16307\,
            carryout => \c0.n16308\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_6_lut_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41065\,
            in2 => \_gnd_net_\,
            in3 => \N__39947\,
            lcout => \c0.n7271\,
            ltout => OPEN,
            carryin => \c0.n16308\,
            carryout => \c0.n16309\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_7_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42555\,
            in1 => \_gnd_net_\,
            in2 => \N__42302\,
            in3 => \N__39944\,
            lcout => \c0.n18012\,
            ltout => OPEN,
            carryin => \c0.n16309\,
            carryout => \c0.n16310\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_8_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41960\,
            in2 => \_gnd_net_\,
            in3 => \N__39935\,
            lcout => \c0.n7269\,
            ltout => OPEN,
            carryin => \c0.n16310\,
            carryout => \c0.n16311\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_9_lut_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42380\,
            in2 => \_gnd_net_\,
            in3 => \N__40034\,
            lcout => \c0.n7268\,
            ltout => OPEN,
            carryin => \c0.n16311\,
            carryout => \c0.n16312\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_10_lut_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42575\,
            in1 => \N__42333\,
            in2 => \_gnd_net_\,
            in3 => \N__40022\,
            lcout => \c0.n18011\,
            ltout => OPEN,
            carryin => \bfn_12_25_0_\,
            carryout => \c0.n16313\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_11_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41927\,
            in2 => \_gnd_net_\,
            in3 => \N__40013\,
            lcout => \c0.n7266\,
            ltout => OPEN,
            carryin => \c0.n16313\,
            carryout => \c0.n16314\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_12_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41743\,
            in2 => \_gnd_net_\,
            in3 => \N__39998\,
            lcout => \c0.n7265\,
            ltout => OPEN,
            carryin => \c0.n16314\,
            carryout => \c0.n16315\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_13_lut_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42355\,
            in2 => \_gnd_net_\,
            in3 => \N__39995\,
            lcout => \c0.n7264\,
            ltout => OPEN,
            carryin => \c0.n16315\,
            carryout => \c0.n16316\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_14_lut_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42574\,
            in1 => \N__42082\,
            in2 => \_gnd_net_\,
            in3 => \N__39992\,
            lcout => \c0.n18009\,
            ltout => OPEN,
            carryin => \c0.n16316\,
            carryout => \c0.n16317\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_15_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__42551\,
            in1 => \N__41009\,
            in2 => \_gnd_net_\,
            in3 => \N__39989\,
            lcout => \c0.n18008\,
            ltout => OPEN,
            carryin => \c0.n16317\,
            carryout => \c0.n16318\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3777_16_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__40982\,
            in1 => \N__42552\,
            in2 => \_gnd_net_\,
            in3 => \N__39986\,
            lcout => \c0.n18105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__41282\,
            in1 => \N__42730\,
            in2 => \N__42692\,
            in3 => \N__41267\,
            lcout => byte_transmit_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15852_3_lut_4_lut_4_lut_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001110000000"
        )
    port map (
            in0 => \N__40413\,
            in1 => \N__40239\,
            in2 => \N__40162\,
            in3 => \N__42984\,
            lcout => OPEN,
            ltout => \n4_adj_2653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111010"
        )
    port map (
            in0 => \N__42914\,
            in1 => \N__40153\,
            in2 => \N__40379\,
            in3 => \N__40338\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i241_2_lut_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40061\,
            in2 => \_gnd_net_\,
            in3 => \N__42913\,
            lcout => \c0.n251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_4_lut_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40337\,
            in1 => \N__40238\,
            in2 => \N__40161\,
            in3 => \N__42983\,
            lcout => n7734,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_3508_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__43052\,
            in1 => \N__47930\,
            in2 => \N__42707\,
            in3 => \N__40055\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46950\,
            in1 => \N__40847\,
            in2 => \_gnd_net_\,
            in3 => \N__48376\,
            lcout => \c0.n2_adj_2476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15940_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__40043\,
            in1 => \N__48106\,
            in2 => \N__47969\,
            in3 => \N__41384\,
            lcout => OPEN,
            ltout => \c0.n18390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18390_bdd_4_lut_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48107\,
            in1 => \N__41360\,
            in2 => \N__40037\,
            in3 => \N__40508\,
            lcout => OPEN,
            ltout => \c0.n18393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11421_4_lut_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__45524\,
            in1 => \N__48815\,
            in2 => \N__40517\,
            in3 => \N__48755\,
            lcout => \tx_data_3_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15744_2_lut_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43408\,
            lcout => \c0.n18095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41656\,
            in1 => \N__43300\,
            in2 => \_gnd_net_\,
            in3 => \N__48312\,
            lcout => \c0.n5_adj_2447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43407\,
            in1 => \N__40728\,
            in2 => \N__40697\,
            in3 => \N__46441\,
            lcout => \c0.n17641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1__I_638_2_lut_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44013\,
            lcout => \c0.data_out_6__1__N_849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__40501\,
            in1 => \N__40451\,
            in2 => \_gnd_net_\,
            in3 => \N__40471\,
            lcout => \r_Bit_Index_0_adj_2627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__0__3581_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100010000"
        )
    port map (
            in0 => \N__47039\,
            in1 => \N__46872\,
            in2 => \N__47465\,
            in3 => \N__40686\,
            lcout => data_out_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_834_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40849\,
            lcout => \c0.n17445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15782_2_lut_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40526\,
            in2 => \_gnd_net_\,
            in3 => \N__48395\,
            lcout => \c0.n18062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__2__3579_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001001110"
        )
    port map (
            in0 => \N__47434\,
            in1 => \N__40729\,
            in2 => \N__46915\,
            in3 => \N__47040\,
            lcout => \data_out_6__6__N_729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__5__3568_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__46949\,
            in1 => \N__46873\,
            in2 => \N__47078\,
            in3 => \N__47435\,
            lcout => data_out_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_895_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47767\,
            in1 => \N__43949\,
            in2 => \N__43421\,
            in3 => \N__40850\,
            lcout => \c0.data_out_6__7__N_675\,
            ltout => \c0.data_out_6__7__N_675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15683_3_lut_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010000010"
        )
    port map (
            in0 => \N__49435\,
            in1 => \N__45658\,
            in2 => \N__40595\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n17928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__7__3534_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47398\,
            in1 => \N__40592\,
            in2 => \N__40571\,
            in3 => \N__46871\,
            lcout => \c0.data_out_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50407\,
            ce => \N__44187\,
            sr => \_gnd_net_\
        );

    \c0.i15763_2_lut_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47397\,
            lcout => OPEN,
            ltout => \c0.n17906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6__3535_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__49383\,
            in1 => \N__40550\,
            in2 => \N__40541\,
            in3 => \N__46870\,
            lcout => \c0.data_out_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50407\,
            ce => \N__44187\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_878_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48198\,
            in1 => \N__47799\,
            in2 => \_gnd_net_\,
            in3 => \N__41821\,
            lcout => \c0.n8950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2__3539_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__46869\,
            in1 => \N__43121\,
            in2 => \N__49449\,
            in3 => \N__40538\,
            lcout => \c0.data_out_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50407\,
            ce => \N__44187\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__6__3511_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43945\,
            in1 => \N__40745\,
            in2 => \N__46219\,
            in3 => \N__48570\,
            lcout => \c0.data_out_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50413\,
            ce => \N__46047\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40743\,
            in1 => \N__41623\,
            in2 => \_gnd_net_\,
            in3 => \N__48460\,
            lcout => \c0.n2_adj_2483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_835_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44268\,
            in2 => \_gnd_net_\,
            in3 => \N__43651\,
            lcout => \c0.n8634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1104_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__49866\,
            in1 => \_gnd_net_\,
            in2 => \N__41254\,
            in3 => \N__41624\,
            lcout => \c0.n17389\,
            ltout => \c0.n17389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1052_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41541\,
            in1 => \N__43562\,
            in2 => \N__40637\,
            in3 => \N__45717\,
            lcout => \c0.n17600\,
            ltout => \c0.n17600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_728_i1_4_lut_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__40744\,
            in1 => \N__43944\,
            in2 => \N__40634\,
            in3 => \N__49417\,
            lcout => \c0.n9658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1060_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43750\,
            in1 => \N__41621\,
            in2 => \N__41546\,
            in3 => \N__44140\,
            lcout => \c0.n17398\,
            ltout => \c0.n17398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_780_i1_4_lut_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__41689\,
            in1 => \N__46382\,
            in2 => \N__40619\,
            in3 => \N__49420\,
            lcout => OPEN,
            ltout => \c0.n2146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4__3545_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47436\,
            in1 => \N__40616\,
            in2 => \N__40598\,
            in3 => \N__46896\,
            lcout => \c0.data_out_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50418\,
            ce => \N__46557\,
            sr => \_gnd_net_\
        );

    \c0.data_out_1__1__3588_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__46894\,
            in1 => \N__49421\,
            in2 => \_gnd_net_\,
            in3 => \N__47437\,
            lcout => \c0.data_out_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50418\,
            ce => \N__46557\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1088_LC_12_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43749\,
            in1 => \N__43796\,
            in2 => \_gnd_net_\,
            in3 => \N__44000\,
            lcout => \c0.data_out_5__3__N_964\,
            ltout => \c0.data_out_5__3__N_964_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1069_LC_12_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43647\,
            in2 => \N__40772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.data_out_6__3__N_785_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_806_i1_4_lut_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__49419\,
            in1 => \N__45749\,
            in2 => \N__40769\,
            in3 => \N__49791\,
            lcout => OPEN,
            ltout => \c0.n2181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3__3546_LC_12_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46895\,
            in1 => \N__40766\,
            in2 => \N__40748\,
            in3 => \N__47438\,
            lcout => \c0.data_out_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50418\,
            ce => \N__46557\,
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6__3591_LC_12_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__49422\,
            in1 => \N__47766\,
            in2 => \N__46918\,
            in3 => \N__46523\,
            lcout => \c0.data_out_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__2__3571_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__47126\,
            in1 => \N__41615\,
            in2 => \N__47461\,
            in3 => \N__47488\,
            lcout => \data_out_5__4__N_959\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1067_LC_12_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40742\,
            in1 => \N__43394\,
            in2 => \N__40703\,
            in3 => \N__41755\,
            lcout => \c0.n17653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3__3578_LC_12_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__46524\,
            in1 => \N__46907\,
            in2 => \N__43409\,
            in3 => \N__49423\,
            lcout => \c0.data_out_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__7__3574_LC_12_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001110"
        )
    port map (
            in0 => \N__47450\,
            in1 => \N__43994\,
            in2 => \N__47141\,
            in3 => \N__46898\,
            lcout => \data_out_6__1__N_850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__5__3576_LC_12_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111110000"
        )
    port map (
            in0 => \N__46897\,
            in1 => \N__47122\,
            in2 => \N__40846\,
            in3 => \N__47451\,
            lcout => \data_out_6__7__N_678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_990_LC_12_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40831\,
            in1 => \N__44128\,
            in2 => \N__44001\,
            in3 => \N__41614\,
            lcout => \c0.n8964\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15704_4_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__47295\,
            in1 => \N__42571\,
            in2 => \N__42893\,
            in3 => \N__42050\,
            lcout => n17958,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_889_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46799\,
            lcout => n2615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1007_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__42888\,
            in1 => \N__42570\,
            in2 => \N__41453\,
            in3 => \N__42049\,
            lcout => n8488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1025_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__43010\,
            in1 => \N__42839\,
            in2 => \N__42892\,
            in3 => \N__42184\,
            lcout => n96,
            ltout => \n96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__49253\,
            in1 => \N__47229\,
            in2 => \N__40814\,
            in3 => \N__42126\,
            lcout => n17709,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_1147_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__46788\,
            in1 => \N__41988\,
            in2 => \_gnd_net_\,
            in3 => \N__42108\,
            lcout => OPEN,
            ltout => \n47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1148_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__49254\,
            in1 => \N__40807\,
            in2 => \N__40811\,
            in3 => \N__42003\,
            lcout => OPEN,
            ltout => \n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i2_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__42004\,
            in1 => \N__40808\,
            in2 => \N__40796\,
            in3 => \N__40907\,
            lcout => \UART_TRANSMITTER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i64_4_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__41989\,
            in1 => \N__46787\,
            in2 => \N__40916\,
            in3 => \N__42142\,
            lcout => n43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i4_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__41066\,
            in1 => \N__42567\,
            in2 => \N__40901\,
            in3 => \N__42430\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__1__3596_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101010"
        )
    port map (
            in0 => \N__47619\,
            in1 => \N__46789\,
            in2 => \N__47127\,
            in3 => \N__47241\,
            lcout => data_out_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i14_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__42431\,
            in1 => \_gnd_net_\,
            in2 => \N__40892\,
            in3 => \N__40974\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i5_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40880\,
            in1 => \N__42301\,
            in2 => \_gnd_net_\,
            in3 => \N__42432\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1001_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__42838\,
            in1 => \N__42185\,
            in2 => \N__42985\,
            in3 => \N__42930\,
            lcout => \c0.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15731_2_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43588\,
            in2 => \_gnd_net_\,
            in3 => \N__48426\,
            lcout => \c0.n17936\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i0_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001111"
        )
    port map (
            in0 => \N__41047\,
            in1 => \N__40865\,
            in2 => \N__42580\,
            in3 => \N__42433\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i1_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__42435\,
            in1 => \N__41101\,
            in2 => \N__40859\,
            in3 => \N__42566\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i13_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41132\,
            in1 => \_gnd_net_\,
            in2 => \N__41011\,
            in3 => \N__42436\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_912_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41122\,
            in1 => \N__41100\,
            in2 => \N__41087\,
            in3 => \N__41064\,
            lcout => \c0.n17387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1042_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42224\,
            in1 => \N__41036\,
            in2 => \N__41010\,
            in3 => \N__40968\,
            lcout => n29,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i11_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__42434\,
            in1 => \N__40952\,
            in2 => \N__40946\,
            in3 => \N__42356\,
            lcout => \c0.delay_counter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i103_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45495\,
            in1 => \N__44540\,
            in2 => \_gnd_net_\,
            in3 => \N__40942\,
            lcout => data_in_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i149_2_lut_3_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__43069\,
            in1 => \N__43051\,
            in2 => \_gnd_net_\,
            in3 => \N__43027\,
            lcout => \c0.n149\,
            ltout => \c0.n149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_915_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__42828\,
            in1 => \_gnd_net_\,
            in2 => \N__40931\,
            in3 => \N__42175\,
            lcout => n119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1019_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__42176\,
            in1 => \N__42870\,
            in2 => \N__42590\,
            in3 => \N__42829\,
            lcout => \c0.n93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1126_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__46627\,
            in1 => \N__47242\,
            in2 => \_gnd_net_\,
            in3 => \N__42240\,
            lcout => n8529,
            ltout => \n8529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_917_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__49255\,
            in1 => \N__43002\,
            in2 => \N__41180\,
            in3 => \N__41174\,
            lcout => \c0.n16450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_905_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41299\,
            in1 => \N__42628\,
            in2 => \N__41210\,
            in3 => \N__41266\,
            lcout => \c0.n8550\,
            ltout => \c0.n8550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_908_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41177\,
            in3 => \N__42827\,
            lcout => n121_adj_2606,
            ltout => \n121_adj_2606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__41423\,
            in1 => \N__41168\,
            in2 => \N__41162\,
            in3 => \N__49256\,
            lcout => n13_adj_2652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_2_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41150\,
            in2 => \N__48398\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_transmit_N_2239_0\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \c0.n16350\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_3_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47890\,
            in2 => \_gnd_net_\,
            in3 => \N__41144\,
            lcout => \c0.tx_transmit_N_2239_1\,
            ltout => OPEN,
            carryin => \c0.n16350\,
            carryout => \c0.n16351\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_4_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48112\,
            in2 => \_gnd_net_\,
            in3 => \N__41141\,
            lcout => \tx_transmit_N_2239_2\,
            ltout => OPEN,
            carryin => \c0.n16351\,
            carryout => \c0.n16352\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_5_lut_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48720\,
            in2 => \_gnd_net_\,
            in3 => \N__41138\,
            lcout => \tx_transmit_N_2239_3\,
            ltout => OPEN,
            carryin => \c0.n16352\,
            carryout => \c0.n16353\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_6_lut_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48804\,
            in2 => \_gnd_net_\,
            in3 => \N__41135\,
            lcout => \tx_transmit_N_2239_4\,
            ltout => OPEN,
            carryin => \c0.n16353\,
            carryout => \c0.n16354\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_7_lut_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41324\,
            in2 => \_gnd_net_\,
            in3 => \N__41288\,
            lcout => \tx_transmit_N_2239_5\,
            ltout => OPEN,
            carryin => \c0.n16354\,
            carryout => \c0.n16355\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_8_lut_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42617\,
            in3 => \N__41285\,
            lcout => \tx_transmit_N_2239_6\,
            ltout => OPEN,
            carryin => \c0.n16355\,
            carryout => \c0.n16356\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_3776_9_lut_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41281\,
            in2 => \_gnd_net_\,
            in3 => \N__41270\,
            lcout => \tx_transmit_N_2239_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15743_2_lut_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48401\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41255\,
            lcout => OPEN,
            ltout => \c0.n18093_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18396_bdd_4_lut_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__41366\,
            in1 => \N__41186\,
            in2 => \N__41216\,
            in3 => \N__48133\,
            lcout => OPEN,
            ltout => \c0.n18399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11416_4_lut_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__41390\,
            in1 => \N__48811\,
            in2 => \N__41213\,
            in3 => \N__48724\,
            lcout => \tx_data_4_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__42749\,
            in1 => \N__42706\,
            in2 => \N__48833\,
            in3 => \N__41209\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15689_2_lut_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43231\,
            lcout => OPEN,
            ltout => \c0.n17941_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15945_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__41195\,
            in1 => \N__48129\,
            in2 => \N__41189\,
            in3 => \N__47956\,
            lcout => \c0.n18396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15796_4_lut_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__47957\,
            in1 => \N__41372\,
            in2 => \N__48156\,
            in3 => \N__44447\,
            lcout => \c0.n18068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46086\,
            in1 => \N__43269\,
            in2 => \_gnd_net_\,
            in3 => \N__48400\,
            lcout => \c0.n5_adj_2490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__4__3513_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46087\,
            in1 => \N__41672\,
            in2 => \N__46365\,
            in3 => \N__43461\,
            lcout => \c0.data_out_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50408\,
            ce => \N__46029\,
            sr => \_gnd_net_\
        );

    \c0.i15822_2_lut_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41378\,
            lcout => \c0.n18067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15742_2_lut_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49874\,
            in2 => \_gnd_net_\,
            in3 => \N__48411\,
            lcout => \c0.n18092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15794_2_lut_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__47696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48412\,
            lcout => \c0.n18094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15798_2_lut_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43772\,
            lcout => \c0.n18096\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15815_2_lut_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47577\,
            in2 => \_gnd_net_\,
            in3 => \N__48415\,
            lcout => \c0.n18088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15875_2_lut_3_lut_4_lut_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__46696\,
            in1 => \N__49322\,
            in2 => \N__47077\,
            in3 => \N__47300\,
            lcout => \c0.n9518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11502_2_lut_3_lut_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__47299\,
            in1 => \N__49324\,
            in2 => \_gnd_net_\,
            in3 => \N__46695\,
            lcout => n4430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43708\,
            in1 => \N__44046\,
            in2 => \N__48527\,
            in3 => \N__41759\,
            lcout => \c0.n9276\,
            ltout => \c0.n9276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_827_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41545\,
            in1 => \N__44084\,
            in2 => \N__41525\,
            in3 => \N__45722\,
            lcout => \c0.n17623\,
            ltout => \c0.n17623_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15771_4_lut_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100000000"
        )
    port map (
            in0 => \N__47529\,
            in1 => \N__41522\,
            in2 => \N__41510\,
            in3 => \N__49323\,
            lcout => OPEN,
            ltout => \c0.n17916_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0__3541_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47301\,
            in1 => \N__41507\,
            in2 => \N__41483\,
            in3 => \N__46697\,
            lcout => \c0.data_out_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50414\,
            ce => \N__44173\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1055_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__46694\,
            in1 => \N__49321\,
            in2 => \_gnd_net_\,
            in3 => \N__47298\,
            lcout => \c0.n8486\,
            ltout => \c0.n8486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_920_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__42248\,
            in1 => \N__42047\,
            in2 => \N__41435\,
            in3 => \N__41432\,
            lcout => n4_adj_2612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15690_2_lut_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47402\,
            lcout => OPEN,
            ltout => \c0.n17925_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5__3536_LC_13_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__44368\,
            in1 => \N__49328\,
            in2 => \N__41393\,
            in3 => \N__46878\,
            lcout => \c0.data_out_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50419\,
            ce => \N__44188\,
            sr => \_gnd_net_\
        );

    \c0.i15673_2_lut_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41717\,
            in2 => \_gnd_net_\,
            in3 => \N__47401\,
            lcout => OPEN,
            ltout => \c0.n17931_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4__3537_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__41668\,
            in1 => \N__49327\,
            in2 => \N__41699\,
            in3 => \N__46877\,
            lcout => \c0.data_out_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50419\,
            ce => \N__44188\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_833_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41648\,
            in2 => \_gnd_net_\,
            in3 => \N__45590\,
            lcout => \c0.n8812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43413\,
            in1 => \N__46448\,
            in2 => \N__47711\,
            in3 => \N__44051\,
            lcout => \c0.n17499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_871_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46449\,
            in1 => \N__43230\,
            in2 => \N__41696\,
            in3 => \N__48526\,
            lcout => \c0.data_out_7__4__N_550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_890_LC_13_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46079\,
            lcout => \c0.n6_adj_2451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15713_4_lut_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111001"
        )
    port map (
            in0 => \N__44123\,
            in1 => \N__41622\,
            in2 => \N__49445\,
            in3 => \N__43769\,
            lcout => OPEN,
            ltout => \c0.n17967_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__4__3553_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__41591\,
            in1 => \N__46899\,
            in2 => \N__41570\,
            in3 => \N__47404\,
            lcout => \c0.data_out_7__4__N_556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50424\,
            ce => \N__46564\,
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1114_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49808\,
            in1 => \N__43648\,
            in2 => \N__41567\,
            in3 => \N__41555\,
            lcout => \c0.n17662\,
            ltout => \c0.n17662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_702_i1_4_lut_LC_13_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__49418\,
            in1 => \N__45779\,
            in2 => \N__41888\,
            in3 => \N__49519\,
            lcout => OPEN,
            ltout => \c0.n2041_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7__3542_LC_13_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47403\,
            in1 => \N__41885\,
            in2 => \N__41864\,
            in3 => \N__46914\,
            lcout => \c0.data_out_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50424\,
            ce => \N__46564\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1084_LC_13_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45625\,
            in1 => \N__48590\,
            in2 => \_gnd_net_\,
            in3 => \N__43226\,
            lcout => \c0.n17611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__7__3550_LC_13_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__49326\,
            in1 => \N__49730\,
            in2 => \N__46919\,
            in3 => \N__41861\,
            lcout => \c0.data_out_7__7__N_519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50427\,
            ce => \N__46565\,
            sr => \_gnd_net_\
        );

    \c0.mux_884_i1_4_lut_LC_13_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47753\,
            in1 => \N__49325\,
            in2 => \N__47537\,
            in3 => \N__44069\,
            lcout => OPEN,
            ltout => \c0.n17693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0__3549_LC_13_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000001111"
        )
    port map (
            in0 => \N__47405\,
            in1 => \N__41849\,
            in2 => \N__41828\,
            in3 => \N__46900\,
            lcout => \c0.data_out_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50427\,
            ce => \N__46565\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1123_LC_13_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43672\,
            lcout => \c0.n17578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4518_2_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42127\,
            lcout => n6878,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1039_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42065\,
            in1 => \N__41935\,
            in2 => \N__41975\,
            in3 => \N__41744\,
            lcout => \c0.n14_adj_2533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_1152_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47235\,
            in1 => \N__42572\,
            in2 => \_gnd_net_\,
            in3 => \N__42154\,
            lcout => n17364,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1030_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101111111"
        )
    port map (
            in0 => \N__46785\,
            in1 => \N__42143\,
            in2 => \N__49364\,
            in3 => \N__42110\,
            lcout => OPEN,
            ltout => \n17672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i0_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__47240\,
            in1 => \N__42778\,
            in2 => \N__42131\,
            in3 => \N__42011\,
            lcout => \UART_TRANSMITTER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5065_3_lut_4_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__42553\,
            in1 => \N__42128\,
            in2 => \N__49363\,
            in3 => \N__42109\,
            lcout => \c0.n7428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i12_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42448\,
            in1 => \N__42095\,
            in2 => \_gnd_net_\,
            in3 => \N__42081\,
            lcout => \c0.delay_counter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1005_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42932\,
            in1 => \N__42554\,
            in2 => \N__42986\,
            in3 => \N__42048\,
            lcout => OPEN,
            ltout => \UART_TRANSMITTER_state_7_N_1749_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15721_4_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__46724\,
            in1 => \N__49304\,
            in2 => \N__42014\,
            in3 => \N__47236\,
            lcout => n18032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1027_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__46723\,
            in1 => \N__42005\,
            in2 => \N__47142\,
            in3 => \N__41990\,
            lcout => n16485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15304_4_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42379\,
            in1 => \N__42354\,
            in2 => \N__41974\,
            in3 => \N__41931\,
            lcout => \c0.n17753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_i0_i7_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__42375\,
            in1 => \N__42568\,
            in2 => \N__42461\,
            in3 => \N__42449\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1037_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42374\,
            in2 => \_gnd_net_\,
            in3 => \N__42353\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1040_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42335\,
            in1 => \N__42296\,
            in2 => \N__42275\,
            in3 => \N__42272\,
            lcout => n17306,
            ltout => \n17306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1041_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42251\,
            in3 => \N__42241\,
            lcout => \c0.n6_adj_2534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48675\,
            in1 => \N__42205\,
            in2 => \_gnd_net_\,
            in3 => \N__42218\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_873_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__49291\,
            in1 => \N__46672\,
            in2 => \_gnd_net_\,
            in3 => \N__43006\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_874_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__43079\,
            in1 => \N__42602\,
            in2 => \N__42191\,
            in3 => \N__42836\,
            lcout => OPEN,
            ltout => \c0.n19_adj_2446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_3509_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__47276\,
            in1 => \N__42874\,
            in2 => \N__42188\,
            in3 => \N__42183\,
            lcout => \c0.tx_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50396\,
            ce => 'H',
            sr => \N__47144\
        );

    \c0.i11059_2_lut_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49290\,
            lcout => \c0.n2650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1112_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__43068\,
            in1 => \N__43050\,
            in2 => \_gnd_net_\,
            in3 => \N__43026\,
            lcout => \c0.n97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11030_2_lut_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42950\,
            in2 => \_gnd_net_\,
            in3 => \N__42931\,
            lcout => n13415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15888_2_lut_3_lut_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__46670\,
            in1 => \N__49289\,
            in2 => \_gnd_net_\,
            in3 => \N__47275\,
            lcout => \data_out_10__7__N_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__48738\,
            in1 => \N__42837\,
            in2 => \N__42713\,
            in3 => \N__42744\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48661\,
            in1 => \N__42793\,
            in2 => \_gnd_net_\,
            in3 => \N__44339\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state_i0_i1_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__42779\,
            in1 => \N__46646\,
            in2 => \N__42764\,
            in3 => \N__47341\,
            lcout => \UART_TRANSMITTER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__42745\,
            in1 => \N__42712\,
            in2 => \N__42635\,
            in3 => \N__42616\,
            lcout => byte_transmit_counter_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15292_2_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46645\,
            in2 => \_gnd_net_\,
            in3 => \N__42601\,
            lcout => \c0.n17741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48660\,
            in1 => \N__43180\,
            in2 => \_gnd_net_\,
            in3 => \N__44318\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47635\,
            in1 => \N__43810\,
            in2 => \_gnd_net_\,
            in3 => \N__48429\,
            lcout => \c0.n1_adj_2522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15800_2_lut_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43106\,
            lcout => \c0.n18071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43100\,
            in1 => \N__43333\,
            in2 => \_gnd_net_\,
            in3 => \N__48416\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15802_4_lut_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__43166\,
            in1 => \N__48134\,
            in2 => \N__43160\,
            in3 => \N__47974\,
            lcout => \c0.n18072\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_858_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49792\,
            in1 => \N__48589\,
            in2 => \N__43145\,
            in3 => \N__43589\,
            lcout => \c0.data_out_7__2__N_574\,
            ltout => \c0.data_out_7__2__N_574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__2__3515_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43490\,
            in1 => \N__46310\,
            in2 => \N__43109\,
            in3 => \N__45834\,
            lcout => \c0.data_out_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50409\,
            ce => \N__46008\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__2__3523_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__43811\,
            in1 => \N__49637\,
            in2 => \_gnd_net_\,
            in3 => \N__44138\,
            lcout => \c0.data_out_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50409\,
            ce => \N__46008\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43094\,
            in1 => \N__49566\,
            in2 => \_gnd_net_\,
            in3 => \N__48402\,
            lcout => \c0.n8_adj_2531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15803_2_lut_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45800\,
            lcout => OPEN,
            ltout => \c0.n18073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15828_4_lut_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__44453\,
            in1 => \N__48163\,
            in2 => \N__43358\,
            in3 => \N__47985\,
            lcout => \c0.n18014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__3__3530_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49567\,
            in1 => \N__46022\,
            in2 => \_gnd_net_\,
            in3 => \N__43355\,
            lcout => data_out_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1063_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43334\,
            in1 => \N__49565\,
            in2 => \_gnd_net_\,
            in3 => \N__43301\,
            lcout => \c0.n9091\,
            ltout => \c0.n9091_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1064_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43280\,
            in3 => \N__43466\,
            lcout => OPEN,
            ltout => \c0.n17566_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1066_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44512\,
            in1 => \N__48591\,
            in2 => \N__43277\,
            in3 => \N__43270\,
            lcout => \c0.n9195\,
            ltout => \c0.n9195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1070_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43235\,
            in3 => \N__43232\,
            lcout => \c0.n17608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15806_4_lut_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__48155\,
            in1 => \N__43427\,
            in2 => \N__43190\,
            in3 => \N__47983\,
            lcout => \c0.n18015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43439\,
            in1 => \N__47833\,
            in2 => \_gnd_net_\,
            in3 => \N__48418\,
            lcout => \c0.n8_adj_2516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1073_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49633\,
            in2 => \_gnd_net_\,
            in3 => \N__43528\,
            lcout => \c0.n17668\,
            ltout => \c0.n17668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__43499\,
            in1 => \_gnd_net_\,
            in2 => \N__43493\,
            in3 => \N__43486\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__0__3517_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46112\,
            in1 => \N__47533\,
            in2 => \N__43475\,
            in3 => \N__43472\,
            lcout => \c0.data_out_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50420\,
            ce => \N__46035\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__0__3525_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__47769\,
            in1 => \N__44419\,
            in2 => \_gnd_net_\,
            in3 => \N__43465\,
            lcout => \c0.data_out_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50420\,
            ce => \N__46035\,
            sr => \_gnd_net_\
        );

    \c0.i15843_2_lut_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48419\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43433\,
            lcout => \c0.n18016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1056_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49872\,
            in1 => \N__43584\,
            in2 => \N__44272\,
            in3 => \N__43655\,
            lcout => \c0.data_out_6__5__N_752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1097_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47703\,
            in2 => \_gnd_net_\,
            in3 => \N__46447\,
            lcout => OPEN,
            ltout => \c0.n4_adj_2543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_754_i1_4_lut_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__46255\,
            in1 => \N__43420\,
            in2 => \N__43361\,
            in3 => \N__49414\,
            lcout => OPEN,
            ltout => \c0.n9656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5__3544_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101100000011"
        )
    port map (
            in0 => \N__43889\,
            in1 => \N__46902\,
            in2 => \N__43868\,
            in3 => \N__47410\,
            lcout => \c0.data_out_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50425\,
            ce => \N__46547\,
            sr => \_gnd_net_\
        );

    \c0.mux_858_i1_4_lut_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100101"
        )
    port map (
            in0 => \N__43661\,
            in1 => \N__43825\,
            in2 => \N__49487\,
            in3 => \N__49415\,
            lcout => OPEN,
            ltout => \c0.n2251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1__3548_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__43865\,
            in1 => \N__46901\,
            in2 => \N__43841\,
            in3 => \N__47409\,
            lcout => \c0.data_out_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50425\,
            ce => \N__46547\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1065_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44388\,
            in2 => \_gnd_net_\,
            in3 => \N__46275\,
            lcout => \c0.n17510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1__3556_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__49416\,
            in1 => \N__43838\,
            in2 => \N__43829\,
            in3 => \N__46903\,
            lcout => \c0.data_out_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50425\,
            ce => \N__46547\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_892_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43797\,
            in1 => \N__47768\,
            in2 => \N__43771\,
            in3 => \N__43947\,
            lcout => \c0.n8767\,
            ltout => \c0.n8767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_836_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43721\,
            in3 => \N__49868\,
            lcout => \c0.n17457\,
            ltout => \c0.n17457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43718\,
            in1 => \N__43709\,
            in2 => \N__43682\,
            in3 => \N__43679\,
            lcout => \c0.n17415\,
            ltout => \c0.n17415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_999_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43646\,
            in1 => \N__44264\,
            in2 => \N__43592\,
            in3 => \N__43580\,
            lcout => \c0.n17659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__1__3540_LC_14_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__49163\,
            in1 => \N__46786\,
            in2 => \N__44219\,
            in3 => \N__47411\,
            lcout => \c0.data_out_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50428\,
            ce => \N__44186\,
            sr => \_gnd_net_\
        );

    \c0.data_out_3__0__3573_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__47110\,
            in1 => \N__44124\,
            in2 => \N__47449\,
            in3 => \N__47476\,
            lcout => \data_out_6__2__N_804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1068_LC_14_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46378\,
            in1 => \N__44080\,
            in2 => \_gnd_net_\,
            in3 => \N__49744\,
            lcout => \c0.n17654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15781_4_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__45875\,
            in1 => \N__48148\,
            in2 => \N__43961\,
            in3 => \N__47970\,
            lcout => \c0.n18061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15694_2_lut_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44050\,
            in2 => \_gnd_net_\,
            in3 => \N__48430\,
            lcout => \c0.n17943\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48431\,
            in1 => \N__46440\,
            in2 => \_gnd_net_\,
            in3 => \N__44015\,
            lcout => \c0.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15746_2_lut_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45758\,
            in2 => \_gnd_net_\,
            in3 => \N__48432\,
            lcout => \c0.n18060\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15784_2_lut_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__43948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48428\,
            lcout => \c0.n18091\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15791_4_lut_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__46235\,
            in1 => \N__48151\,
            in2 => \N__45857\,
            in3 => \N__47968\,
            lcout => OPEN,
            ltout => \c0.n18065_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11411_4_lut_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__48840\,
            in1 => \N__44279\,
            in2 => \N__44342\,
            in3 => \N__48736\,
            lcout => \tx_data_5_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1029_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__48737\,
            in1 => \N__44225\,
            in2 => \N__44330\,
            in3 => \N__48839\,
            lcout => \tx_data_1_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45596\,
            in1 => \N__46280\,
            in2 => \_gnd_net_\,
            in3 => \N__48427\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2481_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15955_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__44312\,
            in1 => \N__48149\,
            in2 => \N__44303\,
            in3 => \N__47967\,
            lcout => OPEN,
            ltout => \c0.n18402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18402_bdd_4_lut_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48150\,
            in1 => \N__44300\,
            in2 => \N__44294\,
            in3 => \N__44291\,
            lcout => \c0.n18405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i59_3_lut_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46309\,
            in1 => \N__44395\,
            in2 => \_gnd_net_\,
            in3 => \N__48464\,
            lcout => OPEN,
            ltout => \c0.n45_adj_2518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i60_4_lut_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__48466\,
            in1 => \N__44273\,
            in2 => \N__44240\,
            in3 => \N__47972\,
            lcout => OPEN,
            ltout => \c0.n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i58_4_lut_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__47973\,
            in1 => \N__44237\,
            in2 => \N__44228\,
            in3 => \N__48136\,
            lcout => \c0.n44_adj_2524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_840_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47704\,
            in2 => \_gnd_net_\,
            in3 => \N__47636\,
            lcout => \c0.n8777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15797_2_lut_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48465\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45542\,
            lcout => OPEN,
            ltout => \c0.n18069_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15799_4_lut_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__47971\,
            in1 => \N__45533\,
            in2 => \N__45527\,
            in3 => \N__48135\,
            lcout => \c0.n18070\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i111_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44944\,
            in1 => \N__44533\,
            in2 => \_gnd_net_\,
            in3 => \N__44561\,
            lcout => data_in_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__1__3524_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49549\,
            in1 => \N__44522\,
            in2 => \N__47783\,
            in3 => \N__44513\,
            lcout => \c0.data_out_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50421\,
            ce => \N__46015\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44495\,
            in1 => \N__44488\,
            in2 => \_gnd_net_\,
            in3 => \N__48467\,
            lcout => \c0.n8_adj_2519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44402\,
            in1 => \N__49616\,
            in2 => \_gnd_net_\,
            in3 => \N__48468\,
            lcout => \c0.n8_adj_2535\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__4__3521_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45913\,
            in1 => \N__44435\,
            in2 => \N__44423\,
            in3 => \N__45838\,
            lcout => \c0.data_out_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50421\,
            ce => \N__46015\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__5__3512_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__47779\,
            in1 => \N__44396\,
            in2 => \N__44375\,
            in3 => \N__44354\,
            lcout => \c0.data_out_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50421\,
            ce => \N__46015\,
            sr => \_gnd_net_\
        );

    \c0.i15788_2_lut_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45863\,
            in2 => \_gnd_net_\,
            in3 => \N__48469\,
            lcout => \c0.n18064\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45599\,
            in1 => \N__45845\,
            in2 => \N__45839\,
            in3 => \N__45657\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__1__3516_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49476\,
            in1 => \N__49505\,
            in2 => \N__45803\,
            in3 => \N__46198\,
            lcout => \c0.data_out_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50426\,
            ce => \N__46036\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__7__3510_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45557\,
            in1 => \N__45794\,
            in2 => \_gnd_net_\,
            in3 => \N__45778\,
            lcout => \c0.data_out_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50426\,
            ce => \N__46036\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_863_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49783\,
            in1 => \N__45745\,
            in2 => \_gnd_net_\,
            in3 => \N__45721\,
            lcout => \c0.n17635\,
            ltout => \c0.n17635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15674_3_lut_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45655\,
            in2 => \N__45680\,
            in3 => \N__49397\,
            lcout => \c0.n17922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1032_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45656\,
            in1 => \N__45598\,
            in2 => \_gnd_net_\,
            in3 => \N__48208\,
            lcout => \c0.n17492\,
            ltout => \c0.n17492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__3__3514_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46286\,
            in1 => \N__45551\,
            in2 => \N__45545\,
            in3 => \N__46364\,
            lcout => \c0.data_out_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50426\,
            ce => \N__46036\,
            sr => \_gnd_net_\
        );

    \c0.data_out_9__6__3519_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46183\,
            in1 => \N__46367\,
            in2 => \N__46328\,
            in3 => \N__49708\,
            lcout => \c0.data_out_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50429\,
            ce => \N__46037\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46316\,
            in1 => \N__46150\,
            in2 => \_gnd_net_\,
            in3 => \N__48458\,
            lcout => \c0.n8_adj_2539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_997_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45912\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46302\,
            lcout => \c0.n17454\,
            ltout => \c0.n17454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__5__3520_LC_15_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__46279\,
            in1 => \N__46256\,
            in2 => \N__46244\,
            in3 => \N__49550\,
            lcout => \c0.data_out_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50429\,
            ce => \N__46037\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48459\,
            in1 => \N__46241\,
            in2 => \_gnd_net_\,
            in3 => \N__49707\,
            lcout => \c0.n8_adj_2537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_949_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46223\,
            in1 => \N__46199\,
            in2 => \N__46184\,
            in3 => \N__46163\,
            lcout => OPEN,
            ltout => \c0.n12_adj_2482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__7__3518_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46151\,
            in1 => \N__46105\,
            in2 => \N__46091\,
            in3 => \N__46088\,
            lcout => \c0.data_out_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50429\,
            ce => \N__46037\,
            sr => \_gnd_net_\
        );

    \c0.i10536_3_lut_LC_15_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45920\,
            in1 => \N__45911\,
            in2 => \_gnd_net_\,
            in3 => \N__48457\,
            lcout => \c0.n8_adj_2538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46978\,
            in1 => \N__47770\,
            in2 => \_gnd_net_\,
            in3 => \N__48473\,
            lcout => \c0.n1_adj_2484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1124_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47695\,
            in1 => \N__47640\,
            in2 => \_gnd_net_\,
            in3 => \N__47578\,
            lcout => \c0.n8926\,
            ltout => \c0.n8926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1109_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47507\,
            in2 => \N__47501\,
            in3 => \N__46976\,
            lcout => \c0.n17438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_1207_i1_3_lut_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49384\,
            in1 => \N__46800\,
            in2 => \_gnd_net_\,
            in3 => \N__47412\,
            lcout => n2720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__6__3583_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__47413\,
            in1 => \N__46977\,
            in2 => \N__47134\,
            in3 => \N__46804\,
            lcout => data_out_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46955\,
            in1 => \N__48502\,
            in2 => \_gnd_net_\,
            in3 => \N__46451\,
            lcout => \c0.data_out_6__3__N_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__6__3567_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__48503\,
            in1 => \N__49385\,
            in2 => \N__46881\,
            in3 => \N__46531\,
            lcout => data_out_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4__I_567_2_lut_LC_15_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48501\,
            in2 => \_gnd_net_\,
            in3 => \N__46450\,
            lcout => \c0.data_out_6__4__N_765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15965_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__48533\,
            in1 => \N__48158\,
            in2 => \N__48182\,
            in3 => \N__47987\,
            lcout => OPEN,
            ltout => \c0.n18414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18414_bdd_4_lut_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48159\,
            in1 => \N__48860\,
            in2 => \N__48848\,
            in3 => \N__48479\,
            lcout => OPEN,
            ltout => \c0.n18417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11407_4_lut_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__48838\,
            in1 => \N__47846\,
            in2 => \N__48764\,
            in3 => \N__48760\,
            lcout => OPEN,
            ltout => \tx_data_6_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__48682\,
            in1 => \_gnd_net_\,
            in2 => \N__48617\,
            in3 => \N__48607\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15698_2_lut_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48593\,
            in2 => \_gnd_net_\,
            in3 => \N__48461\,
            lcout => \c0.n17949\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15720_2_lut_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48522\,
            lcout => \c0.n18090\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48462\,
            in1 => \N__49663\,
            in2 => \_gnd_net_\,
            in3 => \N__48209\,
            lcout => \c0.n5_adj_2444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15787_4_lut_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__48173\,
            in1 => \N__48157\,
            in2 => \N__47999\,
            in3 => \N__47986\,
            lcout => \c0.n18063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_888_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47840\,
            in2 => \_gnd_net_\,
            in3 => \N__47807\,
            lcout => \c0.n17638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i0_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48932\,
            in2 => \_gnd_net_\,
            in3 => \N__48926\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_16_29_0_\,
            carryout => n16380,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i1_LC_16_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48923\,
            in2 => \_gnd_net_\,
            in3 => \N__48917\,
            lcout => n25,
            ltout => OPEN,
            carryin => n16380,
            carryout => n16381,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i2_LC_16_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48914\,
            in2 => \_gnd_net_\,
            in3 => \N__48908\,
            lcout => n24,
            ltout => OPEN,
            carryin => n16381,
            carryout => n16382,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i3_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48905\,
            in2 => \_gnd_net_\,
            in3 => \N__48899\,
            lcout => n23,
            ltout => OPEN,
            carryin => n16382,
            carryout => n16383,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i4_LC_16_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48896\,
            in2 => \_gnd_net_\,
            in3 => \N__48890\,
            lcout => n22_adj_2655,
            ltout => OPEN,
            carryin => n16383,
            carryout => n16384,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i5_LC_16_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48887\,
            in2 => \_gnd_net_\,
            in3 => \N__48881\,
            lcout => n21,
            ltout => OPEN,
            carryin => n16384,
            carryout => n16385,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i6_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48878\,
            in2 => \_gnd_net_\,
            in3 => \N__48872\,
            lcout => n20,
            ltout => OPEN,
            carryin => n16385,
            carryout => n16386,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i7_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48869\,
            in2 => \_gnd_net_\,
            in3 => \N__48863\,
            lcout => n19,
            ltout => OPEN,
            carryin => n16386,
            carryout => n16387,
            clk => \N__50430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i8_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49010\,
            in2 => \_gnd_net_\,
            in3 => \N__49004\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_16_30_0_\,
            carryout => n16388,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i9_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49001\,
            in2 => \_gnd_net_\,
            in3 => \N__48995\,
            lcout => n17,
            ltout => OPEN,
            carryin => n16388,
            carryout => n16389,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i10_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48992\,
            in2 => \_gnd_net_\,
            in3 => \N__48986\,
            lcout => n16,
            ltout => OPEN,
            carryin => n16389,
            carryout => n16390,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i11_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48983\,
            in2 => \_gnd_net_\,
            in3 => \N__48977\,
            lcout => n15,
            ltout => OPEN,
            carryin => n16390,
            carryout => n16391,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i12_LC_16_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48974\,
            in2 => \_gnd_net_\,
            in3 => \N__48968\,
            lcout => n14,
            ltout => OPEN,
            carryin => n16391,
            carryout => n16392,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i13_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48965\,
            in2 => \_gnd_net_\,
            in3 => \N__48959\,
            lcout => n13,
            ltout => OPEN,
            carryin => n16392,
            carryout => n16393,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i14_LC_16_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48956\,
            in2 => \_gnd_net_\,
            in3 => \N__48950\,
            lcout => n12,
            ltout => OPEN,
            carryin => n16393,
            carryout => n16394,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i15_LC_16_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48947\,
            in2 => \_gnd_net_\,
            in3 => \N__48941\,
            lcout => n11,
            ltout => OPEN,
            carryin => n16394,
            carryout => n16395,
            clk => \N__50433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i16_LC_16_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48938\,
            in2 => \_gnd_net_\,
            in3 => \N__49151\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_16_31_0_\,
            carryout => n16396,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i17_LC_16_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49148\,
            in2 => \_gnd_net_\,
            in3 => \N__49142\,
            lcout => n9,
            ltout => OPEN,
            carryin => n16396,
            carryout => n16397,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i18_LC_16_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49139\,
            in2 => \_gnd_net_\,
            in3 => \N__49133\,
            lcout => n8_adj_2617,
            ltout => OPEN,
            carryin => n16397,
            carryout => n16398,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i19_LC_16_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49130\,
            in2 => \_gnd_net_\,
            in3 => \N__49124\,
            lcout => n7,
            ltout => OPEN,
            carryin => n16398,
            carryout => n16399,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i20_LC_16_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49121\,
            in2 => \_gnd_net_\,
            in3 => \N__49115\,
            lcout => n6,
            ltout => OPEN,
            carryin => n16399,
            carryout => n16400,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i21_LC_16_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49102\,
            in2 => \_gnd_net_\,
            in3 => \N__49091\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n16400,
            carryout => n16401,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i22_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49078\,
            in2 => \_gnd_net_\,
            in3 => \N__49067\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n16401,
            carryout => n16402,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i23_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49057\,
            in2 => \_gnd_net_\,
            in3 => \N__49046\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n16402,
            carryout => n16403,
            clk => \N__50434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i24_LC_16_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49024\,
            in2 => \_gnd_net_\,
            in3 => \N__49013\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_16_32_0_\,
            carryout => n16404,
            clk => \N__50435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2271__i25_LC_16_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50446\,
            in2 => \_gnd_net_\,
            in3 => \N__50462\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15672_4_lut_LC_16_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49873\,
            in1 => \N__49807\,
            in2 => \N__49793\,
            in3 => \N__49748\,
            lcout => \c0.n17976\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1054_LC_17_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49610\,
            in1 => \N__49721\,
            in2 => \N__49709\,
            in3 => \N__49667\,
            lcout => \c0.n8922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_929_LC_17_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49611\,
            in2 => \_gnd_net_\,
            in3 => \N__49574\,
            lcout => \c0.n17620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15663_4_lut_LC_18_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100000000"
        )
    port map (
            in0 => \N__49526\,
            in1 => \N__49504\,
            in2 => \N__49486\,
            in3 => \N__49436\,
            lcout => \c0.n17918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
